magic
tech scmos
magscale 1 2
timestamp 1720180704
<< metal1 >>
rect -63 6258 -3 6518
rect 6930 6502 7023 6518
rect 6507 6417 6593 6423
rect 3987 6357 4073 6363
rect 4947 6357 4993 6363
rect 6387 6357 6453 6363
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 277 6223 283 6243
rect 247 6217 283 6223
rect 5507 6157 5613 6163
rect 1687 6137 1733 6143
rect 2507 6137 2593 6143
rect 3087 6137 3233 6143
rect 4447 6137 4513 6143
rect 6067 6137 6113 6143
rect 5707 6117 5733 6123
rect 2667 6057 2733 6063
rect 3947 6057 3973 6063
rect 6327 6057 6393 6063
rect 4827 6037 4873 6043
rect 6963 5998 7023 6502
rect 6930 5982 7023 5998
rect 4947 5957 4993 5963
rect 4627 5937 4693 5943
rect 5147 5937 5173 5943
rect 3407 5917 3453 5923
rect 2987 5897 3033 5903
rect 3287 5897 3333 5903
rect 3427 5903 3440 5907
rect 3427 5893 3443 5903
rect 4247 5897 4273 5903
rect 1567 5877 1633 5883
rect 3437 5867 3443 5893
rect 3427 5857 3443 5867
rect 3427 5853 3440 5857
rect 4787 5857 4833 5863
rect 3547 5837 3693 5843
rect 3887 5837 3933 5843
rect 4027 5837 4093 5843
rect 4227 5837 4333 5843
rect 4587 5837 4693 5843
rect 5247 5837 5272 5843
rect 5307 5837 5373 5843
rect 5967 5837 6053 5843
rect 6527 5837 6593 5843
rect 6347 5817 6453 5823
rect 6307 5797 6413 5803
rect 5307 5777 5333 5783
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 1927 5637 2073 5643
rect 2127 5637 2233 5643
rect 2127 5617 2193 5623
rect 2747 5617 2793 5623
rect 4627 5617 4673 5623
rect 4787 5617 4873 5623
rect 6167 5617 6213 5623
rect 6540 5623 6553 5627
rect 6537 5614 6553 5623
rect 6537 5613 6560 5614
rect 1000 5603 1013 5607
rect 997 5593 1013 5603
rect 3107 5603 3120 5607
rect 3107 5593 3123 5603
rect 6467 5603 6480 5607
rect 6537 5603 6543 5613
rect 6467 5593 6483 5603
rect 997 5567 1003 5593
rect 3117 5567 3123 5593
rect 6477 5567 6483 5593
rect 997 5557 1013 5567
rect 1000 5553 1013 5557
rect 3107 5557 3123 5567
rect 3107 5553 3120 5557
rect 4847 5557 4893 5563
rect 5647 5557 5673 5563
rect 5767 5557 5793 5563
rect 6467 5557 6483 5567
rect 6517 5597 6543 5603
rect 6517 5567 6523 5597
rect 6517 5557 6533 5567
rect 6467 5553 6480 5557
rect 6520 5553 6533 5557
rect 3947 5537 4013 5543
rect 4127 5537 4173 5543
rect 4847 5537 4993 5543
rect 867 5517 893 5523
rect 6963 5478 7023 5982
rect 6930 5462 7023 5478
rect 3167 5437 3193 5443
rect 2627 5417 2653 5423
rect 3927 5397 3993 5403
rect 5507 5397 5593 5403
rect 5867 5397 5933 5403
rect 5987 5397 6073 5403
rect 667 5383 680 5387
rect 667 5373 683 5383
rect 5307 5383 5320 5387
rect 6380 5383 6393 5387
rect 5307 5373 5323 5383
rect 677 5343 683 5373
rect 677 5337 733 5343
rect 1667 5337 1693 5343
rect 2087 5317 2113 5323
rect 4727 5317 4793 5323
rect 5317 5323 5323 5373
rect 6377 5373 6393 5383
rect 6667 5383 6680 5387
rect 6667 5373 6683 5383
rect 6377 5347 6383 5373
rect 6677 5347 6683 5373
rect 6377 5337 6393 5347
rect 6380 5333 6393 5337
rect 6667 5337 6683 5347
rect 6667 5333 6680 5337
rect 5317 5317 5393 5323
rect 5487 5317 5573 5323
rect 5667 5317 5773 5323
rect 5887 5317 5933 5323
rect 6287 5317 6353 5323
rect 6697 5323 6703 5393
rect 6720 5383 6733 5387
rect 6717 5373 6733 5383
rect 6847 5383 6860 5387
rect 6847 5373 6863 5383
rect 6717 5347 6723 5373
rect 6717 5337 6733 5347
rect 6720 5333 6733 5337
rect 6697 5317 6753 5323
rect 6857 5323 6863 5373
rect 6827 5317 6863 5323
rect 2367 5297 2393 5303
rect 5433 5303 5447 5313
rect 5327 5300 5447 5303
rect 5327 5297 5443 5300
rect 6447 5297 6533 5303
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 5787 5117 5833 5123
rect 1367 5097 1393 5103
rect 3007 5097 3073 5103
rect 3907 5097 3933 5103
rect 2877 5077 2933 5083
rect 367 5017 513 5023
rect 627 5017 793 5023
rect 2877 5026 2883 5077
rect 4707 5083 4720 5087
rect 4707 5073 4723 5083
rect 5007 5083 5020 5087
rect 5007 5073 5023 5083
rect 5667 5077 5713 5083
rect 4717 5047 4723 5073
rect 4707 5037 4723 5047
rect 5017 5043 5023 5073
rect 5017 5037 5073 5043
rect 4707 5033 4720 5037
rect 5467 5037 5513 5043
rect 3167 5017 3193 5023
rect 3547 5017 3613 5023
rect 6137 5007 6143 5113
rect 6467 5097 6513 5103
rect 6427 5077 6483 5083
rect 6453 5043 6467 5053
rect 6427 5040 6467 5043
rect 6477 5047 6483 5077
rect 6597 5077 6653 5083
rect 6597 5047 6603 5077
rect 6427 5037 6463 5040
rect 6477 5037 6493 5047
rect 6480 5033 6493 5037
rect 6587 5037 6603 5047
rect 6587 5033 6600 5037
rect 6797 5007 6803 5093
rect 667 4997 773 5003
rect 6797 5006 6820 5007
rect 6797 4997 6813 5006
rect 6800 4993 6813 4997
rect 6963 4958 7023 5462
rect 6930 4942 7023 4958
rect 5067 4917 5113 4923
rect 5907 4897 5973 4903
rect 787 4877 893 4883
rect 1627 4877 1733 4883
rect 2127 4877 2173 4883
rect 4167 4877 4273 4883
rect 5907 4877 5973 4883
rect 6047 4877 6133 4883
rect 6407 4877 6473 4883
rect 6567 4877 6613 4883
rect 2567 4857 2613 4863
rect 3547 4857 3573 4863
rect 4397 4857 4453 4863
rect 4397 4827 4403 4857
rect 5047 4863 5060 4867
rect 5280 4863 5293 4867
rect 5047 4853 5063 4863
rect 4877 4837 4913 4843
rect 4877 4827 4883 4837
rect 5057 4827 5063 4853
rect 5277 4853 5293 4863
rect 6217 4857 6273 4863
rect 5277 4827 5283 4853
rect 6217 4827 6223 4857
rect 6527 4857 6583 4863
rect 3867 4817 3913 4823
rect 4387 4817 4403 4827
rect 4387 4813 4400 4817
rect 4867 4817 4883 4827
rect 4867 4813 4880 4817
rect 5047 4817 5063 4827
rect 5047 4813 5060 4817
rect 5087 4817 5113 4823
rect 5277 4817 5293 4827
rect 5280 4813 5293 4817
rect 6207 4817 6223 4827
rect 6577 4827 6583 4857
rect 6847 4863 6860 4867
rect 6847 4853 6863 4863
rect 6857 4843 6863 4853
rect 6857 4837 6893 4843
rect 6577 4817 6593 4827
rect 6207 4813 6220 4817
rect 6580 4813 6593 4817
rect 2907 4797 2953 4803
rect 4347 4797 4473 4803
rect 4867 4797 4933 4803
rect 5367 4797 5513 4803
rect 5867 4797 5933 4803
rect 6027 4797 6133 4803
rect 6187 4797 6273 4803
rect 5067 4777 5133 4783
rect 5147 4777 5173 4783
rect 5227 4777 5293 4783
rect 6207 4777 6253 4783
rect 2547 4757 2613 4763
rect 4427 4757 4473 4763
rect 5227 4737 5273 4743
rect 3007 4717 3073 4723
rect 4387 4717 4453 4723
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 4207 4657 4273 4663
rect 4407 4657 4433 4663
rect 4927 4657 4973 4663
rect 4727 4617 4793 4623
rect 4747 4597 4813 4603
rect 5847 4597 5973 4603
rect 967 4577 1113 4583
rect 3227 4577 3253 4583
rect 4347 4577 4433 4583
rect 4507 4577 4573 4583
rect 4667 4577 4813 4583
rect 4867 4577 4973 4583
rect 5247 4577 5283 4583
rect 3027 4563 3040 4567
rect 4080 4563 4093 4567
rect 3027 4553 3043 4563
rect 3037 4527 3043 4553
rect 4077 4553 4093 4563
rect 4547 4563 4560 4567
rect 4600 4563 4613 4567
rect 4547 4553 4563 4563
rect 3027 4517 3043 4527
rect 3027 4513 3040 4517
rect 4077 4523 4083 4553
rect 4557 4527 4563 4553
rect 4027 4517 4083 4523
rect 4547 4517 4563 4527
rect 4597 4553 4613 4563
rect 4780 4563 4793 4567
rect 4777 4553 4793 4563
rect 5277 4563 5283 4577
rect 6067 4577 6093 4583
rect 6247 4577 6363 4583
rect 5277 4557 5313 4563
rect 5620 4563 5633 4567
rect 5617 4553 5633 4563
rect 5727 4563 5740 4567
rect 5727 4553 5743 4563
rect 4597 4527 4603 4553
rect 4777 4527 4783 4553
rect 5617 4543 5623 4553
rect 5587 4537 5623 4543
rect 5737 4527 5743 4553
rect 4597 4517 4613 4527
rect 4547 4513 4560 4517
rect 4600 4513 4613 4517
rect 4777 4517 4793 4527
rect 4780 4513 4793 4517
rect 5727 4517 5743 4527
rect 5757 4557 5793 4563
rect 5727 4513 5740 4517
rect 3647 4497 3673 4503
rect 3687 4497 3713 4503
rect 4907 4497 4953 4503
rect 5247 4497 5353 4503
rect 5407 4497 5493 4503
rect 5757 4503 5763 4557
rect 6327 4563 6340 4567
rect 6327 4553 6343 4563
rect 6337 4527 6343 4553
rect 6087 4517 6173 4523
rect 6327 4517 6343 4527
rect 6357 4523 6363 4577
rect 6847 4563 6860 4567
rect 6847 4553 6863 4563
rect 6857 4527 6863 4553
rect 6357 4517 6413 4523
rect 6327 4513 6340 4517
rect 6847 4517 6863 4527
rect 6847 4513 6860 4517
rect 5707 4497 5763 4503
rect 6227 4497 6353 4503
rect 6487 4497 6513 4503
rect 4907 4477 4973 4483
rect 5407 4477 5453 4483
rect 5727 4477 5793 4483
rect 6527 4477 6593 4483
rect 1027 4457 1053 4463
rect 6963 4438 7023 4942
rect 6930 4422 7023 4438
rect 5887 4377 5913 4383
rect 2087 4357 2173 4363
rect 2827 4357 2873 4363
rect 5487 4357 5553 4363
rect 5713 4363 5727 4373
rect 5647 4360 5727 4363
rect 5647 4357 5723 4360
rect 6100 4363 6113 4367
rect 5807 4357 5863 4363
rect 1947 4337 1973 4343
rect 2327 4337 2373 4343
rect 4987 4337 5013 4343
rect 5400 4343 5413 4347
rect 5397 4333 5413 4343
rect 5507 4343 5520 4347
rect 5507 4333 5523 4343
rect 5687 4343 5700 4347
rect 5857 4343 5863 4357
rect 6097 4353 6113 4363
rect 6167 4357 6213 4363
rect 6357 4357 6433 4363
rect 6097 4343 6103 4353
rect 5687 4333 5703 4343
rect 5857 4337 5883 4343
rect 5397 4303 5403 4333
rect 5517 4323 5523 4333
rect 5517 4317 5563 4323
rect 5347 4297 5403 4303
rect 5557 4307 5563 4317
rect 5697 4307 5703 4333
rect 5557 4297 5573 4307
rect 5560 4293 5573 4297
rect 5687 4297 5703 4307
rect 5877 4303 5883 4337
rect 6077 4337 6103 4343
rect 5877 4297 5933 4303
rect 5687 4293 5700 4297
rect 6077 4303 6083 4337
rect 6027 4297 6083 4303
rect 6187 4297 6213 4303
rect 6357 4303 6363 4357
rect 6400 4343 6413 4347
rect 6337 4297 6363 4303
rect 6397 4333 6413 4343
rect 6507 4343 6520 4347
rect 6507 4333 6523 4343
rect 6547 4343 6560 4347
rect 6547 4333 6563 4343
rect 1527 4277 1693 4283
rect 4647 4277 4673 4283
rect 4727 4277 4833 4283
rect 4927 4277 5053 4283
rect 5127 4277 5233 4283
rect 5807 4277 5893 4283
rect 6167 4277 6273 4283
rect 6337 4283 6343 4297
rect 6397 4287 6403 4333
rect 6517 4327 6523 4333
rect 6517 4326 6540 4327
rect 6517 4317 6533 4326
rect 6520 4313 6533 4317
rect 6557 4307 6563 4333
rect 6557 4297 6573 4307
rect 6560 4293 6573 4297
rect 6667 4297 6713 4303
rect 6317 4280 6343 4283
rect 6313 4277 6343 4280
rect 4767 4257 4813 4263
rect 6313 4266 6327 4277
rect 6397 4283 6413 4287
rect 6367 4277 6413 4283
rect 6400 4273 6413 4277
rect 6487 4277 6593 4283
rect 6187 4257 6273 4263
rect 6007 4237 6073 4243
rect 5867 4217 5893 4223
rect 5147 4197 5213 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 2767 4077 2813 4083
rect 6127 4077 6233 4083
rect 6767 4077 6833 4083
rect 227 4057 273 4063
rect 1047 4057 1133 4063
rect 1547 4057 1593 4063
rect 1727 4057 1793 4063
rect 2687 4057 2833 4063
rect 3507 4057 3613 4063
rect 4727 4057 4753 4063
rect 4797 4057 4853 4063
rect 2367 4037 2393 4043
rect 4547 4043 4560 4047
rect 4547 4040 4563 4043
rect 4547 4033 4567 4040
rect 4553 4027 4567 4033
rect 4797 4007 4803 4057
rect 6427 4057 6513 4063
rect 6587 4057 6633 4063
rect 5360 4043 5373 4047
rect 5357 4033 5373 4043
rect 5627 4043 5640 4047
rect 5627 4033 5643 4043
rect 5827 4037 5853 4043
rect 6307 4037 6363 4043
rect 5357 4007 5363 4033
rect 5637 4007 5643 4033
rect 4740 4003 4753 4007
rect 4547 3997 4623 4003
rect 187 3977 213 3983
rect 1467 3977 1573 3983
rect 4327 3977 4353 3983
rect 4527 3977 4593 3983
rect 4617 3967 4623 3997
rect 4737 3993 4753 4003
rect 4797 3997 4813 4007
rect 4800 3993 4813 3997
rect 5357 3997 5373 4007
rect 5360 3993 5373 3997
rect 5507 3997 5533 4003
rect 5627 3997 5643 4007
rect 6357 4007 6363 4037
rect 6607 4037 6653 4043
rect 6357 3997 6373 4007
rect 5627 3993 5640 3997
rect 6360 3993 6373 3997
rect 4737 3963 4743 3993
rect 4767 3977 4853 3983
rect 5107 3977 5193 3983
rect 5447 3977 5553 3983
rect 5607 3977 5673 3983
rect 6737 3980 6773 3983
rect 6733 3977 6773 3980
rect 6733 3967 6747 3977
rect 6887 3977 6933 3983
rect 4737 3957 4813 3963
rect 5127 3957 5153 3963
rect 5467 3937 5533 3943
rect 5647 3937 5693 3943
rect 6963 3918 7023 4422
rect 6930 3902 7023 3918
rect 907 3837 953 3843
rect 2587 3837 2613 3843
rect 3067 3837 3153 3843
rect 3327 3837 3393 3843
rect 3447 3837 3553 3843
rect 6160 3843 6173 3847
rect 6157 3833 6173 3843
rect 2167 3817 2213 3823
rect 5607 3817 5653 3823
rect 5947 3823 5960 3827
rect 6157 3823 6163 3833
rect 6180 3823 6193 3827
rect 5947 3820 5963 3823
rect 5947 3813 5967 3820
rect 4380 3803 4393 3807
rect 4377 3793 4393 3803
rect 5953 3806 5967 3813
rect 3127 3777 3153 3783
rect 687 3757 793 3763
rect 1607 3757 1733 3763
rect 2047 3757 2113 3763
rect 2927 3757 2993 3763
rect 3067 3757 3173 3763
rect 4377 3766 4383 3793
rect 6137 3817 6163 3823
rect 6137 3787 6143 3817
rect 6127 3777 6143 3787
rect 6177 3813 6193 3823
rect 6497 3817 6553 3823
rect 6177 3787 6183 3813
rect 6497 3787 6503 3817
rect 6647 3817 6703 3823
rect 6177 3777 6193 3787
rect 6127 3773 6140 3777
rect 6180 3773 6193 3777
rect 6487 3777 6503 3787
rect 6697 3787 6703 3817
rect 6697 3777 6713 3787
rect 6487 3773 6500 3777
rect 6700 3773 6713 3777
rect 5707 3757 5853 3763
rect 5967 3757 6033 3763
rect 6087 3757 6123 3763
rect 5407 3737 5433 3743
rect 6117 3743 6123 3757
rect 6167 3757 6233 3763
rect 6117 3737 6213 3743
rect 6427 3737 6513 3743
rect 1847 3677 1893 3683
rect 4547 3677 4613 3683
rect 6647 3677 6673 3683
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 1307 3617 1353 3623
rect 1827 3597 1873 3603
rect 4627 3597 4693 3603
rect 6087 3597 6113 3603
rect 6587 3577 6613 3583
rect 2147 3557 2253 3563
rect 2767 3557 2793 3563
rect 5927 3557 6013 3563
rect 6467 3557 6493 3563
rect 6727 3557 6873 3563
rect 607 3537 753 3543
rect 3347 3537 3413 3543
rect 4467 3537 4513 3543
rect 4587 3537 4633 3543
rect 4807 3537 4893 3543
rect 5617 3537 5653 3543
rect 1180 3523 1193 3527
rect 1177 3513 1193 3523
rect 1467 3517 1513 3523
rect 4447 3517 4483 3523
rect 1177 3487 1183 3513
rect 4477 3503 4483 3517
rect 4477 3497 4503 3503
rect 4497 3487 4503 3497
rect 1177 3477 1193 3487
rect 1180 3473 1193 3477
rect 2047 3477 2073 3483
rect 3207 3477 3233 3483
rect 4497 3477 4513 3487
rect 4500 3473 4513 3477
rect 5227 3477 5293 3483
rect 5407 3477 5453 3483
rect 3147 3457 3213 3463
rect 5207 3457 5313 3463
rect 5577 3463 5583 3533
rect 5617 3487 5623 3537
rect 6227 3537 6333 3543
rect 6547 3537 6573 3543
rect 6587 3537 6653 3543
rect 6877 3543 6883 3553
rect 6727 3537 6783 3543
rect 6120 3523 6133 3527
rect 6117 3513 6133 3523
rect 6480 3523 6493 3527
rect 6477 3513 6493 3523
rect 6777 3523 6783 3537
rect 6837 3537 6883 3543
rect 6777 3517 6803 3523
rect 6117 3487 6123 3513
rect 6477 3487 6483 3513
rect 6797 3487 6803 3517
rect 5617 3477 5633 3487
rect 5620 3473 5633 3477
rect 6117 3477 6133 3487
rect 6120 3473 6133 3477
rect 6247 3477 6313 3483
rect 6477 3477 6493 3487
rect 6480 3473 6493 3477
rect 6787 3477 6803 3487
rect 6837 3487 6843 3537
rect 6837 3477 6853 3487
rect 6787 3473 6800 3477
rect 6840 3473 6853 3477
rect 5547 3457 5583 3463
rect 5607 3417 5633 3423
rect 6963 3398 7023 3902
rect 6930 3382 7023 3398
rect 6567 3357 6613 3363
rect 1267 3337 1293 3343
rect 1707 3337 1773 3343
rect 6427 3340 6483 3343
rect 6427 3337 6487 3340
rect 1127 3317 1153 3323
rect 1167 3317 1313 3323
rect 3147 3317 3253 3323
rect 4067 3317 4093 3323
rect 6473 3326 6487 3337
rect 5487 3317 5573 3323
rect 47 3297 93 3303
rect 1207 3297 1293 3303
rect 1687 3297 1733 3303
rect 2167 3297 2233 3303
rect 5457 3263 5463 3293
rect 5487 3297 5553 3303
rect 6387 3303 6400 3307
rect 6387 3293 6403 3303
rect 6427 3297 6453 3303
rect 6397 3283 6403 3293
rect 6397 3277 6443 3283
rect 6437 3267 6443 3277
rect 5457 3257 5553 3263
rect 6437 3257 6453 3267
rect 6440 3253 6453 3257
rect 767 3237 813 3243
rect 1147 3237 1233 3243
rect 1507 3237 1533 3243
rect 3367 3237 3453 3243
rect 5687 3237 5713 3243
rect 6247 3237 6273 3243
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 6847 3077 6913 3083
rect 5407 3057 5473 3063
rect 2507 3037 2533 3043
rect 2147 3017 2173 3023
rect 2827 3017 2853 3023
rect 3027 3017 3073 3023
rect 3327 3017 3393 3023
rect 4327 3017 4393 3023
rect 6807 3017 6913 3023
rect 4540 3003 4553 3007
rect 4537 3000 4553 3003
rect 4533 2993 4553 3000
rect 4700 3003 4713 3007
rect 4697 2993 4713 3003
rect 5277 2997 5353 3003
rect 4533 2987 4547 2993
rect 4697 2947 4703 2993
rect 5277 2966 5283 2997
rect 5427 3003 5440 3007
rect 5427 2993 5443 3003
rect 5607 3003 5620 3007
rect 5607 2993 5623 3003
rect 6847 3003 6860 3007
rect 6847 2993 6863 3003
rect 1867 2937 1933 2943
rect 3167 2937 3213 2943
rect 3847 2937 3913 2943
rect 5437 2946 5443 2993
rect 5617 2967 5623 2993
rect 6857 2967 6863 2993
rect 5607 2957 5623 2967
rect 5607 2953 5620 2957
rect 6847 2957 6863 2967
rect 6847 2953 6860 2957
rect 6467 2897 6513 2903
rect 6963 2878 7023 3382
rect 6930 2862 7023 2878
rect 1647 2837 1713 2843
rect 3087 2837 3153 2843
rect 5827 2837 5853 2843
rect 1827 2797 1893 2803
rect 2187 2797 2213 2803
rect 3907 2797 3993 2803
rect 4067 2797 4193 2803
rect 5067 2797 5153 2803
rect 6367 2797 6433 2803
rect 1497 2743 1503 2793
rect 6507 2777 6533 2783
rect 4717 2757 4753 2763
rect 4717 2747 4723 2757
rect 1497 2737 1533 2743
rect 4707 2737 4723 2747
rect 4707 2733 4720 2737
rect 6367 2737 6393 2743
rect 2747 2717 2773 2723
rect 2867 2717 2893 2723
rect 2947 2717 3013 2723
rect 5547 2717 5653 2723
rect 1267 2697 1373 2703
rect 2567 2657 2593 2663
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 6077 2583 6083 2603
rect 6027 2577 6083 2583
rect 307 2497 353 2503
rect 647 2497 793 2503
rect 1967 2497 2013 2503
rect 4407 2497 4493 2503
rect 5007 2497 5033 2503
rect 6547 2497 6653 2503
rect 1327 2477 1373 2483
rect 1467 2483 1480 2487
rect 1467 2473 1483 2483
rect 1477 2467 1483 2473
rect 4777 2477 4853 2483
rect 1477 2466 1500 2467
rect 1477 2457 1493 2466
rect 1480 2453 1493 2457
rect 1307 2417 1333 2423
rect 2387 2417 2493 2423
rect 4207 2417 4293 2423
rect 4597 2407 4603 2433
rect 4777 2383 4783 2477
rect 4957 2477 5013 2483
rect 4957 2447 4963 2477
rect 6007 2477 6093 2483
rect 6187 2477 6233 2483
rect 6367 2477 6413 2483
rect 6567 2477 6593 2483
rect 6907 2457 6933 2463
rect 4947 2437 4963 2447
rect 4947 2433 4960 2437
rect 6007 2417 6073 2423
rect 4807 2397 4873 2403
rect 4777 2377 4853 2383
rect 6963 2358 7023 2862
rect 6930 2342 7023 2358
rect 4827 2317 4873 2323
rect 4807 2277 4873 2283
rect 6407 2277 6493 2283
rect 1067 2257 1113 2263
rect 5167 2257 5213 2263
rect 6057 2257 6113 2263
rect 1387 2223 1400 2227
rect 1387 2213 1403 2223
rect 1397 2183 1403 2213
rect 1867 2217 1913 2223
rect 6057 2223 6063 2257
rect 6037 2217 6063 2223
rect 1413 2203 1427 2213
rect 1413 2200 1453 2203
rect 1417 2197 1453 2200
rect 1907 2197 1973 2203
rect 5747 2197 5793 2203
rect 6037 2203 6043 2217
rect 6007 2197 6043 2203
rect 6207 2197 6273 2203
rect 6287 2197 6353 2203
rect 1397 2177 1433 2183
rect 2387 2177 2413 2183
rect 4987 2157 5013 2163
rect 5027 2137 5053 2143
rect 5507 2117 5573 2123
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 5817 2043 5823 2083
rect 5847 2057 5893 2063
rect 5817 2037 5873 2043
rect 5127 2017 5193 2023
rect 6407 2017 6453 2023
rect 6587 2017 6613 2023
rect 1747 1997 1813 2003
rect 6027 1997 6053 2003
rect 1427 1977 1513 1983
rect 4607 1977 4653 1983
rect 4967 1977 5073 1983
rect 5887 1977 5933 1983
rect 5987 1977 6033 1983
rect 4687 1957 4713 1963
rect 4987 1957 5043 1963
rect 5037 1927 5043 1957
rect 6587 1957 6653 1963
rect 2567 1917 2633 1923
rect 5037 1917 5053 1927
rect 5040 1913 5053 1917
rect 87 1897 133 1903
rect 1307 1897 1353 1903
rect 2867 1897 2933 1903
rect 1767 1877 1853 1883
rect 6427 1877 6473 1883
rect 1927 1857 1973 1863
rect 6963 1838 7023 2342
rect 6930 1822 7023 1838
rect 3847 1777 3873 1783
rect 3727 1757 3793 1763
rect 6177 1757 6213 1763
rect 1087 1737 1133 1743
rect 1567 1737 1633 1743
rect 5927 1737 6013 1743
rect 6177 1707 6183 1757
rect 6787 1757 6843 1763
rect 6660 1743 6673 1747
rect 6657 1733 6673 1743
rect 6657 1707 6663 1733
rect 6837 1707 6843 1757
rect 927 1697 973 1703
rect 6177 1697 6193 1707
rect 6180 1693 6193 1697
rect 6657 1697 6673 1707
rect 6660 1693 6673 1697
rect 6837 1697 6853 1707
rect 6840 1693 6853 1697
rect 1547 1677 1573 1683
rect 6407 1677 6493 1683
rect 6587 1677 6633 1683
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 947 1477 1033 1483
rect 527 1457 573 1463
rect 6347 1457 6393 1463
rect 827 1443 840 1447
rect 827 1433 843 1443
rect 2347 1443 2360 1447
rect 2347 1433 2363 1443
rect 837 1407 843 1433
rect 827 1397 843 1407
rect 2357 1403 2363 1433
rect 2357 1397 2413 1403
rect 827 1393 840 1397
rect 327 1377 353 1383
rect 5647 1377 5693 1383
rect 6963 1318 7023 1822
rect 6930 1302 7023 1318
rect 6647 1237 6693 1243
rect 2407 1223 2420 1227
rect 2407 1213 2423 1223
rect 2907 1223 2920 1227
rect 2907 1213 2923 1223
rect 2417 1187 2423 1213
rect 2407 1177 2423 1187
rect 2917 1183 2923 1213
rect 2917 1177 2973 1183
rect 2407 1173 2420 1177
rect 5967 1177 6013 1183
rect 827 1157 873 1163
rect 887 1157 913 1163
rect 967 1157 1033 1163
rect 1187 1157 1253 1163
rect 1987 1157 2053 1163
rect 2527 1157 2553 1163
rect 2567 1157 2653 1163
rect 2747 1157 2813 1163
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 4207 977 4233 983
rect 4447 957 4473 963
rect 4527 957 4593 963
rect 6307 957 6353 963
rect 187 937 313 943
rect 3447 937 3473 943
rect 4547 937 4613 943
rect 5527 937 5593 943
rect 727 917 773 923
rect 6307 917 6373 923
rect 1607 857 1673 863
rect 3847 857 3893 863
rect 3907 857 3933 863
rect 4407 857 4473 863
rect 1367 837 1393 843
rect 2607 837 2653 843
rect 6963 798 7023 1302
rect 6930 782 7023 798
rect 567 637 653 643
rect 1747 637 1793 643
rect 3427 637 3573 643
rect 4027 637 4093 643
rect 4607 637 4693 643
rect -63 522 30 538
rect -63 18 -3 522
rect 2487 477 2533 483
rect 627 417 673 423
rect 1947 417 2053 423
rect 2707 417 2733 423
rect 4487 417 4513 423
rect 4807 417 4913 423
rect 2167 337 2193 343
rect 2387 337 2433 343
rect 3387 297 3413 303
rect 6963 278 7023 782
rect 6930 262 7023 278
rect 6847 117 6893 123
rect 4707 97 4853 103
rect -63 2 30 18
rect 6963 2 7023 262
<< m2contact >>
rect 6493 6413 6507 6427
rect 6593 6413 6607 6427
rect 3973 6353 3987 6367
rect 4073 6353 4087 6367
rect 4933 6353 4947 6367
rect 4993 6353 5007 6367
rect 6373 6353 6387 6367
rect 6453 6353 6467 6367
rect 233 6213 247 6227
rect 533 6233 547 6247
rect 953 6233 967 6247
rect 1513 6233 1527 6247
rect 1953 6233 1967 6247
rect 5493 6153 5507 6167
rect 5613 6153 5627 6167
rect 1673 6133 1687 6147
rect 1733 6133 1747 6147
rect 2493 6133 2507 6147
rect 2593 6133 2607 6147
rect 3073 6133 3087 6147
rect 3233 6133 3247 6147
rect 4433 6133 4447 6147
rect 4513 6133 4527 6147
rect 6053 6133 6067 6147
rect 6113 6133 6127 6147
rect 5693 6113 5707 6127
rect 5733 6113 5747 6127
rect 2653 6053 2667 6067
rect 2733 6053 2747 6067
rect 3933 6053 3947 6067
rect 3973 6053 3987 6067
rect 6313 6053 6327 6067
rect 6393 6053 6407 6067
rect 4813 6033 4827 6047
rect 4873 6033 4887 6047
rect 4933 5953 4947 5967
rect 4993 5953 5007 5967
rect 4613 5933 4627 5947
rect 4693 5933 4707 5947
rect 5133 5933 5147 5947
rect 5173 5933 5187 5947
rect 3393 5912 3407 5926
rect 3453 5913 3467 5927
rect 2973 5893 2987 5907
rect 3033 5893 3047 5907
rect 3273 5893 3287 5907
rect 3333 5893 3347 5907
rect 3413 5893 3427 5907
rect 4233 5893 4247 5907
rect 4273 5893 4287 5907
rect 1553 5873 1567 5887
rect 1633 5873 1647 5887
rect 3413 5853 3427 5867
rect 4773 5853 4787 5867
rect 4833 5853 4847 5867
rect 3533 5833 3547 5847
rect 3693 5833 3707 5847
rect 3873 5833 3887 5847
rect 3933 5833 3947 5847
rect 4013 5833 4027 5847
rect 4093 5833 4107 5847
rect 4213 5833 4227 5847
rect 4333 5833 4347 5847
rect 4573 5833 4587 5847
rect 4693 5833 4707 5847
rect 5233 5833 5247 5847
rect 5272 5833 5286 5847
rect 5293 5833 5307 5847
rect 5373 5833 5387 5847
rect 5953 5833 5967 5847
rect 6053 5833 6067 5847
rect 6513 5833 6527 5847
rect 6593 5833 6607 5847
rect 6333 5813 6347 5827
rect 6453 5813 6467 5827
rect 6293 5793 6307 5807
rect 6413 5793 6427 5807
rect 5293 5773 5307 5787
rect 5333 5772 5347 5786
rect 1153 5713 1167 5727
rect 1193 5713 1207 5727
rect 1913 5633 1927 5647
rect 2073 5633 2087 5647
rect 2113 5633 2127 5647
rect 2233 5632 2247 5646
rect 2113 5612 2127 5626
rect 2193 5613 2207 5627
rect 2733 5613 2747 5627
rect 2793 5613 2807 5627
rect 4613 5613 4627 5627
rect 4673 5613 4687 5627
rect 4773 5613 4787 5627
rect 4873 5613 4887 5627
rect 6153 5613 6167 5627
rect 6213 5613 6227 5627
rect 6553 5614 6567 5628
rect 1013 5593 1027 5607
rect 3093 5593 3107 5607
rect 6453 5593 6467 5607
rect 1013 5553 1027 5567
rect 3093 5553 3107 5567
rect 4833 5553 4847 5567
rect 4893 5553 4907 5567
rect 5633 5553 5647 5567
rect 5673 5553 5687 5567
rect 5753 5553 5767 5567
rect 5793 5553 5807 5567
rect 6453 5553 6467 5567
rect 6533 5553 6547 5567
rect 3933 5533 3947 5547
rect 4013 5533 4027 5547
rect 4113 5533 4127 5547
rect 4173 5533 4187 5547
rect 4833 5532 4847 5546
rect 4993 5533 5007 5547
rect 853 5513 867 5527
rect 893 5513 907 5527
rect 3153 5433 3167 5447
rect 3193 5433 3207 5447
rect 2613 5413 2627 5427
rect 2653 5413 2667 5427
rect 3913 5393 3927 5407
rect 3993 5393 4007 5407
rect 5493 5393 5507 5407
rect 5593 5393 5607 5407
rect 5853 5393 5867 5407
rect 5933 5393 5947 5407
rect 5973 5393 5987 5407
rect 6073 5393 6087 5407
rect 6693 5393 6707 5407
rect 653 5373 667 5387
rect 5293 5373 5307 5387
rect 733 5333 747 5347
rect 1653 5333 1667 5347
rect 1693 5333 1707 5347
rect 2073 5313 2087 5327
rect 2113 5313 2127 5327
rect 4713 5313 4727 5327
rect 4793 5313 4807 5327
rect 6393 5373 6407 5387
rect 6653 5373 6667 5387
rect 6393 5333 6407 5347
rect 6653 5333 6667 5347
rect 5393 5313 5407 5327
rect 5433 5313 5447 5327
rect 5473 5313 5487 5327
rect 5573 5313 5587 5327
rect 5653 5313 5667 5327
rect 5773 5313 5787 5327
rect 5873 5313 5887 5327
rect 5933 5313 5947 5327
rect 6273 5313 6287 5327
rect 6353 5313 6367 5327
rect 6733 5373 6747 5387
rect 6833 5373 6847 5387
rect 6733 5333 6747 5347
rect 6753 5313 6767 5327
rect 6813 5313 6827 5327
rect 2353 5293 2367 5307
rect 2393 5293 2407 5307
rect 5313 5293 5327 5307
rect 6433 5293 6447 5307
rect 6533 5293 6547 5307
rect 93 5193 107 5207
rect 253 5193 267 5207
rect 1193 5193 1207 5207
rect 5773 5113 5787 5127
rect 5833 5113 5847 5127
rect 6133 5113 6147 5127
rect 1353 5093 1367 5107
rect 1393 5093 1407 5107
rect 2993 5093 3007 5107
rect 3073 5093 3087 5107
rect 3893 5093 3907 5107
rect 3933 5093 3947 5107
rect 353 5013 367 5027
rect 513 5013 527 5027
rect 613 5013 627 5027
rect 793 5013 807 5027
rect 2933 5073 2947 5087
rect 4693 5073 4707 5087
rect 4993 5073 5007 5087
rect 5653 5073 5667 5087
rect 5713 5073 5727 5087
rect 4693 5033 4707 5047
rect 5073 5033 5087 5047
rect 5453 5033 5467 5047
rect 5513 5033 5527 5047
rect 2873 5012 2887 5026
rect 3153 5011 3167 5025
rect 3193 5013 3207 5027
rect 3533 5013 3547 5027
rect 3613 5013 3627 5027
rect 6453 5093 6467 5107
rect 6513 5093 6527 5107
rect 6793 5093 6807 5107
rect 6413 5073 6427 5087
rect 6453 5053 6467 5067
rect 6413 5033 6427 5047
rect 6653 5073 6667 5087
rect 6493 5033 6507 5047
rect 6573 5033 6587 5047
rect 653 4993 667 5007
rect 773 4993 787 5007
rect 6133 4993 6147 5007
rect 6813 4992 6827 5006
rect 5053 4913 5067 4927
rect 5113 4913 5127 4927
rect 5893 4893 5907 4907
rect 5973 4893 5987 4907
rect 773 4873 787 4887
rect 893 4873 907 4887
rect 1613 4873 1627 4887
rect 1733 4873 1747 4887
rect 2113 4873 2127 4887
rect 2173 4873 2187 4887
rect 4153 4873 4167 4887
rect 4273 4874 4287 4888
rect 5893 4872 5907 4886
rect 5973 4872 5987 4886
rect 6033 4873 6047 4887
rect 6133 4873 6147 4887
rect 6393 4873 6407 4887
rect 6473 4874 6487 4888
rect 6553 4873 6567 4887
rect 6613 4873 6627 4887
rect 2553 4853 2567 4867
rect 2613 4853 2627 4867
rect 3533 4853 3547 4867
rect 3573 4853 3587 4867
rect 4453 4853 4467 4867
rect 5033 4853 5047 4867
rect 4913 4833 4927 4847
rect 5293 4853 5307 4867
rect 6273 4853 6287 4867
rect 6513 4853 6527 4867
rect 3853 4813 3867 4827
rect 3913 4813 3927 4827
rect 4373 4813 4387 4827
rect 4853 4813 4867 4827
rect 5033 4813 5047 4827
rect 5073 4813 5087 4827
rect 5113 4813 5127 4827
rect 5293 4813 5307 4827
rect 6193 4813 6207 4827
rect 6833 4853 6847 4867
rect 6893 4832 6907 4846
rect 6593 4813 6607 4827
rect 2893 4793 2907 4807
rect 2953 4793 2967 4807
rect 4333 4791 4347 4805
rect 4473 4793 4487 4807
rect 4853 4792 4867 4806
rect 4933 4793 4947 4807
rect 5353 4793 5367 4807
rect 5513 4793 5527 4807
rect 5853 4793 5867 4807
rect 5933 4793 5947 4807
rect 6013 4793 6027 4807
rect 6133 4793 6147 4807
rect 6173 4793 6187 4807
rect 6273 4793 6287 4807
rect 5053 4773 5067 4787
rect 5133 4773 5147 4787
rect 5173 4772 5187 4786
rect 5213 4773 5227 4787
rect 5293 4773 5307 4787
rect 6193 4772 6207 4786
rect 6253 4773 6267 4787
rect 2533 4753 2547 4767
rect 2613 4753 2627 4767
rect 4413 4752 4427 4766
rect 4473 4753 4487 4767
rect 5213 4733 5227 4747
rect 5273 4733 5287 4747
rect 2993 4713 3007 4727
rect 3073 4713 3087 4727
rect 4373 4713 4387 4727
rect 4453 4713 4467 4727
rect 4193 4653 4207 4667
rect 4273 4653 4287 4667
rect 4393 4653 4407 4667
rect 4433 4653 4447 4667
rect 4913 4653 4927 4667
rect 4973 4653 4987 4667
rect 4713 4613 4727 4627
rect 4793 4613 4807 4627
rect 4733 4593 4747 4607
rect 4813 4593 4827 4607
rect 5833 4593 5847 4607
rect 5973 4593 5987 4607
rect 953 4573 967 4587
rect 1113 4573 1127 4587
rect 3213 4573 3227 4587
rect 3253 4573 3267 4587
rect 4333 4573 4347 4587
rect 4433 4573 4447 4587
rect 4493 4573 4507 4587
rect 4573 4573 4587 4587
rect 4653 4573 4667 4587
rect 4813 4572 4827 4586
rect 4853 4573 4867 4587
rect 4973 4573 4987 4587
rect 5233 4573 5247 4587
rect 3013 4553 3027 4567
rect 4093 4553 4107 4567
rect 4533 4553 4547 4567
rect 3013 4513 3027 4527
rect 4013 4513 4027 4527
rect 4533 4513 4547 4527
rect 4613 4553 4627 4567
rect 4793 4553 4807 4567
rect 6053 4573 6067 4587
rect 6093 4573 6107 4587
rect 6233 4573 6247 4587
rect 5313 4553 5327 4567
rect 5633 4553 5647 4567
rect 5713 4553 5727 4567
rect 5573 4533 5587 4547
rect 4613 4513 4627 4527
rect 4793 4513 4807 4527
rect 5713 4513 5727 4527
rect 3633 4493 3647 4507
rect 3673 4493 3687 4507
rect 3713 4493 3727 4507
rect 4893 4493 4907 4507
rect 4953 4493 4967 4507
rect 5233 4493 5247 4507
rect 5353 4493 5367 4507
rect 5393 4493 5407 4507
rect 5493 4493 5507 4507
rect 5693 4493 5707 4507
rect 5793 4553 5807 4567
rect 6313 4553 6327 4567
rect 6073 4513 6087 4527
rect 6173 4513 6187 4527
rect 6313 4513 6327 4527
rect 6833 4553 6847 4567
rect 6413 4513 6427 4527
rect 6833 4513 6847 4527
rect 6213 4493 6227 4507
rect 6353 4493 6367 4507
rect 6473 4493 6487 4507
rect 6513 4493 6527 4507
rect 4893 4472 4907 4486
rect 4973 4473 4987 4487
rect 5393 4472 5407 4486
rect 5453 4473 5467 4487
rect 5713 4473 5727 4487
rect 5793 4473 5807 4487
rect 6513 4472 6527 4486
rect 6593 4473 6607 4487
rect 1013 4453 1027 4467
rect 1053 4453 1067 4467
rect 5713 4373 5727 4387
rect 5873 4373 5887 4387
rect 5913 4373 5927 4387
rect 2073 4353 2087 4367
rect 2173 4353 2187 4367
rect 2813 4353 2827 4367
rect 2873 4354 2887 4368
rect 5473 4353 5487 4367
rect 5553 4353 5567 4367
rect 5633 4353 5647 4367
rect 5793 4353 5807 4367
rect 1933 4333 1947 4347
rect 1973 4333 1987 4347
rect 2313 4333 2327 4347
rect 2373 4333 2387 4347
rect 4973 4332 4987 4346
rect 5013 4333 5027 4347
rect 5413 4333 5427 4347
rect 5493 4333 5507 4347
rect 5673 4333 5687 4347
rect 6113 4353 6127 4367
rect 6153 4353 6167 4367
rect 6213 4353 6227 4367
rect 5333 4293 5347 4307
rect 5573 4293 5587 4307
rect 5673 4293 5687 4307
rect 5933 4293 5947 4307
rect 6013 4293 6027 4307
rect 6173 4293 6187 4307
rect 6213 4293 6227 4307
rect 6433 4353 6447 4367
rect 6413 4333 6427 4347
rect 6493 4333 6507 4347
rect 6533 4333 6547 4347
rect 1513 4271 1527 4285
rect 1693 4273 1707 4287
rect 4633 4273 4647 4287
rect 4673 4273 4687 4287
rect 4713 4273 4727 4287
rect 4833 4271 4847 4285
rect 4913 4273 4927 4287
rect 5053 4273 5067 4287
rect 5113 4273 5127 4287
rect 5233 4271 5247 4285
rect 5793 4273 5807 4287
rect 5893 4273 5907 4287
rect 6153 4273 6167 4287
rect 6273 4273 6287 4287
rect 6533 4312 6547 4326
rect 6573 4293 6587 4307
rect 6653 4293 6667 4307
rect 6713 4293 6727 4307
rect 4753 4253 4767 4267
rect 4813 4253 4827 4267
rect 6173 4253 6187 4267
rect 6353 4272 6367 4286
rect 6413 4273 6427 4287
rect 6473 4273 6487 4287
rect 6593 4273 6607 4287
rect 6273 4252 6287 4266
rect 6313 4252 6327 4266
rect 5993 4233 6007 4247
rect 6073 4233 6087 4247
rect 5853 4213 5867 4227
rect 5893 4213 5907 4227
rect 5133 4192 5147 4206
rect 5213 4193 5227 4207
rect 813 4153 827 4167
rect 2753 4073 2767 4087
rect 2813 4073 2827 4087
rect 6113 4073 6127 4087
rect 6233 4073 6247 4087
rect 6753 4073 6767 4087
rect 6833 4073 6847 4087
rect 213 4053 227 4067
rect 273 4054 287 4068
rect 1033 4053 1047 4067
rect 1133 4053 1147 4067
rect 1533 4053 1547 4067
rect 1593 4053 1607 4067
rect 1713 4053 1727 4067
rect 1793 4054 1807 4068
rect 2673 4053 2687 4067
rect 2833 4053 2847 4067
rect 3493 4053 3507 4067
rect 3613 4052 3627 4066
rect 4713 4053 4727 4067
rect 4753 4053 4767 4067
rect 2353 4033 2367 4047
rect 2393 4033 2407 4047
rect 4533 4033 4547 4047
rect 4553 4013 4567 4027
rect 4853 4053 4867 4067
rect 6413 4053 6427 4067
rect 6513 4053 6527 4067
rect 6573 4053 6587 4067
rect 6633 4053 6647 4067
rect 5373 4033 5387 4047
rect 5613 4033 5627 4047
rect 5813 4033 5827 4047
rect 5853 4033 5867 4047
rect 6293 4033 6307 4047
rect 4533 3993 4547 4007
rect 173 3973 187 3987
rect 213 3973 227 3987
rect 1453 3973 1467 3987
rect 1573 3973 1587 3987
rect 4313 3973 4327 3987
rect 4353 3972 4367 3986
rect 4513 3973 4527 3987
rect 4593 3973 4607 3987
rect 4753 3993 4767 4007
rect 4813 3993 4827 4007
rect 5373 3993 5387 4007
rect 5493 3993 5507 4007
rect 5533 3993 5547 4007
rect 5613 3993 5627 4007
rect 6593 4033 6607 4047
rect 6653 4033 6667 4047
rect 6373 3993 6387 4007
rect 4613 3953 4627 3967
rect 4753 3972 4767 3986
rect 4853 3971 4867 3985
rect 5093 3973 5107 3987
rect 5193 3973 5207 3987
rect 5433 3973 5447 3987
rect 5553 3973 5567 3987
rect 5593 3973 5607 3987
rect 5673 3973 5687 3987
rect 6773 3973 6787 3987
rect 6873 3973 6887 3987
rect 6933 3973 6947 3987
rect 4813 3953 4827 3967
rect 5113 3953 5127 3967
rect 5153 3953 5167 3967
rect 6733 3953 6747 3967
rect 5453 3933 5467 3947
rect 5533 3933 5547 3947
rect 5633 3932 5647 3946
rect 5693 3933 5707 3947
rect 893 3833 907 3847
rect 953 3833 967 3847
rect 2573 3833 2587 3847
rect 2613 3833 2627 3847
rect 3053 3833 3067 3847
rect 3153 3833 3167 3847
rect 3313 3833 3327 3847
rect 3393 3834 3407 3848
rect 3433 3833 3447 3847
rect 3553 3833 3567 3847
rect 6173 3833 6187 3847
rect 2153 3813 2167 3827
rect 2213 3813 2227 3827
rect 5593 3813 5607 3827
rect 5653 3813 5667 3827
rect 5933 3813 5947 3827
rect 4393 3793 4407 3807
rect 3113 3773 3127 3787
rect 3153 3773 3167 3787
rect 673 3753 687 3767
rect 793 3753 807 3767
rect 1593 3753 1607 3767
rect 1733 3753 1747 3767
rect 2033 3753 2047 3767
rect 2113 3753 2127 3767
rect 2913 3753 2927 3767
rect 2993 3753 3007 3767
rect 3053 3753 3067 3767
rect 3173 3753 3187 3767
rect 5953 3792 5967 3806
rect 6113 3773 6127 3787
rect 6193 3813 6207 3827
rect 6553 3813 6567 3827
rect 6633 3813 6647 3827
rect 6193 3773 6207 3787
rect 6473 3773 6487 3787
rect 6713 3773 6727 3787
rect 4373 3752 4387 3766
rect 5693 3753 5707 3767
rect 5853 3753 5867 3767
rect 5953 3753 5967 3767
rect 6033 3753 6047 3767
rect 6073 3753 6087 3767
rect 5393 3732 5407 3746
rect 5433 3733 5447 3747
rect 6153 3753 6167 3767
rect 6233 3753 6247 3767
rect 6213 3732 6227 3746
rect 6413 3733 6427 3747
rect 6513 3733 6527 3747
rect 1833 3673 1847 3687
rect 1893 3673 1907 3687
rect 4533 3673 4547 3687
rect 4613 3673 4627 3687
rect 6633 3673 6647 3687
rect 6673 3673 6687 3687
rect 653 3633 667 3647
rect 1193 3633 1207 3647
rect 4053 3633 4067 3647
rect 4293 3633 4307 3647
rect 4813 3633 4827 3647
rect 5893 3633 5907 3647
rect 1293 3613 1307 3627
rect 1353 3613 1367 3627
rect 1813 3593 1827 3607
rect 1873 3593 1887 3607
rect 4613 3593 4627 3607
rect 4693 3592 4707 3606
rect 6073 3593 6087 3607
rect 6113 3593 6127 3607
rect 6573 3573 6587 3587
rect 6613 3573 6627 3587
rect 2133 3553 2147 3567
rect 2253 3553 2267 3567
rect 2753 3553 2767 3567
rect 2793 3553 2807 3567
rect 5913 3553 5927 3567
rect 6013 3553 6027 3567
rect 6453 3553 6467 3567
rect 6493 3553 6507 3567
rect 6713 3553 6727 3567
rect 6873 3553 6887 3567
rect 593 3533 607 3547
rect 753 3533 767 3547
rect 3333 3533 3347 3547
rect 3413 3533 3427 3547
rect 4453 3533 4467 3547
rect 4513 3533 4527 3547
rect 4573 3533 4587 3547
rect 4633 3533 4647 3547
rect 4793 3532 4807 3546
rect 4893 3533 4907 3547
rect 5573 3533 5587 3547
rect 1193 3513 1207 3527
rect 1453 3513 1467 3527
rect 1513 3513 1527 3527
rect 4433 3513 4447 3527
rect 1193 3473 1207 3487
rect 2033 3473 2047 3487
rect 2073 3473 2087 3487
rect 3193 3473 3207 3487
rect 3233 3473 3247 3487
rect 4513 3473 4527 3487
rect 5213 3473 5227 3487
rect 5293 3473 5307 3487
rect 5393 3473 5407 3487
rect 5453 3473 5467 3487
rect 3133 3453 3147 3467
rect 3213 3452 3227 3466
rect 5193 3453 5207 3467
rect 5313 3453 5327 3467
rect 5533 3453 5547 3467
rect 5653 3533 5667 3547
rect 6213 3533 6227 3547
rect 6333 3534 6347 3548
rect 6533 3534 6547 3548
rect 6573 3533 6587 3547
rect 6653 3533 6667 3547
rect 6713 3532 6727 3546
rect 6133 3513 6147 3527
rect 6493 3513 6507 3527
rect 5633 3473 5647 3487
rect 6133 3473 6147 3487
rect 6233 3473 6247 3487
rect 6313 3473 6327 3487
rect 6493 3473 6507 3487
rect 6773 3473 6787 3487
rect 6853 3473 6867 3487
rect 5593 3413 5607 3427
rect 5633 3413 5647 3427
rect 6553 3353 6567 3367
rect 6613 3353 6627 3367
rect 1253 3333 1267 3347
rect 1293 3333 1307 3347
rect 1693 3333 1707 3347
rect 1773 3332 1787 3346
rect 6413 3333 6427 3347
rect 1113 3313 1127 3327
rect 1153 3313 1167 3327
rect 1313 3314 1327 3328
rect 3133 3313 3147 3327
rect 3253 3312 3267 3326
rect 4053 3313 4067 3327
rect 4093 3313 4107 3327
rect 5473 3313 5487 3327
rect 5573 3312 5587 3326
rect 6473 3312 6487 3326
rect 33 3293 47 3307
rect 93 3293 107 3307
rect 1193 3293 1207 3307
rect 1293 3293 1307 3307
rect 1673 3293 1687 3307
rect 1733 3293 1747 3307
rect 2153 3293 2167 3307
rect 2233 3293 2247 3307
rect 5452 3293 5466 3307
rect 5473 3292 5487 3306
rect 5553 3293 5567 3307
rect 6373 3293 6387 3307
rect 6413 3293 6427 3307
rect 6453 3293 6467 3307
rect 5553 3253 5567 3267
rect 6453 3253 6467 3267
rect 753 3233 767 3247
rect 813 3233 827 3247
rect 1133 3233 1147 3247
rect 1233 3233 1247 3247
rect 1493 3233 1507 3247
rect 1533 3233 1547 3247
rect 3353 3233 3367 3247
rect 3453 3233 3467 3247
rect 5673 3233 5687 3247
rect 5713 3233 5727 3247
rect 6233 3233 6247 3247
rect 6273 3233 6287 3247
rect 3973 3113 3987 3127
rect 5273 3113 5287 3127
rect 6833 3073 6847 3087
rect 6913 3073 6927 3087
rect 5393 3053 5407 3067
rect 5473 3053 5487 3067
rect 2493 3033 2507 3047
rect 2533 3033 2547 3047
rect 2133 3013 2147 3027
rect 2173 3013 2187 3027
rect 2813 3013 2827 3027
rect 2853 3013 2867 3027
rect 3013 3013 3027 3027
rect 3073 3013 3087 3027
rect 3313 3013 3327 3027
rect 3393 3013 3407 3027
rect 4313 3013 4327 3027
rect 4393 3013 4407 3027
rect 6793 3013 6807 3027
rect 6913 3013 6927 3027
rect 4553 2993 4567 3007
rect 4713 2993 4727 3007
rect 4533 2973 4547 2987
rect 5353 2993 5367 3007
rect 5413 2993 5427 3007
rect 5593 2993 5607 3007
rect 6833 2993 6847 3007
rect 5273 2952 5287 2966
rect 1853 2933 1867 2947
rect 1933 2933 1947 2947
rect 3153 2933 3167 2947
rect 3213 2933 3227 2947
rect 3833 2933 3847 2947
rect 3913 2931 3927 2945
rect 4693 2933 4707 2947
rect 5593 2953 5607 2967
rect 6833 2953 6847 2967
rect 5433 2932 5447 2946
rect 6453 2893 6467 2907
rect 6513 2893 6527 2907
rect 1633 2833 1647 2847
rect 1713 2833 1727 2847
rect 3073 2833 3087 2847
rect 3153 2833 3167 2847
rect 5813 2833 5827 2847
rect 5853 2833 5867 2847
rect 1493 2793 1507 2807
rect 1813 2793 1827 2807
rect 1893 2793 1907 2807
rect 2173 2793 2187 2807
rect 2213 2793 2227 2807
rect 3893 2793 3907 2807
rect 3993 2793 4007 2807
rect 4053 2793 4067 2807
rect 4193 2793 4207 2807
rect 5053 2793 5067 2807
rect 5153 2793 5167 2807
rect 6353 2793 6367 2807
rect 6433 2793 6447 2807
rect 6493 2773 6507 2787
rect 6533 2773 6547 2787
rect 4753 2753 4767 2767
rect 1533 2733 1547 2747
rect 4693 2733 4707 2747
rect 6353 2733 6367 2747
rect 6393 2733 6407 2747
rect 2733 2713 2747 2727
rect 2773 2713 2787 2727
rect 2853 2713 2867 2727
rect 2893 2711 2907 2725
rect 2933 2711 2947 2725
rect 3013 2713 3027 2727
rect 5533 2713 5547 2727
rect 5653 2713 5667 2727
rect 1253 2693 1267 2707
rect 1373 2693 1387 2707
rect 2553 2653 2567 2667
rect 2593 2653 2607 2667
rect 353 2593 367 2607
rect 673 2593 687 2607
rect 6013 2573 6027 2587
rect 293 2493 307 2507
rect 353 2493 367 2507
rect 633 2493 647 2507
rect 793 2493 807 2507
rect 1953 2493 1967 2507
rect 2013 2493 2027 2507
rect 4393 2493 4407 2507
rect 4493 2493 4507 2507
rect 4993 2493 5007 2507
rect 5033 2493 5047 2507
rect 6533 2493 6547 2507
rect 6653 2493 6667 2507
rect 1313 2473 1327 2487
rect 1373 2473 1387 2487
rect 1453 2473 1467 2487
rect 1493 2452 1507 2466
rect 4593 2433 4607 2447
rect 1293 2413 1307 2427
rect 1333 2413 1347 2427
rect 2373 2413 2387 2427
rect 2493 2413 2507 2427
rect 4193 2411 4207 2425
rect 4293 2413 4307 2427
rect 4593 2393 4607 2407
rect 4853 2473 4867 2487
rect 5013 2473 5027 2487
rect 5993 2473 6007 2487
rect 6093 2473 6107 2487
rect 6173 2473 6187 2487
rect 6233 2473 6247 2487
rect 6353 2473 6367 2487
rect 6413 2473 6427 2487
rect 6553 2473 6567 2487
rect 6593 2473 6607 2487
rect 6893 2453 6907 2467
rect 6933 2453 6947 2467
rect 4933 2433 4947 2447
rect 5993 2413 6007 2427
rect 6073 2413 6087 2427
rect 4793 2393 4807 2407
rect 4873 2393 4887 2407
rect 4853 2373 4867 2387
rect 4813 2313 4827 2327
rect 4873 2313 4887 2327
rect 4793 2273 4807 2287
rect 4873 2273 4887 2287
rect 6393 2273 6407 2287
rect 6493 2273 6507 2287
rect 1053 2253 1067 2267
rect 1113 2253 1127 2267
rect 5153 2253 5167 2267
rect 5213 2253 5227 2267
rect 1373 2213 1387 2227
rect 1413 2213 1427 2227
rect 1853 2213 1867 2227
rect 1913 2213 1927 2227
rect 6113 2253 6127 2267
rect 1453 2193 1467 2207
rect 1893 2193 1907 2207
rect 1973 2191 1987 2205
rect 5733 2193 5747 2207
rect 5793 2193 5807 2207
rect 5993 2193 6007 2207
rect 6193 2193 6207 2207
rect 6273 2193 6287 2207
rect 6353 2193 6367 2207
rect 1433 2173 1447 2187
rect 2373 2173 2387 2187
rect 2413 2173 2427 2187
rect 4973 2153 4987 2167
rect 5013 2153 5027 2167
rect 5013 2132 5027 2146
rect 5053 2133 5067 2147
rect 5493 2113 5507 2127
rect 5573 2113 5587 2127
rect 93 2073 107 2087
rect 2573 2073 2587 2087
rect 2833 2073 2847 2087
rect 2893 2073 2907 2087
rect 3913 2073 3927 2087
rect 5833 2053 5847 2067
rect 5893 2053 5907 2067
rect 5873 2033 5887 2047
rect 5113 2013 5127 2027
rect 5193 2013 5207 2027
rect 6393 2013 6407 2027
rect 6453 2013 6467 2027
rect 6573 2013 6587 2027
rect 6613 2012 6627 2026
rect 1733 1993 1747 2007
rect 1813 1993 1827 2007
rect 6013 1993 6027 2007
rect 6053 1993 6067 2007
rect 1413 1973 1427 1987
rect 1513 1973 1527 1987
rect 4593 1974 4607 1988
rect 4653 1973 4667 1987
rect 4953 1973 4967 1987
rect 5073 1973 5087 1987
rect 5873 1973 5887 1987
rect 5933 1973 5947 1987
rect 5973 1973 5987 1987
rect 6033 1973 6047 1987
rect 4673 1953 4687 1967
rect 4713 1953 4727 1967
rect 4973 1953 4987 1967
rect 6573 1953 6587 1967
rect 6653 1953 6667 1967
rect 2553 1913 2567 1927
rect 2633 1913 2647 1927
rect 5053 1913 5067 1927
rect 73 1893 87 1907
rect 133 1893 147 1907
rect 1293 1893 1307 1907
rect 1353 1893 1367 1907
rect 2853 1893 2867 1907
rect 2933 1893 2947 1907
rect 1753 1873 1767 1887
rect 1853 1873 1867 1887
rect 6413 1873 6427 1887
rect 6473 1873 6487 1887
rect 1913 1853 1927 1867
rect 1973 1853 1987 1867
rect 3833 1773 3847 1787
rect 3873 1773 3887 1787
rect 3713 1753 3727 1767
rect 3793 1753 3807 1767
rect 1073 1733 1087 1747
rect 1133 1733 1147 1747
rect 1553 1733 1567 1747
rect 1633 1733 1647 1747
rect 5913 1733 5927 1747
rect 6013 1733 6027 1747
rect 6213 1753 6227 1767
rect 6773 1753 6787 1767
rect 6673 1733 6687 1747
rect 913 1693 927 1707
rect 973 1693 987 1707
rect 6193 1693 6207 1707
rect 6673 1693 6687 1707
rect 6853 1693 6867 1707
rect 1533 1671 1547 1685
rect 1573 1673 1587 1687
rect 6393 1673 6407 1687
rect 6493 1673 6507 1687
rect 6573 1673 6587 1687
rect 6633 1673 6647 1687
rect 2953 1553 2967 1567
rect 2973 1553 2987 1567
rect 3153 1553 3167 1567
rect 3353 1553 3367 1567
rect 4893 1553 4907 1567
rect 5593 1553 5607 1567
rect 5653 1553 5667 1567
rect 933 1473 947 1487
rect 1033 1473 1047 1487
rect 513 1453 527 1467
rect 573 1454 587 1468
rect 6333 1454 6347 1468
rect 6393 1453 6407 1467
rect 813 1433 827 1447
rect 2333 1433 2347 1447
rect 813 1393 827 1407
rect 2413 1393 2427 1407
rect 313 1373 327 1387
rect 353 1373 367 1387
rect 5633 1373 5647 1387
rect 5693 1373 5707 1387
rect 6633 1233 6647 1247
rect 6693 1233 6707 1247
rect 2393 1213 2407 1227
rect 2893 1213 2907 1227
rect 2393 1173 2407 1187
rect 2973 1173 2987 1187
rect 5953 1173 5967 1187
rect 6013 1173 6027 1187
rect 813 1153 827 1167
rect 873 1153 887 1167
rect 913 1153 927 1167
rect 953 1153 967 1167
rect 1033 1153 1047 1167
rect 1173 1153 1187 1167
rect 1253 1153 1267 1167
rect 1973 1153 1987 1167
rect 2053 1153 2067 1167
rect 2513 1153 2527 1167
rect 2553 1153 2567 1167
rect 2653 1153 2667 1167
rect 2733 1153 2747 1167
rect 2813 1153 2827 1167
rect 2353 1033 2367 1047
rect 3113 1033 3127 1047
rect 5573 1033 5587 1047
rect 5833 1033 5847 1047
rect 6093 1033 6107 1047
rect 4193 973 4207 987
rect 4233 973 4247 987
rect 4433 953 4447 967
rect 4473 953 4487 967
rect 4513 953 4527 967
rect 4593 953 4607 967
rect 6293 953 6307 967
rect 6353 953 6367 967
rect 173 933 187 947
rect 313 933 327 947
rect 3433 933 3447 947
rect 3473 933 3487 947
rect 4533 933 4547 947
rect 4613 933 4627 947
rect 5513 933 5527 947
rect 5593 933 5607 947
rect 713 913 727 927
rect 773 913 787 927
rect 6293 913 6307 927
rect 6373 913 6387 927
rect 1593 853 1607 867
rect 1673 853 1687 867
rect 3833 853 3847 867
rect 3893 853 3907 867
rect 3933 853 3947 867
rect 4393 853 4407 867
rect 4473 853 4487 867
rect 1353 833 1367 847
rect 1393 833 1407 847
rect 2593 833 2607 847
rect 2653 833 2667 847
rect 553 633 567 647
rect 653 633 667 647
rect 1733 633 1747 647
rect 1793 633 1807 647
rect 3413 633 3427 647
rect 3573 633 3587 647
rect 4013 633 4027 647
rect 4093 633 4107 647
rect 4593 633 4607 647
rect 4693 633 4707 647
rect 2013 513 2027 527
rect 2193 513 2207 527
rect 5073 513 5087 527
rect 6453 513 6467 527
rect 2473 473 2487 487
rect 2533 473 2547 487
rect 613 413 627 427
rect 673 413 687 427
rect 1933 413 1947 427
rect 2053 413 2067 427
rect 2693 413 2707 427
rect 2733 413 2747 427
rect 4473 413 4487 427
rect 4513 413 4527 427
rect 4793 413 4807 427
rect 4913 413 4927 427
rect 2153 331 2167 345
rect 2193 333 2207 347
rect 2373 333 2387 347
rect 2433 333 2447 347
rect 3373 292 3387 306
rect 3413 293 3427 307
rect 6833 113 6847 127
rect 6893 113 6907 127
rect 4693 93 4707 107
rect 4853 93 4867 107
<< metal2 >>
rect 296 6527 303 6563
rect 336 6383 343 6513
rect 436 6447 443 6563
rect 476 6556 503 6563
rect 427 6416 443 6423
rect 316 6376 343 6383
rect 16 6086 23 6113
rect 16 5367 23 6072
rect 236 5876 243 6213
rect 356 6116 363 6313
rect 256 6086 263 6114
rect 256 5908 263 6072
rect 416 6067 423 6414
rect 496 6407 503 6556
rect 2987 6456 3013 6463
rect 6467 6456 6503 6463
rect 556 6396 583 6403
rect 476 6116 483 6333
rect 516 6247 523 6363
rect 576 6327 583 6396
rect 576 6287 583 6313
rect 676 6247 683 6403
rect 516 6236 533 6247
rect 520 6233 533 6236
rect 536 6083 543 6114
rect 716 6087 723 6233
rect 816 6227 823 6413
rect 856 6396 883 6403
rect 913 6400 927 6413
rect 916 6396 923 6400
rect 876 6347 883 6396
rect 833 6120 847 6133
rect 836 6116 843 6120
rect 516 6076 543 6083
rect 116 5860 123 5863
rect 113 5846 127 5860
rect 196 5727 203 5832
rect 56 5367 63 5713
rect 196 5616 203 5713
rect 156 5507 163 5563
rect 236 5467 243 5583
rect 256 5487 263 5894
rect 356 5787 363 5883
rect 356 5576 363 5613
rect 496 5503 503 6053
rect 536 5883 543 5973
rect 536 5876 563 5883
rect 556 5583 563 5876
rect 536 5576 563 5583
rect 496 5496 513 5503
rect 76 5356 103 5363
rect 16 5287 23 5313
rect 16 3927 23 4293
rect 36 3548 43 4673
rect 56 3727 63 5273
rect 96 5207 103 5356
rect 196 5307 203 5363
rect 336 5207 343 5453
rect 396 5287 403 5473
rect 436 5356 463 5363
rect 176 5023 183 5074
rect 156 5016 183 5023
rect 156 4856 163 5016
rect 76 4307 83 4753
rect 196 4576 203 4673
rect 236 4607 243 4993
rect 256 4543 263 5193
rect 356 5076 363 5113
rect 336 5007 343 5043
rect 316 4687 323 4823
rect 236 4536 263 4543
rect 336 4543 343 4593
rect 356 4567 363 5013
rect 396 5007 403 5043
rect 436 4868 443 5273
rect 456 5167 463 5356
rect 476 5307 483 5413
rect 476 4787 483 4823
rect 496 4807 503 5354
rect 516 5027 523 5493
rect 636 5487 643 6083
rect 676 5867 683 6083
rect 856 5967 863 6083
rect 896 6007 903 6133
rect 916 5987 923 6333
rect 936 6247 943 6393
rect 976 6287 983 6363
rect 936 6236 953 6247
rect 940 6233 953 6236
rect 936 6128 943 6213
rect 976 6207 983 6273
rect 1016 6116 1023 6153
rect 1076 6136 1083 6193
rect 1136 6147 1143 6403
rect 1316 6396 1333 6403
rect 1373 6400 1387 6413
rect 1376 6396 1383 6400
rect 1476 6396 1503 6403
rect 1336 6347 1343 6394
rect 936 6047 943 6114
rect 1036 6047 1043 6083
rect 536 5346 543 5393
rect 596 5376 603 5413
rect 640 5383 653 5387
rect 636 5376 653 5383
rect 640 5373 653 5376
rect 616 5076 623 5113
rect 676 5083 683 5773
rect 796 5627 803 5863
rect 753 5600 767 5613
rect 756 5596 763 5600
rect 736 5527 743 5563
rect 736 5383 743 5513
rect 776 5447 783 5552
rect 716 5376 743 5383
rect 816 5403 823 5853
rect 916 5608 923 5863
rect 956 5687 963 5863
rect 996 5827 1003 6033
rect 1036 5787 1043 6033
rect 1056 6007 1063 6053
rect 1076 5967 1083 5993
rect 1096 5896 1103 6033
rect 1116 5967 1123 6103
rect 1236 6096 1243 6173
rect 1376 6047 1383 6333
rect 1436 6287 1443 6363
rect 1436 6227 1443 6273
rect 1496 6247 1503 6396
rect 1596 6283 1603 6403
rect 1576 6276 1603 6283
rect 1496 6236 1513 6247
rect 1500 6233 1513 6236
rect 1416 6047 1423 6103
rect 1176 5956 1193 5963
rect 1176 5876 1183 5956
rect 1096 5787 1103 5813
rect 836 5566 843 5593
rect 753 5380 767 5393
rect 796 5396 823 5403
rect 796 5388 803 5396
rect 756 5376 763 5380
rect 696 5346 703 5373
rect 696 5147 703 5332
rect 676 5076 703 5083
rect 696 5046 703 5076
rect 596 5023 603 5043
rect 596 5016 613 5023
rect 616 4856 623 5013
rect 596 4767 603 4823
rect 636 4820 663 4823
rect 636 4816 667 4820
rect 653 4807 667 4816
rect 336 4536 363 4543
rect 176 4003 183 4093
rect 156 3996 183 4003
rect 176 3816 183 3973
rect 196 3967 203 4334
rect 216 4107 223 4512
rect 236 4407 243 4493
rect 256 4447 263 4536
rect 316 4336 323 4393
rect 216 3987 223 4053
rect 236 4007 243 4253
rect 256 4047 263 4292
rect 336 4267 343 4303
rect 287 4056 323 4063
rect 376 4056 383 4433
rect 496 4347 503 4593
rect 536 4527 543 4543
rect 536 4307 543 4513
rect 436 4067 443 4253
rect 536 4207 543 4293
rect 556 4287 563 4653
rect 596 4487 603 4543
rect 616 4527 623 4793
rect 636 4347 643 4773
rect 656 4526 663 4793
rect 696 4727 703 5032
rect 716 5027 723 5376
rect 776 5227 783 5343
rect 856 5343 863 5433
rect 876 5367 883 5493
rect 936 5447 943 5552
rect 976 5387 983 5713
rect 996 5567 1003 5613
rect 1016 5607 1023 5633
rect 1096 5596 1103 5773
rect 1136 5727 1143 5843
rect 1196 5727 1203 5953
rect 1156 5647 1163 5713
rect 1016 5363 1023 5553
rect 1036 5427 1043 5552
rect 1053 5463 1067 5473
rect 1076 5463 1083 5563
rect 1156 5487 1163 5594
rect 1176 5566 1183 5693
rect 1296 5607 1303 5883
rect 1436 5827 1443 6133
rect 1476 5967 1483 6033
rect 1476 5876 1483 5953
rect 1236 5527 1243 5563
rect 1316 5547 1323 5773
rect 1496 5747 1503 6153
rect 1516 6087 1523 6173
rect 1576 5987 1583 6276
rect 1736 6207 1743 6413
rect 1836 6396 1863 6403
rect 1936 6396 1963 6403
rect 1856 6287 1863 6396
rect 1633 6120 1647 6133
rect 1673 6120 1687 6133
rect 1636 6116 1643 6120
rect 1676 6116 1683 6120
rect 1616 6007 1623 6083
rect 1716 6027 1723 6133
rect 1736 6087 1743 6133
rect 1796 6128 1803 6253
rect 1896 6227 1903 6363
rect 1956 6247 1963 6396
rect 2047 6403 2060 6407
rect 2047 6396 2063 6403
rect 2236 6396 2263 6403
rect 2296 6396 2323 6403
rect 2047 6393 2060 6396
rect 1836 6116 1843 6153
rect 1996 6116 2003 6153
rect 2033 6120 2047 6133
rect 2036 6116 2043 6120
rect 1616 5908 1623 5993
rect 1676 5908 1683 5933
rect 1716 5896 1723 5973
rect 1540 5883 1553 5887
rect 1536 5876 1553 5883
rect 1540 5873 1553 5876
rect 1616 5867 1623 5894
rect 1856 5896 1863 6072
rect 1416 5596 1423 5633
rect 1336 5566 1343 5593
rect 1053 5460 1083 5463
rect 1056 5456 1083 5460
rect 1036 5387 1043 5413
rect 1016 5356 1043 5363
rect 856 5336 923 5343
rect 816 5207 823 5332
rect 736 5003 743 5093
rect 716 4996 743 5003
rect 716 4807 723 4996
rect 756 4927 763 5074
rect 796 5040 803 5043
rect 793 5027 807 5040
rect 876 4903 883 5133
rect 896 5127 903 5313
rect 956 5287 963 5343
rect 896 5046 903 5113
rect 856 4896 883 4903
rect 773 4860 787 4873
rect 776 4856 783 4860
rect 756 4820 763 4823
rect 753 4807 767 4820
rect 836 4487 843 4854
rect 856 4587 863 4896
rect 916 4887 923 5213
rect 1016 5103 1023 5293
rect 1056 5287 1063 5456
rect 1136 5307 1143 5353
rect 933 5083 947 5093
rect 996 5096 1023 5103
rect 933 5080 963 5083
rect 936 5076 963 5080
rect 996 5076 1003 5096
rect 1056 5046 1063 5233
rect 1156 5207 1163 5363
rect 1296 5247 1303 5473
rect 1336 5363 1343 5493
rect 1396 5427 1403 5563
rect 1436 5560 1443 5563
rect 1433 5547 1447 5560
rect 1447 5536 1463 5543
rect 1336 5356 1363 5363
rect 1396 5356 1423 5363
rect 1076 5087 1083 5193
rect 976 5007 983 5043
rect 893 4868 907 4873
rect 976 4767 983 4854
rect 916 4607 923 4753
rect 856 4526 863 4573
rect 916 4556 923 4593
rect 953 4560 967 4573
rect 956 4556 963 4560
rect 896 4520 903 4523
rect 893 4507 907 4520
rect 936 4423 943 4512
rect 996 4447 1003 5013
rect 1016 4743 1023 4953
rect 1076 4883 1083 5073
rect 1096 5047 1103 5153
rect 1056 4876 1083 4883
rect 1056 4856 1063 4876
rect 1136 4867 1143 5032
rect 1196 4836 1203 5193
rect 1236 5007 1243 5193
rect 1356 5107 1363 5356
rect 1293 5080 1307 5093
rect 1296 5076 1303 5080
rect 1376 5047 1383 5074
rect 1276 4967 1283 5043
rect 1316 5007 1323 5043
rect 1396 4967 1403 5093
rect 1416 5087 1423 5356
rect 1436 5107 1443 5373
rect 1456 5207 1463 5536
rect 1496 5247 1503 5733
rect 1636 5707 1643 5873
rect 1776 5866 1783 5893
rect 1976 5867 1983 6072
rect 1636 5566 1643 5693
rect 1536 5447 1543 5533
rect 1556 5487 1563 5513
rect 1576 5376 1583 5453
rect 1496 5076 1503 5233
rect 1556 5127 1563 5343
rect 1596 5340 1603 5343
rect 1593 5327 1607 5340
rect 1636 5167 1643 5552
rect 1656 5347 1663 5853
rect 1696 5627 1703 5863
rect 1876 5747 1883 5863
rect 1916 5727 1923 5863
rect 1776 5596 1783 5653
rect 1676 5388 1683 5594
rect 1816 5566 1823 5673
rect 1716 5527 1723 5563
rect 1836 5543 1843 5594
rect 1856 5567 1863 5613
rect 1956 5596 1963 5753
rect 1996 5563 2003 5953
rect 2096 5908 2103 6273
rect 2196 6207 2203 6273
rect 2216 6116 2223 6213
rect 2156 6027 2163 6083
rect 2196 6063 2203 6083
rect 2196 6056 2223 6063
rect 2216 5896 2223 6056
rect 2256 5967 2263 6396
rect 2316 6327 2323 6396
rect 2276 6128 2283 6153
rect 1976 5556 2003 5563
rect 1816 5536 1843 5543
rect 1676 5323 1683 5374
rect 1716 5340 1723 5343
rect 1656 5316 1683 5323
rect 1656 5076 1663 5316
rect 1696 5083 1703 5333
rect 1713 5327 1727 5340
rect 1696 5076 1713 5083
rect 1556 5047 1563 5074
rect 1016 4736 1043 4743
rect 1016 4467 1023 4554
rect 1036 4527 1043 4736
rect 1076 4727 1083 4823
rect 1096 4587 1103 4793
rect 1116 4707 1123 4823
rect 1156 4800 1163 4803
rect 1153 4787 1167 4800
rect 1113 4560 1127 4573
rect 1116 4556 1123 4560
rect 1176 4527 1183 4793
rect 936 4416 963 4423
rect 576 4267 583 4333
rect 696 4316 723 4323
rect 816 4320 823 4323
rect 596 4300 603 4303
rect 593 4287 607 4300
rect 656 4280 663 4283
rect 653 4267 667 4280
rect 716 4167 723 4316
rect 813 4307 827 4320
rect 316 4036 323 4056
rect 436 4023 443 4053
rect 416 4016 443 4023
rect 336 3847 343 4003
rect 356 3816 363 3953
rect 396 3887 403 4013
rect 116 3647 123 3783
rect 76 3500 83 3503
rect 73 3487 87 3500
rect 96 3307 103 3533
rect 176 3503 183 3553
rect 196 3527 203 3772
rect 256 3767 263 3814
rect 176 3496 203 3503
rect 36 3028 43 3293
rect 136 3260 143 3263
rect 133 3247 147 3260
rect 176 3207 183 3294
rect 256 3127 263 3263
rect 336 3247 343 3751
rect 356 3567 363 3713
rect 356 3223 363 3493
rect 376 3347 383 3503
rect 396 3447 403 3833
rect 416 3687 423 3913
rect 436 3647 443 3973
rect 676 3927 683 4014
rect 476 3816 483 3913
rect 436 3447 443 3503
rect 456 3487 463 3613
rect 476 3427 483 3633
rect 496 3607 503 3783
rect 416 3296 423 3373
rect 396 3260 403 3263
rect 393 3247 407 3260
rect 336 3216 363 3223
rect 56 2976 83 2983
rect 56 2847 63 2976
rect 76 2707 83 2953
rect 96 2827 103 3013
rect 196 2976 203 3113
rect 336 2967 343 3216
rect 436 3127 443 3263
rect 376 2927 383 2983
rect 116 2667 123 2713
rect 136 2707 143 2743
rect 196 2707 203 2813
rect 116 2476 123 2513
rect 136 2407 143 2443
rect 176 2407 183 2653
rect 196 2347 203 2693
rect 216 2647 223 2774
rect 236 2667 243 2833
rect 396 2767 403 3053
rect 476 3047 483 3333
rect 496 3187 503 3553
rect 416 2976 443 2983
rect 416 2847 423 2976
rect 416 2756 423 2793
rect 256 2527 263 2733
rect 276 2476 283 2713
rect 296 2627 303 2743
rect 436 2727 443 2953
rect 476 2927 483 3033
rect 516 2967 523 3633
rect 536 3487 543 3913
rect 616 3816 623 3873
rect 636 3767 643 3783
rect 676 3780 683 3783
rect 673 3767 687 3780
rect 596 3547 603 3593
rect 596 3516 603 3533
rect 636 3528 643 3753
rect 716 3747 723 3814
rect 736 3766 743 4053
rect 776 3987 783 4023
rect 796 3947 803 4113
rect 653 3627 667 3633
rect 756 3607 763 3933
rect 816 3923 823 4073
rect 796 3916 823 3923
rect 796 3828 803 3916
rect 836 3816 843 4133
rect 856 4026 863 4193
rect 856 3927 863 4012
rect 776 3707 783 3773
rect 816 3767 823 3783
rect 807 3756 823 3767
rect 807 3753 820 3756
rect 856 3747 863 3773
rect 676 3487 683 3573
rect 616 3463 623 3483
rect 596 3456 623 3463
rect 596 3308 603 3456
rect 656 3266 663 3373
rect 616 3260 623 3263
rect 613 3247 627 3260
rect 696 3247 703 3593
rect 753 3547 767 3553
rect 756 3480 763 3483
rect 753 3467 767 3480
rect 756 3427 763 3453
rect 836 3447 843 3593
rect 836 3267 843 3294
rect 756 3260 763 3263
rect 753 3247 767 3260
rect 776 3067 783 3233
rect 796 3223 803 3263
rect 856 3243 863 3653
rect 876 3567 883 4173
rect 956 4127 963 4416
rect 1016 4147 1023 4453
rect 1056 4328 1063 4453
rect 1076 4227 1083 4493
rect 1096 4203 1103 4512
rect 1136 4487 1143 4523
rect 1196 4487 1203 4593
rect 1216 4527 1223 4913
rect 1456 4846 1463 4893
rect 1476 4868 1483 4933
rect 1496 4836 1503 4953
rect 1516 4947 1523 5043
rect 1516 4727 1523 4933
rect 1556 4836 1563 4973
rect 1636 4903 1643 5032
rect 1676 4987 1683 5043
rect 1636 4896 1663 4903
rect 1253 4560 1267 4573
rect 1256 4556 1263 4560
rect 1296 4556 1303 4593
rect 1416 4556 1423 4693
rect 1076 4196 1103 4203
rect 1116 4476 1133 4483
rect 916 4036 923 4113
rect 956 4036 963 4073
rect 1076 4067 1083 4196
rect 1116 4087 1123 4476
rect 1156 4348 1163 4433
rect 1276 4387 1283 4523
rect 1196 4336 1203 4373
rect 1156 4167 1163 4334
rect 1316 4303 1323 4513
rect 1316 4296 1343 4303
rect 1376 4300 1383 4303
rect 1036 4007 1043 4053
rect 1133 4040 1147 4053
rect 1136 4036 1143 4040
rect 976 3887 983 4003
rect 1056 3887 1063 4034
rect 896 3607 903 3833
rect 916 3727 923 3833
rect 953 3820 967 3833
rect 993 3820 1007 3833
rect 1076 3828 1083 3933
rect 1116 3907 1123 4003
rect 1156 3947 1163 4003
rect 1196 3907 1203 4073
rect 1216 3967 1223 4213
rect 1293 4040 1307 4053
rect 1296 4036 1303 4040
rect 1276 4000 1283 4003
rect 1273 3987 1287 4000
rect 1336 3987 1343 4296
rect 1373 4287 1387 4300
rect 1416 4247 1423 4334
rect 1436 4328 1443 4523
rect 1476 4347 1483 4553
rect 1576 4487 1583 4523
rect 1496 4336 1503 4373
rect 1436 4207 1443 4314
rect 1500 4285 1520 4287
rect 1507 4273 1513 4285
rect 1556 4227 1563 4303
rect 1576 4247 1583 4293
rect 1596 4127 1603 4373
rect 1356 4007 1363 4093
rect 1616 4087 1623 4873
rect 1656 4767 1663 4896
rect 1716 4868 1723 5074
rect 1736 4887 1743 5293
rect 1756 5047 1763 5332
rect 1816 5127 1823 5536
rect 1876 5376 1883 5453
rect 1896 5336 1923 5343
rect 1916 5267 1923 5336
rect 1856 5076 1863 5113
rect 1756 4856 1763 4893
rect 1796 4826 1803 5043
rect 1836 5023 1843 5043
rect 1816 5016 1843 5023
rect 1696 4820 1703 4823
rect 1693 4807 1707 4820
rect 1816 4807 1823 5016
rect 1916 4987 1923 5253
rect 1916 4887 1923 4973
rect 1956 4927 1963 5374
rect 1976 5343 1983 5556
rect 2016 5388 2023 5853
rect 2096 5727 2103 5894
rect 2116 5867 2123 5894
rect 2116 5687 2123 5853
rect 2136 5827 2143 5873
rect 2116 5663 2123 5673
rect 2116 5656 2143 5663
rect 2087 5636 2113 5643
rect 2056 5607 2063 5633
rect 2113 5600 2127 5612
rect 2136 5608 2143 5656
rect 2116 5596 2123 5600
rect 2056 5376 2063 5513
rect 1976 5336 2003 5343
rect 1873 4860 1887 4873
rect 1876 4856 1883 4860
rect 1836 4568 1843 4853
rect 1896 4820 1903 4823
rect 1893 4807 1907 4820
rect 1896 4647 1903 4693
rect 1976 4563 1983 5193
rect 1996 5076 2003 5336
rect 2036 5247 2043 5343
rect 2076 5340 2083 5343
rect 2073 5327 2087 5340
rect 2116 5327 2123 5493
rect 2136 5467 2143 5553
rect 2156 5347 2163 5713
rect 2176 5527 2183 5813
rect 2196 5627 2203 5863
rect 2236 5707 2243 5863
rect 2236 5667 2243 5693
rect 2276 5647 2283 6114
rect 2296 6087 2303 6173
rect 2316 6147 2323 6313
rect 2396 5923 2403 6433
rect 2493 6420 2507 6433
rect 2496 6416 2503 6420
rect 2416 6376 2443 6383
rect 2476 6380 2483 6383
rect 2416 6187 2423 6376
rect 2473 6367 2487 6380
rect 2536 6367 2543 6413
rect 2716 6386 2723 6453
rect 2993 6428 3007 6433
rect 3156 6416 3163 6453
rect 2436 6207 2443 6253
rect 2436 6086 2443 6193
rect 2676 6167 2683 6383
rect 2776 6376 2803 6383
rect 2776 6347 2783 6376
rect 2493 6120 2507 6133
rect 2496 6116 2503 6120
rect 2536 6116 2543 6153
rect 2576 6086 2583 6113
rect 2476 6047 2483 6083
rect 2467 6036 2483 6047
rect 2467 6033 2480 6036
rect 2596 6027 2603 6133
rect 2716 6116 2723 6153
rect 2776 6116 2783 6333
rect 2836 6327 2843 6372
rect 2396 5916 2413 5923
rect 2413 5900 2427 5913
rect 2416 5896 2423 5900
rect 2576 5896 2583 5933
rect 2456 5866 2463 5893
rect 2356 5827 2363 5863
rect 2296 5727 2303 5773
rect 2376 5767 2383 5793
rect 2240 5646 2260 5647
rect 2247 5643 2260 5646
rect 2247 5633 2263 5643
rect 2256 5623 2263 5633
rect 2256 5616 2283 5623
rect 2196 5567 2203 5613
rect 2276 5608 2283 5616
rect 2196 5487 2203 5532
rect 2196 5376 2203 5473
rect 2256 5383 2263 5563
rect 2356 5487 2363 5573
rect 2376 5467 2383 5753
rect 2496 5566 2503 5733
rect 2416 5560 2423 5563
rect 2413 5547 2427 5560
rect 2416 5507 2423 5533
rect 2456 5487 2463 5563
rect 2516 5547 2523 5813
rect 2556 5627 2563 5863
rect 2636 5827 2643 5993
rect 2656 5807 2663 6053
rect 2676 5908 2683 6072
rect 2733 6067 2747 6072
rect 2756 5896 2763 5933
rect 2796 5903 2803 6153
rect 2816 6007 2823 6253
rect 2796 5896 2823 5903
rect 2576 5596 2583 5733
rect 2636 5727 2643 5773
rect 2636 5566 2643 5713
rect 2676 5707 2683 5894
rect 2816 5866 2823 5896
rect 2736 5807 2743 5863
rect 2836 5827 2843 6313
rect 2876 6127 2883 6413
rect 3236 6387 3243 6414
rect 2976 6347 2983 6383
rect 2996 6047 3003 6313
rect 2896 5896 2903 6013
rect 2936 5896 2943 6033
rect 3016 6027 3023 6383
rect 3136 6327 3143 6383
rect 3176 6363 3183 6383
rect 3176 6356 3203 6363
rect 3073 6128 3087 6133
rect 3116 6128 3123 6193
rect 2967 5893 2973 5907
rect 2976 5866 2983 5893
rect 2876 5747 2883 5863
rect 3016 5787 3023 6013
rect 3056 5923 3063 6083
rect 3036 5920 3063 5923
rect 3033 5916 3063 5920
rect 3033 5907 3047 5916
rect 3076 5896 3083 6013
rect 2236 5376 2263 5383
rect 2073 5307 2087 5313
rect 2216 5127 2223 5343
rect 2096 5076 2123 5083
rect 2016 4787 2023 4823
rect 2056 4667 2063 4823
rect 2096 4707 2103 5076
rect 2116 4667 2123 4873
rect 2173 4860 2187 4873
rect 2176 4856 2183 4860
rect 1976 4556 2003 4563
rect 1836 4526 1843 4554
rect 1816 4487 1823 4512
rect 1956 4487 1963 4523
rect 1636 4067 1643 4353
rect 1776 4306 1783 4473
rect 1896 4360 1943 4363
rect 1896 4356 1947 4360
rect 1896 4336 1903 4356
rect 1933 4347 1947 4356
rect 1696 4300 1703 4303
rect 1693 4287 1707 4300
rect 1607 4063 1620 4067
rect 1607 4053 1623 4063
rect 1433 4040 1447 4053
rect 1436 4036 1443 4040
rect 1456 4000 1463 4003
rect 1453 3987 1467 4000
rect 1096 3896 1113 3903
rect 956 3816 963 3820
rect 996 3816 1003 3820
rect 1096 3587 1103 3896
rect 1336 3807 1343 3973
rect 1176 3743 1183 3793
rect 1376 3796 1383 3913
rect 1176 3736 1203 3743
rect 1196 3647 1203 3736
rect 1293 3627 1307 3633
rect 1356 3627 1363 3673
rect 1396 3607 1403 3813
rect 1436 3796 1463 3803
rect 1456 3727 1463 3796
rect 1476 3747 1483 3953
rect 916 3516 923 3553
rect 936 3427 943 3483
rect 996 3407 1003 3514
rect 836 3236 863 3243
rect 796 3220 823 3223
rect 793 3216 823 3220
rect 793 3207 807 3216
rect 776 2996 783 3053
rect 676 2823 683 2993
rect 676 2816 703 2823
rect 376 2720 383 2723
rect 373 2707 387 2720
rect 296 2507 303 2613
rect 356 2607 363 2653
rect 316 2476 323 2513
rect 356 2446 363 2493
rect 256 2347 263 2443
rect 56 2247 63 2333
rect 76 2236 103 2243
rect 196 2240 203 2243
rect 96 2087 103 2236
rect 193 2227 207 2240
rect 376 2236 383 2273
rect 256 1927 263 1954
rect 396 1927 403 2713
rect 676 2607 683 2793
rect 696 2766 703 2816
rect 716 2763 723 2913
rect 756 2907 763 2963
rect 716 2756 743 2763
rect 773 2760 787 2773
rect 776 2756 783 2760
rect 736 2603 743 2756
rect 716 2596 743 2603
rect 456 2476 463 2593
rect 620 2503 633 2507
rect 616 2493 633 2503
rect 616 2476 623 2493
rect 436 2407 443 2443
rect 436 2236 443 2393
rect 476 2347 483 2443
rect 476 2127 483 2333
rect 136 1920 143 1923
rect 76 1407 83 1893
rect 96 1787 103 1913
rect 133 1907 147 1920
rect 156 1776 163 1893
rect 256 1867 263 1913
rect 276 1607 283 1692
rect 296 1647 303 1893
rect 316 1807 323 1923
rect 156 1436 163 1513
rect 136 1216 143 1273
rect 116 1180 123 1183
rect 113 1167 127 1180
rect 176 947 183 1213
rect 196 1167 203 1553
rect 216 1287 223 1434
rect 196 967 203 1153
rect 176 916 183 933
rect 216 928 223 1273
rect 236 1227 243 1473
rect 276 1436 283 1593
rect 336 1487 343 1703
rect 336 1443 343 1473
rect 316 1436 343 1443
rect 296 1267 303 1403
rect 356 1387 363 1633
rect 396 1407 403 1793
rect 416 1748 423 2093
rect 496 2047 503 2433
rect 536 2407 543 2473
rect 547 2396 563 2403
rect 436 1706 443 2033
rect 516 1956 523 1993
rect 496 1736 503 1773
rect 436 1567 443 1692
rect 516 1547 523 1703
rect 436 1436 443 1513
rect 516 1507 523 1533
rect 476 1443 483 1493
rect 476 1436 503 1443
rect 256 1216 263 1253
rect 316 1243 323 1373
rect 456 1307 463 1403
rect 496 1307 503 1436
rect 296 1236 323 1243
rect 296 1216 303 1236
rect 356 1186 363 1213
rect 396 1186 403 1273
rect 276 1147 283 1183
rect 516 1047 523 1453
rect 556 1443 563 2396
rect 636 2187 643 2443
rect 676 2226 683 2513
rect 696 2447 703 2573
rect 716 2283 723 2596
rect 796 2547 803 2952
rect 816 2847 823 3216
rect 836 2527 843 3236
rect 916 2996 923 3252
rect 953 3247 967 3252
rect 996 3127 1003 3293
rect 893 2947 907 2952
rect 856 2647 863 2774
rect 793 2480 807 2493
rect 796 2476 803 2480
rect 776 2440 783 2443
rect 773 2427 787 2440
rect 756 2416 773 2423
rect 716 2276 733 2283
rect 736 2223 743 2273
rect 716 2216 743 2223
rect 576 1468 583 2113
rect 676 1956 683 1993
rect 716 1956 723 2153
rect 756 2107 763 2416
rect 596 1867 603 1954
rect 656 1867 663 1923
rect 696 1736 703 1873
rect 636 1527 643 1703
rect 676 1627 683 1703
rect 536 1436 563 1443
rect 536 1247 543 1436
rect 616 1436 623 1473
rect 227 916 243 923
rect 96 703 103 753
rect 116 727 123 883
rect 156 807 163 883
rect 153 708 167 713
rect 96 696 123 703
rect 196 627 203 872
rect 236 767 243 916
rect 313 920 327 933
rect 316 916 323 920
rect 516 916 523 953
rect 536 947 543 1233
rect 556 1187 563 1293
rect 636 1287 643 1403
rect 696 1327 703 1434
rect 596 1216 603 1273
rect 676 1186 683 1214
rect 616 1147 623 1183
rect 276 887 283 914
rect 436 887 443 914
rect 116 396 123 533
rect 216 487 223 694
rect 236 547 243 753
rect 336 696 343 872
rect 456 696 463 793
rect 496 696 503 883
rect 536 807 543 883
rect 276 623 283 663
rect 556 647 563 693
rect 256 616 283 623
rect 156 396 163 473
rect 256 367 263 616
rect 276 396 283 493
rect 336 396 363 403
rect 456 396 463 493
rect 296 360 303 363
rect 293 347 307 360
rect 156 176 163 213
rect 316 176 323 213
rect 356 146 363 396
rect 556 367 563 413
rect 476 360 483 363
rect 473 347 487 360
rect 576 347 583 933
rect 616 847 623 1112
rect 676 987 683 1172
rect 716 1127 723 1693
rect 736 1607 743 1734
rect 756 1707 763 1954
rect 776 1887 783 2353
rect 856 2347 863 2633
rect 876 2427 883 2833
rect 936 2827 943 2963
rect 976 2827 983 2994
rect 996 2907 1003 3113
rect 1016 2963 1023 3453
rect 1076 3447 1083 3483
rect 1076 3323 1083 3433
rect 1156 3327 1163 3573
rect 1207 3523 1220 3527
rect 1207 3516 1223 3523
rect 1207 3513 1220 3516
rect 1176 3327 1183 3513
rect 1196 3347 1203 3473
rect 1236 3407 1243 3483
rect 1296 3347 1303 3592
rect 1396 3516 1403 3572
rect 1456 3527 1463 3713
rect 1336 3467 1343 3514
rect 1056 3316 1083 3323
rect 1056 3207 1063 3316
rect 1113 3300 1127 3313
rect 1180 3303 1193 3307
rect 1116 3296 1123 3300
rect 1176 3296 1193 3303
rect 1180 3293 1193 3296
rect 1136 3260 1143 3263
rect 1133 3247 1147 3260
rect 1236 3247 1243 3293
rect 1016 2956 1043 2963
rect 976 2747 983 2813
rect 996 2587 1003 2774
rect 956 2476 963 2553
rect 936 2407 943 2443
rect 1016 2427 1023 2913
rect 1036 2783 1043 2956
rect 1116 2960 1123 2963
rect 1113 2947 1127 2960
rect 1036 2776 1053 2783
rect 1096 2776 1103 2833
rect 1136 2627 1143 2953
rect 1156 2503 1163 3053
rect 1176 3008 1183 3193
rect 1256 3027 1263 3333
rect 1316 3328 1323 3353
rect 1307 3293 1313 3307
rect 1356 3296 1363 3353
rect 1376 3307 1383 3472
rect 1416 3427 1423 3483
rect 1476 3407 1483 3693
rect 1496 3487 1503 3873
rect 1516 3727 1523 4034
rect 1536 3527 1543 4053
rect 1616 4036 1623 4053
rect 1556 4006 1563 4033
rect 1556 3947 1563 3992
rect 1576 3828 1583 3973
rect 1636 3843 1643 3873
rect 1616 3836 1643 3843
rect 1616 3816 1623 3836
rect 1676 3786 1683 4113
rect 1596 3780 1603 3783
rect 1556 3516 1563 3773
rect 1593 3767 1607 3780
rect 1636 3687 1643 3783
rect 1593 3520 1607 3533
rect 1596 3516 1603 3520
rect 1516 3363 1523 3513
rect 1516 3356 1533 3363
rect 1276 3167 1283 3273
rect 1336 3167 1343 3263
rect 1496 3247 1503 3263
rect 1276 2996 1283 3153
rect 1176 2827 1183 2994
rect 1176 2743 1183 2813
rect 1236 2776 1243 2873
rect 1176 2736 1203 2743
rect 1136 2496 1163 2503
rect 1136 2476 1143 2496
rect 1056 2443 1063 2474
rect 1056 2436 1083 2443
rect 856 2256 863 2333
rect 916 2167 923 2313
rect 936 2227 943 2254
rect 796 1926 803 2053
rect 856 1827 863 1923
rect 896 1907 903 1923
rect 776 1547 783 1753
rect 796 1567 803 1734
rect 816 1527 823 1703
rect 800 1443 813 1447
rect 796 1436 813 1443
rect 800 1433 813 1436
rect 836 1407 843 1473
rect 816 1367 823 1393
rect 776 1216 783 1353
rect 700 923 713 927
rect 696 916 713 923
rect 700 913 713 916
rect 736 863 743 1153
rect 756 887 763 1183
rect 796 1047 803 1183
rect 856 1167 863 1633
rect 876 1627 883 1703
rect 896 1647 903 1893
rect 916 1707 923 1853
rect 876 1367 883 1513
rect 896 1447 903 1573
rect 936 1487 943 2213
rect 956 1707 963 2413
rect 1040 2263 1053 2267
rect 1036 2256 1053 2263
rect 1040 2253 1053 2256
rect 1076 2227 1083 2436
rect 1116 2407 1123 2443
rect 1196 2407 1203 2736
rect 1216 2607 1223 2743
rect 1236 2563 1243 2653
rect 1256 2567 1263 2693
rect 1216 2556 1243 2563
rect 1156 2268 1163 2393
rect 1216 2307 1223 2556
rect 1276 2476 1283 2693
rect 1316 2487 1323 3013
rect 1236 2446 1243 2473
rect 1296 2427 1303 2443
rect 1336 2427 1343 3113
rect 1396 2963 1403 3173
rect 1416 3067 1423 3153
rect 1496 3127 1503 3233
rect 1396 2956 1423 2963
rect 1396 2776 1403 2853
rect 1436 2776 1443 2833
rect 1456 2787 1463 2893
rect 1376 2707 1383 2743
rect 1376 2527 1383 2593
rect 1416 2476 1423 2533
rect 1456 2487 1463 2733
rect 1036 1956 1043 2013
rect 1096 2003 1103 2253
rect 1116 2227 1123 2253
rect 1127 2216 1143 2223
rect 1096 1996 1123 2003
rect 1016 1847 1023 1923
rect 1056 1920 1063 1923
rect 1053 1907 1067 1920
rect 993 1740 1007 1753
rect 996 1736 1003 1740
rect 976 1467 983 1693
rect 1076 1567 1083 1733
rect 1096 1543 1103 1734
rect 1076 1536 1103 1543
rect 996 1443 1003 1533
rect 976 1436 1003 1443
rect 1016 1403 1023 1434
rect 956 1367 963 1403
rect 996 1396 1023 1403
rect 876 1167 883 1353
rect 936 1216 943 1313
rect 916 1180 923 1183
rect 956 1180 963 1183
rect 913 1167 927 1180
rect 953 1167 967 1180
rect 776 887 783 913
rect 736 856 763 863
rect 636 696 643 733
rect 676 696 683 833
rect 656 660 663 663
rect 616 427 623 652
rect 653 647 667 660
rect 633 400 647 413
rect 673 400 687 413
rect 636 396 643 400
rect 676 396 683 400
rect 436 176 443 213
rect 556 147 563 193
rect 596 176 603 393
rect 656 327 663 363
rect 736 307 743 733
rect 756 367 763 856
rect 796 847 803 973
rect 816 916 823 1153
rect 887 916 903 923
rect 896 887 903 916
rect 836 747 843 872
rect 936 867 943 1133
rect 856 736 863 853
rect 776 366 783 453
rect 856 360 863 363
rect 853 347 867 360
rect 636 176 643 293
rect 276 -17 283 143
rect 476 -17 483 143
rect 696 146 703 173
rect 736 146 743 193
rect 756 143 763 313
rect 916 146 923 453
rect 936 447 943 694
rect 956 467 963 1153
rect 996 1147 1003 1396
rect 1036 1167 1043 1473
rect 1056 1406 1063 1473
rect 1076 1447 1083 1536
rect 1116 1527 1123 1996
rect 1136 1747 1143 2216
rect 1216 2107 1223 2293
rect 1296 2268 1303 2413
rect 1336 2256 1343 2293
rect 1256 2223 1263 2254
rect 1376 2227 1383 2473
rect 1436 2263 1443 2443
rect 1476 2327 1483 2933
rect 1496 2807 1503 2994
rect 1496 2487 1503 2772
rect 1496 2387 1503 2452
rect 1416 2256 1443 2263
rect 1476 2256 1483 2313
rect 1516 2287 1523 3253
rect 1536 3247 1543 3353
rect 1536 2787 1543 3073
rect 1556 2807 1563 3393
rect 1576 3308 1583 3483
rect 1616 3327 1623 3483
rect 1676 3307 1683 3513
rect 1696 3347 1703 4193
rect 1716 4006 1723 4053
rect 1756 4036 1763 4113
rect 1796 4068 1803 4333
rect 1956 4306 1963 4373
rect 1876 4300 1883 4303
rect 1873 4287 1887 4300
rect 1776 3816 1783 3992
rect 1816 3907 1823 4003
rect 1813 3820 1827 3833
rect 1816 3816 1823 3820
rect 1736 3647 1743 3753
rect 1856 3687 1863 3833
rect 1876 3828 1883 4034
rect 1716 3547 1723 3613
rect 1756 3516 1763 3573
rect 1816 3487 1823 3593
rect 1736 3447 1743 3483
rect 1776 3367 1783 3483
rect 1696 3266 1703 3312
rect 1776 3308 1783 3332
rect 1816 3296 1823 3393
rect 1836 3303 1843 3673
rect 1876 3607 1883 3814
rect 1896 3687 1903 4073
rect 1976 4048 1983 4333
rect 1996 4087 2003 4556
rect 2136 4556 2143 4853
rect 2236 4823 2243 5173
rect 2316 5103 2323 5413
rect 2416 5376 2423 5453
rect 2456 5427 2463 5473
rect 2356 5307 2363 5343
rect 2396 5323 2403 5332
rect 2396 5316 2423 5323
rect 2356 5267 2363 5293
rect 2316 5096 2343 5103
rect 2253 5080 2267 5093
rect 2256 5076 2263 5080
rect 2296 4967 2303 5043
rect 2336 4907 2343 5096
rect 2356 4987 2363 5074
rect 2376 5046 2383 5093
rect 2216 4816 2243 4823
rect 2156 4567 2163 4613
rect 2076 4407 2083 4523
rect 2073 4340 2087 4353
rect 2076 4336 2083 4340
rect 2056 4300 2063 4303
rect 2053 4287 2067 4300
rect 1956 4000 1963 4003
rect 1953 3987 1967 4000
rect 1856 3327 1863 3533
rect 1893 3520 1907 3533
rect 1896 3516 1903 3520
rect 1936 3516 1943 3713
rect 1976 3516 1983 3653
rect 1996 3547 2003 4003
rect 2036 3767 2043 4033
rect 2076 4006 2083 4233
rect 2136 4036 2143 4393
rect 2176 4367 2183 4653
rect 2216 4563 2223 4816
rect 2256 4747 2263 4854
rect 2207 4556 2223 4563
rect 2236 4736 2253 4743
rect 2196 4387 2203 4553
rect 2236 4526 2243 4736
rect 2276 4587 2283 4893
rect 2356 4856 2363 4933
rect 2396 4867 2403 5293
rect 2416 5247 2423 5316
rect 2436 5267 2443 5313
rect 2456 5076 2463 5332
rect 2496 5187 2503 5393
rect 2553 5380 2567 5393
rect 2593 5380 2607 5393
rect 2616 5387 2623 5413
rect 2556 5376 2563 5380
rect 2596 5376 2603 5380
rect 2433 5027 2447 5032
rect 2376 4787 2383 4812
rect 2316 4556 2323 4613
rect 2336 4526 2343 4693
rect 2176 4306 2183 4353
rect 2236 4348 2243 4413
rect 2256 4287 2263 4303
rect 2267 4276 2283 4283
rect 2276 4223 2283 4276
rect 2296 4247 2303 4293
rect 2316 4223 2323 4333
rect 2276 4216 2323 4223
rect 2176 4167 2183 4213
rect 2176 4036 2183 4153
rect 2116 3987 2123 4003
rect 2116 3843 2123 3973
rect 2216 3887 2223 4173
rect 2316 4036 2323 4093
rect 2356 4047 2363 4573
rect 2416 4563 2423 4873
rect 2436 4826 2443 4853
rect 2456 4707 2463 4953
rect 2536 4887 2543 5153
rect 2636 5147 2643 5493
rect 2656 5427 2663 5633
rect 2676 5507 2683 5653
rect 2916 5623 2923 5733
rect 2956 5647 2963 5673
rect 3056 5667 3063 5852
rect 2896 5616 2923 5623
rect 2733 5608 2747 5613
rect 2716 5447 2723 5563
rect 2796 5507 2803 5613
rect 2896 5596 2903 5616
rect 2656 5346 2663 5392
rect 2676 5287 2683 5433
rect 2736 5376 2743 5413
rect 2816 5347 2823 5594
rect 2876 5560 2883 5563
rect 2873 5547 2887 5560
rect 2756 5327 2763 5343
rect 2556 4867 2563 5133
rect 2576 5116 2593 5123
rect 2576 5046 2583 5116
rect 2596 5076 2603 5113
rect 2616 5040 2623 5043
rect 2613 5027 2627 5040
rect 2496 4767 2503 4823
rect 2536 4820 2543 4823
rect 2533 4807 2547 4820
rect 2396 4556 2423 4563
rect 2376 4347 2383 4553
rect 2396 4348 2403 4556
rect 2436 4336 2443 4433
rect 2516 4363 2523 4613
rect 2536 4447 2543 4753
rect 2576 4563 2583 4973
rect 2596 4947 2603 4993
rect 2676 4967 2683 5233
rect 2696 4863 2703 5293
rect 2756 5287 2763 5313
rect 2676 4856 2703 4863
rect 2596 4747 2603 4853
rect 2616 4767 2623 4853
rect 2556 4556 2583 4563
rect 2616 4556 2623 4693
rect 2656 4587 2663 4823
rect 2676 4747 2683 4793
rect 2660 4563 2673 4567
rect 2656 4556 2673 4563
rect 2556 4526 2563 4556
rect 2660 4553 2673 4556
rect 2496 4356 2523 4363
rect 2416 4048 2423 4303
rect 2496 4187 2503 4356
rect 2536 4347 2543 4393
rect 2516 4147 2523 4333
rect 2636 4167 2643 4523
rect 2513 4040 2527 4053
rect 2516 4036 2523 4040
rect 2396 4006 2403 4033
rect 2536 4006 2543 4093
rect 2296 3947 2303 4003
rect 2096 3836 2123 3843
rect 2096 3816 2103 3836
rect 2140 3823 2153 3827
rect 2136 3816 2153 3823
rect 2140 3813 2153 3816
rect 2416 3816 2423 3893
rect 2456 3816 2463 3853
rect 2067 3783 2080 3787
rect 2067 3776 2083 3783
rect 2116 3780 2123 3783
rect 2067 3773 2080 3776
rect 2113 3767 2127 3780
rect 2036 3487 2043 3732
rect 2176 3667 2183 3793
rect 2216 3786 2223 3813
rect 2356 3786 2363 3813
rect 2133 3567 2147 3573
rect 2156 3516 2203 3523
rect 1836 3296 1863 3303
rect 1656 3207 1663 3263
rect 1596 2823 1603 2963
rect 1636 2847 1643 2963
rect 1587 2816 1603 2823
rect 1576 2776 1583 2813
rect 1616 2776 1623 2833
rect 1536 2487 1543 2733
rect 1556 2667 1563 2732
rect 1656 2607 1663 2853
rect 1676 2747 1683 2953
rect 1696 2847 1703 3252
rect 1736 3227 1743 3293
rect 1716 3008 1723 3133
rect 1756 3007 1763 3253
rect 1796 3027 1803 3193
rect 1856 3187 1863 3296
rect 1876 3207 1883 3473
rect 1916 3303 1923 3483
rect 1956 3427 1963 3483
rect 1896 3296 1923 3303
rect 1896 3027 1903 3296
rect 1973 3300 1987 3313
rect 1976 3296 1983 3300
rect 1956 3227 1963 3263
rect 1716 2947 1723 2994
rect 1793 3000 1807 3013
rect 1796 2996 1803 3000
rect 1956 2996 1963 3192
rect 1996 3187 2003 3263
rect 2036 3023 2043 3313
rect 2016 3016 2043 3023
rect 1776 2887 1783 2952
rect 1816 2867 1823 2963
rect 1713 2847 1727 2853
rect 1696 2707 1703 2812
rect 1736 2776 1743 2813
rect 1556 2567 1563 2593
rect 1676 2547 1683 2633
rect 1573 2480 1587 2493
rect 1576 2476 1583 2480
rect 1556 2440 1563 2443
rect 1536 2307 1543 2433
rect 1553 2427 1567 2440
rect 1556 2283 1563 2373
rect 1536 2276 1563 2283
rect 1536 2263 1543 2276
rect 1516 2256 1543 2263
rect 1416 2227 1423 2256
rect 1596 2263 1603 2443
rect 1636 2343 1643 2433
rect 1656 2367 1663 2453
rect 1676 2427 1683 2474
rect 1636 2336 1663 2343
rect 1576 2256 1603 2263
rect 1256 2216 1283 2223
rect 1176 1736 1183 1873
rect 1216 1867 1223 1923
rect 1276 1767 1283 2216
rect 1316 2147 1323 2223
rect 1447 2223 1460 2227
rect 1447 2216 1463 2223
rect 1447 2213 1460 2216
rect 1296 1747 1303 1893
rect 1316 1887 1323 2093
rect 1413 1967 1427 1973
rect 1356 1920 1363 1923
rect 1353 1907 1367 1920
rect 1316 1876 1333 1887
rect 1320 1873 1333 1876
rect 1396 1807 1403 1923
rect 1156 1663 1163 1703
rect 1173 1663 1187 1673
rect 1156 1660 1187 1663
rect 1156 1656 1183 1660
rect 1113 1440 1127 1453
rect 1116 1436 1123 1440
rect 1176 1407 1183 1656
rect 1256 1647 1263 1734
rect 1416 1747 1423 1853
rect 1296 1706 1303 1733
rect 1336 1700 1343 1703
rect 1333 1687 1347 1700
rect 1256 1436 1263 1553
rect 1316 1527 1323 1573
rect 1136 1327 1143 1403
rect 1093 1220 1107 1233
rect 1096 1216 1103 1220
rect 1076 1107 1083 1183
rect 1156 1183 1163 1273
rect 1147 1176 1163 1183
rect 1176 1167 1183 1233
rect 1096 916 1123 923
rect 976 876 1003 883
rect 976 807 983 876
rect 1116 847 1123 916
rect 1136 787 1143 1093
rect 1196 1087 1203 1434
rect 1216 1167 1223 1213
rect 1256 1180 1263 1183
rect 1253 1167 1267 1180
rect 1176 916 1223 923
rect 1256 916 1263 1132
rect 1296 1107 1303 1183
rect 1056 736 1063 773
rect 976 707 983 733
rect 996 696 1023 703
rect 976 666 983 693
rect 936 367 943 433
rect 976 408 983 613
rect 996 507 1003 696
rect 996 467 1003 493
rect 1176 427 1183 916
rect 1316 787 1323 1073
rect 1276 647 1283 663
rect 1316 647 1323 694
rect 1133 400 1147 413
rect 1136 396 1143 400
rect 1216 366 1223 453
rect 1276 396 1283 633
rect 1336 547 1343 1453
rect 1376 1367 1383 1703
rect 1416 1436 1423 1533
rect 1436 1467 1443 2173
rect 1456 1807 1463 2193
rect 1476 2107 1483 2173
rect 1496 2147 1503 2223
rect 1516 2067 1523 2193
rect 1556 2007 1563 2253
rect 1476 1743 1483 1993
rect 1576 1987 1583 2256
rect 1656 2256 1663 2336
rect 1696 2263 1703 2693
rect 1816 2687 1823 2793
rect 1836 2747 1843 2774
rect 1776 2527 1783 2673
rect 1776 2476 1783 2513
rect 1816 2467 1823 2513
rect 1756 2327 1763 2443
rect 1836 2427 1843 2693
rect 1776 2303 1783 2413
rect 1756 2296 1783 2303
rect 1696 2256 1723 2263
rect 1596 2127 1603 2213
rect 1513 1960 1527 1973
rect 1516 1956 1523 1960
rect 1496 1887 1503 1913
rect 1536 1847 1543 1923
rect 1576 1907 1583 1923
rect 1456 1736 1483 1743
rect 1516 1736 1523 1793
rect 1456 1487 1463 1736
rect 1496 1647 1503 1703
rect 1576 1687 1583 1893
rect 1476 1436 1503 1443
rect 1416 1216 1423 1313
rect 1436 1247 1443 1403
rect 1496 1347 1503 1436
rect 1476 1180 1483 1183
rect 1473 1167 1487 1180
rect 1496 1107 1503 1173
rect 1416 916 1423 1093
rect 1356 847 1363 872
rect 1396 847 1403 883
rect 1336 427 1343 493
rect 1356 467 1363 833
rect 1436 787 1443 883
rect 1456 696 1463 833
rect 1496 666 1503 693
rect 1336 366 1343 413
rect 1396 408 1403 663
rect 1376 396 1393 403
rect 1116 360 1123 363
rect 1113 347 1127 360
rect 756 136 783 143
rect 1036 143 1043 333
rect 1356 227 1363 373
rect 1156 176 1193 183
rect 996 136 1043 143
rect 276 -24 303 -17
rect 456 -24 483 -17
rect 1116 -17 1123 143
rect 1316 -17 1323 143
rect 1376 87 1383 396
rect 1416 307 1423 363
rect 1456 176 1463 352
rect 1496 307 1503 533
rect 1516 366 1523 1473
rect 1536 927 1543 1671
rect 1556 1167 1563 1573
rect 1596 1436 1603 1753
rect 1616 1507 1623 1973
rect 1636 1747 1643 2053
rect 1656 1887 1663 2173
rect 1696 1956 1703 2013
rect 1716 2007 1723 2256
rect 1736 2187 1743 2293
rect 1756 2167 1763 2296
rect 1833 2260 1847 2273
rect 1856 2267 1863 2933
rect 1896 2807 1903 2992
rect 1936 2960 1943 2963
rect 1933 2947 1947 2960
rect 1936 2847 1943 2933
rect 1893 2780 1907 2793
rect 1896 2776 1903 2780
rect 1916 2667 1923 2732
rect 1956 2647 1963 2774
rect 1916 2476 1923 2533
rect 1953 2480 1967 2493
rect 1976 2487 1983 2963
rect 1996 2927 2003 2952
rect 1996 2707 2003 2732
rect 2016 2667 2023 3016
rect 2056 2966 2063 3293
rect 2076 3227 2083 3473
rect 2136 3407 2143 3483
rect 2196 3467 2203 3516
rect 2216 3507 2223 3733
rect 2256 3727 2263 3783
rect 2253 3547 2267 3553
rect 2296 3516 2303 3713
rect 2276 3480 2283 3483
rect 2273 3467 2287 3480
rect 2140 3303 2153 3307
rect 2136 3296 2153 3303
rect 2140 3293 2153 3296
rect 2116 3227 2123 3263
rect 2176 3247 2183 3433
rect 2120 3023 2133 3027
rect 2116 3013 2133 3023
rect 2116 2996 2123 3013
rect 2156 3007 2163 3213
rect 2176 2987 2183 3013
rect 2136 2907 2143 2963
rect 2096 2816 2103 2873
rect 2036 2547 2043 2633
rect 2156 2547 2163 2953
rect 2196 2887 2203 3453
rect 2316 3407 2323 3483
rect 2216 2967 2223 3393
rect 2236 3307 2243 3333
rect 2276 3296 2283 3333
rect 2256 3187 2263 3263
rect 2296 3260 2303 3263
rect 2293 3247 2307 3260
rect 2336 2987 2343 3013
rect 2256 2927 2263 2963
rect 2356 2963 2363 3693
rect 2376 3687 2383 3814
rect 2436 3747 2443 3783
rect 2376 3266 2383 3293
rect 2396 3147 2403 3333
rect 2416 3087 2423 3713
rect 2433 3520 2447 3533
rect 2436 3516 2443 3520
rect 2476 3447 2483 3483
rect 2393 3000 2407 3013
rect 2396 2996 2403 3000
rect 2476 2967 2483 3233
rect 2496 3087 2503 3263
rect 2356 2956 2383 2963
rect 2173 2807 2187 2813
rect 2213 2787 2227 2793
rect 2236 2783 2243 2833
rect 2296 2816 2303 2953
rect 2236 2776 2263 2783
rect 2216 2647 2223 2713
rect 1956 2476 1963 2480
rect 1876 2307 1883 2433
rect 1836 2256 1843 2260
rect 1816 2007 1823 2223
rect 1856 2067 1863 2213
rect 1736 1956 1743 1993
rect 1676 1748 1683 1913
rect 1776 1883 1783 1954
rect 1816 1927 1823 1972
rect 1876 1956 1883 2293
rect 1896 2268 1903 2443
rect 1936 2440 1943 2443
rect 1933 2427 1947 2440
rect 1896 2226 1903 2254
rect 1916 2227 1923 2333
rect 1956 2256 1963 2293
rect 1996 2256 2003 2333
rect 2016 2327 2023 2493
rect 2036 2287 2043 2533
rect 2076 2476 2083 2533
rect 2113 2480 2127 2493
rect 2116 2476 2123 2480
rect 2156 2407 2163 2533
rect 2236 2476 2243 2693
rect 2376 2683 2383 2956
rect 2496 2966 2503 3033
rect 2516 2963 2523 3633
rect 2556 3543 2563 4073
rect 2636 4036 2643 4093
rect 2656 4087 2663 4333
rect 2676 4107 2683 4353
rect 2696 4347 2703 4573
rect 2716 4367 2723 5273
rect 2836 5247 2843 5513
rect 2896 5376 2903 5413
rect 2916 5403 2923 5563
rect 2956 5547 2963 5633
rect 3036 5527 3043 5563
rect 2916 5396 2943 5403
rect 2936 5376 2943 5396
rect 2856 5227 2863 5374
rect 2736 4923 2743 5133
rect 2876 5047 2883 5333
rect 2896 5047 2903 5074
rect 2776 5007 2783 5043
rect 2736 4916 2763 4923
rect 2736 4387 2743 4893
rect 2756 4627 2763 4916
rect 2796 4727 2803 4812
rect 2776 4556 2783 4673
rect 2816 4607 2823 4753
rect 2836 4647 2843 4823
rect 2816 4556 2823 4593
rect 2856 4587 2863 4613
rect 2756 4267 2763 4303
rect 2696 4043 2703 4253
rect 2676 4036 2703 4043
rect 2616 3847 2623 4003
rect 2656 3887 2663 4003
rect 2536 3536 2563 3543
rect 2536 3347 2543 3536
rect 2556 3163 2563 3513
rect 2576 3308 2583 3833
rect 2676 3816 2683 3853
rect 2716 3827 2723 4093
rect 2736 3816 2743 4053
rect 2756 3823 2763 4073
rect 2776 4043 2783 4093
rect 2796 4067 2803 4373
rect 2876 4368 2883 5012
rect 2896 4807 2903 4953
rect 2916 4907 2923 5343
rect 2936 5087 2943 5233
rect 2976 5203 2983 5493
rect 3076 5487 3083 5552
rect 2996 5267 3003 5374
rect 3016 5247 3023 5393
rect 3053 5380 3067 5393
rect 3056 5376 3063 5380
rect 3096 5376 3103 5553
rect 3116 5527 3123 5973
rect 3136 5566 3143 5813
rect 3136 5383 3143 5493
rect 3156 5447 3163 6333
rect 3176 6086 3183 6253
rect 3196 6227 3203 6356
rect 3196 6087 3203 6213
rect 3233 6120 3247 6133
rect 3276 6128 3283 6453
rect 3473 6420 3487 6433
rect 3476 6416 3483 6420
rect 3316 6167 3323 6372
rect 3376 6267 3383 6414
rect 3953 6420 3967 6433
rect 3956 6416 3963 6420
rect 3456 6327 3463 6383
rect 3236 6116 3243 6120
rect 3236 5787 3243 5863
rect 3276 5623 3283 5893
rect 3296 5807 3303 6013
rect 3316 5863 3323 6114
rect 3336 5907 3343 6173
rect 3396 5947 3403 6083
rect 3436 5927 3443 6083
rect 3516 5987 3523 6393
rect 3636 6380 3643 6383
rect 3633 6367 3647 6380
rect 3736 6347 3743 6383
rect 3876 6347 3883 6413
rect 3996 6367 4003 6433
rect 4136 6416 4143 6453
rect 3973 6347 3987 6353
rect 3393 5900 3407 5912
rect 3396 5896 3403 5900
rect 3316 5856 3343 5863
rect 3256 5616 3283 5623
rect 3256 5596 3263 5616
rect 3176 5447 3183 5553
rect 3196 5487 3203 5563
rect 3236 5507 3243 5563
rect 3136 5376 3163 5383
rect 3076 5287 3083 5343
rect 2976 5196 3003 5203
rect 2976 5076 2983 5173
rect 2996 5107 3003 5196
rect 2996 4987 3003 5043
rect 2896 4587 2903 4733
rect 2896 4487 2903 4552
rect 2916 4507 2923 4854
rect 2956 4820 2963 4823
rect 2953 4807 2967 4820
rect 2996 4687 3003 4713
rect 3016 4567 3023 4853
rect 3036 4727 3043 4893
rect 2936 4516 2963 4523
rect 2936 4387 2943 4516
rect 2816 4087 2823 4353
rect 2776 4036 2803 4043
rect 2833 4040 2847 4053
rect 2836 4036 2843 4040
rect 2896 4006 2903 4303
rect 2956 4267 2963 4493
rect 2756 3816 2783 3823
rect 2616 3587 2623 3812
rect 2636 3667 2643 3783
rect 2696 3707 2703 3783
rect 2776 3667 2783 3816
rect 2633 3520 2647 3533
rect 2636 3516 2643 3520
rect 2676 3516 2683 3573
rect 2716 3487 2723 3613
rect 2796 3567 2803 3933
rect 2856 3907 2863 4003
rect 2916 3947 2923 4053
rect 2936 4006 2943 4133
rect 2976 4087 2983 4433
rect 3016 4343 3023 4513
rect 3036 4387 3043 4713
rect 3056 4687 3063 5213
rect 3156 5147 3163 5376
rect 3076 4867 3083 5093
rect 3196 5027 3203 5433
rect 3236 5376 3243 5472
rect 3316 5327 3323 5513
rect 3336 5387 3343 5856
rect 3436 5843 3443 5913
rect 3453 5908 3467 5913
rect 3533 5900 3547 5913
rect 3536 5896 3543 5900
rect 3456 5863 3463 5894
rect 3456 5856 3483 5863
rect 3416 5836 3443 5843
rect 3416 5596 3423 5836
rect 3336 5307 3343 5373
rect 3156 4856 3163 5011
rect 3216 4987 3223 5073
rect 3236 4863 3243 5193
rect 3256 4907 3263 5233
rect 3336 5147 3343 5173
rect 3356 5167 3363 5473
rect 3396 5427 3403 5563
rect 3436 5487 3443 5563
rect 3387 5383 3400 5387
rect 3387 5376 3403 5383
rect 3387 5373 3400 5376
rect 3276 5076 3283 5113
rect 3336 5076 3343 5133
rect 3316 4887 3323 5032
rect 3216 4856 3243 4863
rect 3076 4727 3083 4812
rect 3096 4787 3103 4823
rect 3196 4787 3203 4853
rect 3056 4507 3063 4593
rect 3076 4487 3083 4713
rect 3216 4587 3223 4856
rect 3236 4667 3243 4833
rect 3276 4747 3283 4812
rect 3316 4787 3323 4823
rect 3356 4807 3363 4853
rect 3376 4826 3383 4973
rect 3216 4523 3223 4552
rect 3136 4487 3143 4523
rect 3176 4503 3183 4523
rect 3156 4496 3183 4503
rect 3196 4516 3223 4523
rect 3076 4427 3083 4473
rect 2996 4336 3023 4343
rect 2996 4247 3003 4336
rect 3116 4306 3123 4393
rect 3036 4300 3043 4303
rect 3033 4287 3047 4300
rect 3136 4287 3143 4353
rect 3156 4307 3163 4496
rect 3196 4407 3203 4516
rect 3236 4503 3243 4653
rect 3356 4627 3363 4733
rect 3376 4647 3383 4773
rect 3216 4496 3243 4503
rect 3216 4336 3223 4496
rect 3256 4343 3263 4573
rect 3316 4520 3323 4523
rect 3313 4507 3327 4520
rect 3356 4507 3363 4573
rect 3376 4526 3383 4633
rect 3396 4487 3403 5313
rect 3416 5287 3423 5343
rect 3476 5327 3483 5856
rect 3516 5847 3523 5863
rect 3516 5836 3533 5847
rect 3520 5833 3533 5836
rect 3576 5747 3583 6083
rect 3656 6027 3663 6114
rect 3896 6116 3903 6153
rect 3696 5987 3703 6113
rect 3727 6076 3743 6083
rect 3596 5687 3603 5973
rect 3716 5896 3723 6072
rect 3696 5860 3703 5863
rect 3693 5847 3707 5860
rect 3836 5807 3843 5863
rect 3876 5860 3883 5863
rect 3873 5847 3887 5860
rect 3936 5847 3943 6053
rect 3956 5867 3963 6073
rect 3976 6067 3983 6193
rect 3976 5923 3983 6013
rect 3996 5947 4003 6353
rect 4036 6327 4043 6413
rect 4076 6380 4083 6383
rect 4073 6367 4087 6380
rect 4116 6363 4123 6383
rect 4216 6367 4223 6453
rect 4436 6416 4443 6453
rect 4916 6416 4923 6453
rect 4956 6416 4963 6453
rect 5116 6428 5123 6453
rect 4376 6386 4383 6413
rect 4256 6380 4263 6383
rect 4253 6367 4267 6380
rect 4116 6356 4143 6363
rect 4136 6307 4143 6356
rect 4296 6307 4303 6383
rect 4456 6327 4463 6383
rect 4016 6047 4023 6253
rect 4136 6083 4143 6293
rect 4236 6116 4243 6153
rect 4176 6086 4183 6113
rect 4296 6086 4303 6153
rect 3976 5916 4003 5923
rect 3996 5896 4003 5916
rect 4036 5896 4043 6073
rect 4056 6007 4063 6083
rect 4096 6047 4103 6083
rect 4116 6076 4143 6083
rect 4016 5860 4023 5863
rect 4013 5847 4027 5860
rect 4096 5847 4103 5893
rect 3556 5527 3563 5563
rect 3636 5507 3643 5553
rect 3616 5387 3623 5473
rect 3516 5346 3523 5373
rect 3636 5347 3643 5493
rect 3436 5207 3443 5253
rect 3456 4947 3463 5043
rect 3496 5007 3503 5043
rect 3536 5027 3543 5293
rect 3556 4947 3563 5332
rect 3596 5247 3603 5333
rect 3576 5046 3583 5093
rect 3636 5076 3643 5133
rect 3656 5107 3663 5753
rect 3836 5747 3843 5793
rect 3776 5596 3783 5713
rect 3816 5608 3823 5693
rect 3676 5567 3683 5594
rect 3716 5447 3723 5513
rect 3816 5463 3823 5594
rect 3836 5487 3843 5733
rect 3956 5596 3963 5653
rect 3816 5456 3843 5463
rect 3716 5376 3723 5433
rect 3756 5347 3763 5393
rect 3616 5027 3623 5043
rect 3616 4887 3623 5013
rect 3433 4860 3447 4873
rect 3436 4856 3443 4860
rect 3516 4747 3523 4854
rect 3416 4587 3423 4673
rect 3456 4556 3463 4693
rect 3436 4427 3443 4523
rect 3516 4523 3523 4613
rect 3536 4527 3543 4853
rect 3556 4707 3563 4873
rect 3587 4863 3600 4867
rect 3587 4856 3603 4863
rect 3587 4853 3600 4856
rect 3676 4863 3683 4933
rect 3696 4927 3703 5074
rect 3736 5046 3743 5193
rect 3776 5127 3783 5373
rect 3796 5207 3803 5433
rect 3836 5388 3843 5456
rect 3896 5447 3903 5563
rect 3936 5560 3943 5563
rect 3933 5547 3947 5560
rect 4036 5566 4043 5813
rect 4096 5707 4103 5793
rect 4116 5687 4123 6076
rect 4316 6067 4323 6114
rect 4336 6083 4343 6173
rect 4516 6147 4523 6413
rect 4636 6307 4643 6383
rect 4433 6120 4447 6133
rect 4436 6116 4443 6120
rect 4336 6076 4383 6083
rect 4136 5707 4143 5993
rect 4176 5908 4183 5973
rect 4220 5903 4233 5907
rect 4216 5896 4233 5903
rect 4220 5893 4233 5896
rect 3816 5167 3823 5333
rect 3856 5187 3863 5343
rect 3896 5247 3903 5333
rect 3816 4947 3823 5043
rect 3676 4856 3703 4863
rect 3776 4856 3783 4893
rect 3816 4856 3823 4912
rect 3616 4820 3623 4823
rect 3613 4807 3627 4820
rect 3656 4707 3663 4823
rect 3676 4687 3683 4773
rect 3496 4516 3523 4523
rect 3256 4336 3283 4343
rect 2816 3567 2823 3853
rect 2856 3627 2863 3783
rect 2916 3727 2923 3753
rect 2956 3727 2963 3814
rect 2996 3767 3003 3933
rect 3036 3887 3043 4034
rect 3056 3847 3063 4233
rect 3076 4007 3083 4113
rect 3116 4036 3123 4193
rect 3136 4067 3143 4273
rect 3196 4147 3203 4292
rect 3147 4056 3163 4063
rect 3156 4036 3163 4056
rect 3216 4003 3223 4233
rect 3276 4043 3283 4336
rect 3296 4267 3303 4413
rect 3316 4307 3323 4393
rect 3373 4340 3387 4353
rect 3376 4336 3383 4340
rect 3356 4247 3363 4303
rect 3396 4267 3403 4303
rect 3436 4207 3443 4293
rect 3456 4187 3463 4473
rect 3476 4283 3483 4512
rect 3496 4307 3503 4516
rect 3556 4487 3563 4573
rect 3616 4556 3623 4633
rect 3696 4587 3703 4856
rect 3856 4827 3863 4993
rect 3876 4983 3883 5113
rect 3896 5107 3903 5233
rect 3896 5027 3903 5072
rect 3876 4976 3903 4983
rect 3573 4340 3587 4353
rect 3596 4347 3603 4523
rect 3636 4520 3643 4523
rect 3633 4507 3647 4520
rect 3716 4507 3723 4813
rect 3736 4526 3743 4733
rect 3876 4647 3883 4933
rect 3896 4826 3903 4976
rect 3916 4907 3923 5393
rect 3936 5147 3943 5473
rect 3956 5267 3963 5433
rect 3976 5387 3983 5553
rect 4116 5560 4123 5563
rect 4113 5547 4127 5560
rect 4127 5536 4143 5543
rect 3996 5407 4003 5493
rect 4016 5427 4023 5533
rect 4016 5376 4023 5413
rect 4036 5407 4043 5513
rect 4096 5387 4103 5473
rect 4136 5383 4143 5536
rect 4156 5487 4163 5773
rect 4216 5767 4223 5833
rect 4256 5767 4263 5933
rect 4276 5807 4283 5893
rect 4296 5727 4303 5933
rect 4376 5896 4383 6053
rect 4456 5866 4463 6013
rect 4476 5908 4483 6072
rect 4516 6027 4523 6112
rect 4616 6080 4623 6083
rect 4613 6067 4627 6080
rect 4676 6067 4683 6233
rect 4696 6128 4703 6413
rect 4776 6287 4783 6383
rect 4876 6376 4903 6383
rect 4936 6380 4943 6383
rect 4776 6187 4783 6273
rect 4696 6023 4703 6114
rect 4676 6016 4703 6023
rect 4676 5987 4683 6016
rect 4656 5976 4673 5983
rect 4316 5827 4323 5853
rect 4333 5827 4347 5833
rect 4476 5747 4483 5894
rect 4496 5867 4503 5973
rect 4536 5896 4543 5973
rect 4613 5927 4627 5933
rect 4573 5900 4587 5913
rect 4576 5896 4583 5900
rect 4196 5647 4203 5693
rect 4176 5547 4183 5613
rect 4196 5566 4203 5593
rect 4316 5566 4323 5653
rect 4416 5628 4423 5673
rect 4396 5507 4403 5563
rect 4460 5523 4473 5527
rect 4456 5513 4473 5523
rect 4116 5376 4143 5383
rect 4156 5376 4163 5433
rect 4196 5376 4203 5433
rect 4116 5346 4123 5376
rect 3933 5087 3947 5093
rect 3976 5088 3983 5173
rect 4016 5076 4023 5213
rect 4176 5187 4183 5343
rect 4216 5307 4223 5343
rect 3956 5040 3963 5043
rect 3953 5027 3967 5040
rect 3996 5007 4003 5043
rect 3956 4856 3963 4992
rect 4016 4987 4023 5013
rect 4016 4867 4023 4933
rect 4036 4826 4043 5033
rect 4056 4947 4063 5153
rect 3916 4727 3923 4813
rect 3796 4556 3803 4613
rect 3747 4516 3763 4523
rect 3576 4336 3583 4340
rect 3476 4280 3503 4283
rect 3476 4276 3507 4280
rect 3493 4267 3507 4276
rect 3476 4207 3483 4253
rect 3256 4036 3283 4043
rect 3296 4036 3303 4073
rect 3333 4040 3347 4053
rect 3336 4036 3343 4040
rect 3176 3996 3223 4003
rect 3033 3820 3047 3833
rect 3036 3816 3043 3820
rect 3056 3767 3063 3783
rect 3136 3786 3143 3953
rect 3156 3787 3163 3833
rect 3056 3727 3063 3753
rect 3076 3707 3083 3733
rect 2616 3296 2623 3483
rect 2656 3480 2663 3483
rect 2653 3467 2667 3480
rect 2736 3427 2743 3533
rect 2756 3467 2763 3553
rect 2793 3520 2807 3532
rect 2796 3516 2803 3520
rect 2896 3486 2903 3553
rect 2656 3296 2663 3333
rect 2536 3156 2563 3163
rect 2536 3047 2543 3156
rect 2556 2996 2563 3133
rect 2636 3127 2643 3263
rect 2736 3247 2743 3294
rect 2516 2956 2543 2963
rect 2536 2776 2543 2956
rect 2356 2676 2383 2683
rect 2196 2447 2203 2474
rect 2056 2226 2063 2253
rect 2076 2226 2083 2313
rect 1893 2207 1907 2212
rect 1856 1887 1863 1923
rect 1896 1920 1903 1923
rect 1893 1907 1907 1920
rect 1767 1876 1783 1883
rect 1656 1667 1663 1703
rect 1633 1440 1647 1453
rect 1636 1436 1643 1440
rect 1696 1407 1703 1692
rect 1716 1607 1723 1873
rect 1756 1667 1763 1873
rect 1896 1748 1903 1893
rect 1836 1736 1883 1743
rect 1876 1687 1883 1736
rect 1616 1216 1623 1353
rect 1696 1243 1703 1273
rect 1716 1267 1723 1553
rect 1896 1507 1903 1734
rect 1916 1707 1923 1853
rect 1936 1787 1943 2153
rect 1956 1847 1963 1993
rect 1976 1867 1983 2191
rect 2016 2187 2023 2223
rect 2096 2107 2103 2393
rect 2236 2226 2243 2253
rect 2176 2187 2183 2212
rect 2256 2147 2263 2443
rect 2336 2287 2343 2653
rect 2356 2447 2363 2676
rect 2476 2667 2483 2743
rect 2496 2587 2503 2633
rect 2516 2607 2523 2743
rect 2376 2427 2383 2513
rect 2396 2507 2403 2553
rect 2396 2347 2403 2493
rect 2473 2480 2487 2493
rect 2476 2476 2483 2480
rect 2536 2476 2543 2513
rect 2053 1960 2067 1973
rect 2056 1956 2063 1960
rect 2116 1927 2123 1954
rect 2036 1827 2043 1923
rect 2076 1920 2083 1923
rect 2073 1907 2087 1920
rect 2156 1907 2163 2133
rect 2196 1956 2203 2093
rect 1956 1687 1963 1703
rect 1776 1436 1783 1493
rect 1956 1487 1963 1673
rect 2016 1647 2023 1733
rect 2036 1527 2043 1773
rect 2056 1706 2063 1833
rect 2176 1728 2183 1853
rect 1976 1436 1983 1513
rect 1756 1247 1763 1403
rect 1856 1367 1863 1434
rect 1676 1236 1703 1243
rect 1596 1180 1603 1183
rect 1593 1167 1607 1180
rect 1576 916 1583 953
rect 1596 880 1603 883
rect 1593 867 1607 880
rect 1636 847 1643 1013
rect 1636 723 1643 833
rect 1616 716 1643 723
rect 1616 696 1623 716
rect 1656 703 1663 953
rect 1676 867 1683 1236
rect 1813 1220 1827 1233
rect 1816 1216 1823 1220
rect 1696 1107 1703 1214
rect 1876 1183 1883 1233
rect 1716 928 1723 1172
rect 1796 1107 1803 1183
rect 1836 1147 1843 1183
rect 1856 1176 1883 1183
rect 1756 916 1763 953
rect 1736 847 1743 883
rect 1727 816 1753 823
rect 1796 787 1803 833
rect 1656 696 1683 703
rect 1676 666 1683 696
rect 1536 467 1543 513
rect 1536 367 1543 453
rect 1676 407 1683 533
rect 1716 447 1723 733
rect 1776 696 1783 733
rect 1816 696 1823 973
rect 1836 787 1843 914
rect 1856 887 1863 1176
rect 1896 1027 1903 1434
rect 2036 1406 2043 1473
rect 1956 1347 1963 1403
rect 1996 1216 2003 1253
rect 1976 1180 1983 1183
rect 1973 1167 1987 1180
rect 2016 1147 2023 1183
rect 2056 1167 2063 1213
rect 2076 1186 2083 1633
rect 2136 1627 2143 1703
rect 2156 1667 2163 1693
rect 2116 1436 2123 1473
rect 2136 1467 2143 1613
rect 2156 1448 2163 1513
rect 2196 1403 2203 1513
rect 2136 1367 2143 1403
rect 2176 1396 2203 1403
rect 2096 1163 2103 1313
rect 2116 1247 2123 1273
rect 2136 1267 2143 1353
rect 2176 1327 2183 1396
rect 2196 1287 2203 1373
rect 2196 1216 2203 1273
rect 2216 1247 2223 1833
rect 2233 1720 2247 1733
rect 2236 1716 2243 1720
rect 2236 1387 2243 1653
rect 2276 1587 2283 2173
rect 2296 2107 2303 2223
rect 2376 2187 2383 2293
rect 2436 2268 2443 2443
rect 2496 2440 2503 2443
rect 2493 2427 2507 2440
rect 2396 2187 2403 2254
rect 2496 2236 2503 2353
rect 2516 2247 2523 2333
rect 2296 1847 2303 2093
rect 2416 2007 2423 2173
rect 2536 2147 2543 2333
rect 2556 2236 2563 2653
rect 2576 2307 2583 2732
rect 2596 2667 2603 2833
rect 2536 2047 2543 2133
rect 2596 2107 2603 2632
rect 2616 2347 2623 2963
rect 2656 2887 2663 3073
rect 2676 2907 2683 3033
rect 2676 2847 2683 2893
rect 2696 2883 2703 3193
rect 2776 2996 2783 3113
rect 2696 2876 2723 2883
rect 2696 2803 2703 2853
rect 2676 2796 2703 2803
rect 2676 2776 2683 2796
rect 2716 2776 2723 2876
rect 2696 2707 2703 2743
rect 2736 2740 2743 2743
rect 2733 2727 2747 2740
rect 2776 2727 2783 2833
rect 2796 2746 2803 2933
rect 2816 2847 2823 3013
rect 2836 2867 2843 3133
rect 2856 3027 2863 3373
rect 2916 3308 2923 3653
rect 2936 3486 2943 3613
rect 3036 3487 3043 3533
rect 2996 3296 3003 3413
rect 3056 3387 3063 3593
rect 3116 3547 3123 3773
rect 3176 3767 3183 3793
rect 3196 3767 3203 3996
rect 3236 3828 3243 3992
rect 3256 3847 3263 4036
rect 3296 3783 3303 3953
rect 3376 3927 3383 4053
rect 3396 3848 3403 4053
rect 3416 3847 3423 4173
rect 3480 4063 3493 4067
rect 3476 4053 3493 4063
rect 3476 4036 3483 4053
rect 3536 4006 3543 4113
rect 3596 4067 3603 4293
rect 3616 4087 3623 4473
rect 3636 4147 3643 4413
rect 3656 4247 3663 4353
rect 3676 4347 3683 4493
rect 3696 4348 3703 4413
rect 3613 4040 3627 4052
rect 3676 4043 3683 4293
rect 3716 4247 3723 4303
rect 3616 4036 3623 4040
rect 3656 4036 3683 4043
rect 3636 3883 3643 4003
rect 3696 3947 3703 4093
rect 3756 4047 3763 4516
rect 3876 4467 3883 4573
rect 3896 4547 3903 4713
rect 3776 4207 3783 4333
rect 3796 4107 3803 4433
rect 3776 4036 3783 4073
rect 3816 4036 3823 4193
rect 3916 4127 3923 4653
rect 3956 4556 3963 4593
rect 3996 4556 4003 4593
rect 3936 4306 3943 4393
rect 3796 3967 3803 4003
rect 3636 3876 3663 3883
rect 3436 3847 3443 3873
rect 3553 3847 3567 3853
rect 3216 3707 3223 3783
rect 3276 3776 3303 3783
rect 2936 3147 2943 3252
rect 2936 3027 2943 3133
rect 2976 3127 2983 3263
rect 2856 2827 2863 2992
rect 2936 2887 2943 2963
rect 2916 2776 2923 2833
rect 2816 2567 2823 2774
rect 2856 2740 2863 2743
rect 2853 2727 2867 2740
rect 2907 2715 2933 2722
rect 2876 2488 2883 2653
rect 2936 2527 2943 2573
rect 2736 2476 2763 2483
rect 2756 2347 2763 2476
rect 2956 2446 2963 2733
rect 2976 2488 2983 3013
rect 2996 2788 3003 2993
rect 3016 2927 3023 3013
rect 3036 3007 3043 3333
rect 3056 3266 3063 3293
rect 3076 3187 3083 3533
rect 3173 3520 3187 3533
rect 3176 3516 3183 3520
rect 3216 3487 3223 3653
rect 3236 3487 3243 3713
rect 3256 3347 3263 3553
rect 3296 3516 3303 3633
rect 3316 3547 3323 3833
rect 3336 3747 3343 3793
rect 3356 3567 3363 3833
rect 3433 3820 3447 3833
rect 3436 3816 3443 3820
rect 3333 3520 3347 3533
rect 3336 3516 3343 3520
rect 3316 3480 3323 3483
rect 3276 3427 3283 3473
rect 3313 3467 3327 3480
rect 3120 3323 3133 3327
rect 3116 3313 3133 3323
rect 3116 3296 3123 3313
rect 3176 3256 3203 3263
rect 3196 3247 3203 3256
rect 3073 3000 3087 3013
rect 3176 3008 3183 3113
rect 3076 2996 3083 3000
rect 3116 2996 3163 3003
rect 3056 2887 3063 2963
rect 3156 2947 3163 2996
rect 2996 2507 3003 2774
rect 3036 2727 3043 2743
rect 3027 2716 3043 2727
rect 3027 2713 3040 2716
rect 3096 2667 3103 2913
rect 3116 2747 3123 2873
rect 3156 2847 3163 2912
rect 3176 2847 3183 2994
rect 3196 2967 3203 3233
rect 3236 3008 3243 3273
rect 3256 3266 3263 3312
rect 3316 3296 3323 3333
rect 3356 3308 3363 3393
rect 3336 3260 3343 3263
rect 3333 3247 3347 3260
rect 3316 3236 3333 3243
rect 3316 3027 3323 3236
rect 3356 3207 3363 3233
rect 3396 3227 3403 3753
rect 3416 3467 3423 3533
rect 3436 3407 3443 3733
rect 3476 3667 3483 3813
rect 3496 3787 3503 3833
rect 3556 3816 3563 3833
rect 3476 3516 3483 3613
rect 3516 3607 3523 3793
rect 3636 3787 3643 3853
rect 3576 3780 3583 3783
rect 3573 3767 3587 3780
rect 3656 3703 3663 3876
rect 3676 3707 3683 3813
rect 3636 3696 3663 3703
rect 3516 3516 3523 3593
rect 3496 3480 3503 3483
rect 3436 3207 3443 3333
rect 3456 3247 3463 3473
rect 3493 3467 3507 3480
rect 3536 3427 3543 3483
rect 3416 3067 3423 3133
rect 3393 3000 3407 3013
rect 3396 2996 3403 3000
rect 3256 2960 3263 2963
rect 3253 2947 3267 2960
rect 3296 2907 3303 2953
rect 3356 2867 3363 2993
rect 3416 2927 3423 2963
rect 3456 2887 3463 2933
rect 2896 2268 2903 2443
rect 2976 2387 2983 2474
rect 3096 2443 3103 2513
rect 3056 2436 3103 2443
rect 2736 2240 2743 2243
rect 2733 2227 2747 2240
rect 2836 2236 2863 2243
rect 2316 1907 2323 1953
rect 2376 1867 2383 1923
rect 2416 1867 2423 1993
rect 2456 1867 2463 1953
rect 2540 1923 2553 1927
rect 2496 1920 2503 1923
rect 2493 1907 2507 1920
rect 2536 1916 2553 1923
rect 2540 1913 2553 1916
rect 2576 1907 2583 2073
rect 2676 1963 2683 2093
rect 2836 2087 2843 2236
rect 2936 2227 2943 2293
rect 2976 2226 2983 2333
rect 3076 2256 3083 2293
rect 3116 2256 3123 2313
rect 3136 2263 3143 2813
rect 3196 2776 3203 2813
rect 3436 2743 3443 2853
rect 3476 2847 3483 2994
rect 3496 2927 3503 2994
rect 3516 2967 3523 3133
rect 3556 2996 3563 3053
rect 3596 3047 3603 3433
rect 3616 3276 3623 3653
rect 3636 3627 3643 3696
rect 3656 3547 3663 3673
rect 3756 3647 3763 3783
rect 3836 3627 3843 3893
rect 3856 3747 3863 3873
rect 3876 3687 3883 4053
rect 3936 4036 3943 4213
rect 3956 4187 3963 4493
rect 3976 4347 3983 4523
rect 4013 4507 4027 4513
rect 4036 4447 4043 4753
rect 4016 4336 4023 4413
rect 4056 4347 4063 4673
rect 4036 4296 4063 4303
rect 3976 4036 3983 4073
rect 4056 4027 4063 4296
rect 4076 4227 4083 5133
rect 4096 5046 4103 5073
rect 4127 4876 4153 4883
rect 4096 4747 4103 4823
rect 4156 4747 4163 4823
rect 4093 4567 4107 4573
rect 4136 4556 4143 4613
rect 4176 4587 4183 4853
rect 4216 4767 4223 5173
rect 4236 5046 4243 5213
rect 4256 5127 4263 5473
rect 4296 5346 4303 5433
rect 4353 5380 4367 5393
rect 4356 5376 4363 5380
rect 4456 5367 4463 5513
rect 4336 5307 4343 5343
rect 4476 5187 4483 5453
rect 4496 5427 4503 5594
rect 4536 5563 4543 5773
rect 4576 5608 4583 5833
rect 4596 5627 4603 5813
rect 4616 5747 4623 5913
rect 4613 5600 4627 5613
rect 4636 5603 4643 5933
rect 4656 5847 4663 5976
rect 4696 5947 4703 5993
rect 4716 5947 4723 6173
rect 4816 6167 4823 6213
rect 4776 6116 4783 6152
rect 4836 6086 4843 6133
rect 4756 6063 4763 6083
rect 4756 6056 4783 6063
rect 4716 5923 4723 5933
rect 4716 5916 4743 5923
rect 4736 5896 4743 5916
rect 4776 5867 4783 6056
rect 4676 5787 4683 5853
rect 4756 5807 4763 5853
rect 4616 5596 4623 5600
rect 4636 5596 4663 5603
rect 4536 5556 4563 5563
rect 4556 5407 4563 5556
rect 4576 5343 4583 5473
rect 4596 5347 4603 5374
rect 4496 5307 4503 5343
rect 4556 5336 4583 5343
rect 4476 5076 4483 5173
rect 4516 5076 4523 5133
rect 4256 5007 4263 5053
rect 4296 4927 4303 5043
rect 4416 4947 4423 4973
rect 4287 4874 4293 4887
rect 4280 4873 4300 4874
rect 4356 4856 4403 4863
rect 4173 4560 4187 4573
rect 4196 4567 4203 4653
rect 4176 4556 4183 4560
rect 3956 3947 3963 4003
rect 3996 4000 4003 4003
rect 3993 3987 4007 4000
rect 3916 3816 3923 3873
rect 3936 3667 3943 3783
rect 3636 3496 3663 3503
rect 3636 3307 3643 3333
rect 3656 3283 3663 3496
rect 3676 3347 3683 3494
rect 3916 3387 3923 3613
rect 4016 3563 4023 3913
rect 4056 3816 4063 3873
rect 4076 3847 4083 4173
rect 4096 4167 4103 4373
rect 4116 4247 4123 4393
rect 4156 4336 4163 4433
rect 4196 4336 4203 4453
rect 4216 4427 4223 4593
rect 4236 4568 4243 4813
rect 4296 4803 4303 4823
rect 4276 4796 4303 4803
rect 4276 4667 4283 4796
rect 4236 4347 4243 4554
rect 4096 4007 4103 4113
rect 4136 4107 4143 4293
rect 4216 4247 4223 4303
rect 4133 4040 4147 4053
rect 4136 4036 4143 4040
rect 4156 3823 4163 3992
rect 4136 3816 4183 3823
rect 4076 3707 4083 3783
rect 4116 3763 4123 3772
rect 4096 3756 4123 3763
rect 4016 3556 4043 3563
rect 3656 3276 3683 3283
rect 3616 3067 3623 3213
rect 3636 3123 3643 3233
rect 3656 3147 3663 3276
rect 3716 3267 3723 3293
rect 3996 3287 4003 3373
rect 4016 3303 4023 3534
rect 4036 3327 4043 3556
rect 4056 3507 4063 3633
rect 4076 3527 4083 3613
rect 4056 3327 4063 3453
rect 4076 3427 4083 3473
rect 4096 3427 4103 3756
rect 4116 3607 4123 3713
rect 4176 3647 4183 3816
rect 4196 3587 4203 4153
rect 4256 4143 4263 4633
rect 4296 4607 4303 4773
rect 4336 4667 4343 4791
rect 4376 4787 4383 4813
rect 4367 4713 4373 4727
rect 4333 4560 4347 4573
rect 4336 4556 4343 4560
rect 4376 4487 4383 4692
rect 4396 4667 4403 4856
rect 4416 4787 4423 4933
rect 4416 4687 4423 4752
rect 4436 4707 4443 4913
rect 4456 4867 4463 4993
rect 4476 4947 4483 5013
rect 4473 4807 4487 4812
rect 4516 4787 4523 4823
rect 4476 4727 4483 4753
rect 4456 4687 4463 4713
rect 4396 4526 4403 4573
rect 4276 4147 4283 4333
rect 4296 4307 4303 4433
rect 4416 4343 4423 4652
rect 4436 4607 4443 4653
rect 4516 4647 4523 4773
rect 4433 4587 4447 4593
rect 4453 4560 4467 4573
rect 4493 4560 4507 4573
rect 4536 4567 4543 4733
rect 4456 4556 4463 4560
rect 4496 4556 4503 4560
rect 4396 4336 4423 4343
rect 4436 4307 4443 4334
rect 4376 4300 4383 4303
rect 4373 4287 4387 4300
rect 4236 4136 4263 4143
rect 4216 3583 4223 4093
rect 4236 3887 4243 4136
rect 4276 4067 4283 4133
rect 4296 4036 4303 4272
rect 4316 4127 4323 4253
rect 4356 4007 4363 4053
rect 4316 4000 4323 4003
rect 4313 3987 4327 4000
rect 4256 3816 4263 3913
rect 4316 3727 4323 3783
rect 4356 3767 4363 3972
rect 4376 3927 4383 4013
rect 4376 3787 4383 3814
rect 4396 3807 4403 4153
rect 4436 4048 4443 4093
rect 4456 4067 4463 4473
rect 4476 4467 4483 4523
rect 4536 4467 4543 4513
rect 4556 4447 4563 5093
rect 4576 5046 4583 5133
rect 4576 4587 4583 4873
rect 4596 4643 4603 5153
rect 4616 5087 4623 5533
rect 4656 5383 4663 5596
rect 4676 5507 4683 5613
rect 4696 5547 4703 5733
rect 4756 5596 4763 5653
rect 4796 5607 4803 5633
rect 4816 5566 4823 6033
rect 4836 5907 4843 6072
rect 4856 6007 4863 6213
rect 4876 6086 4883 6376
rect 4933 6367 4947 6380
rect 4996 6367 5003 6414
rect 4936 6147 4943 6313
rect 4933 6120 4947 6133
rect 4996 6128 5003 6353
rect 4936 6116 4943 6120
rect 5116 6116 5123 6173
rect 4876 6047 4883 6072
rect 4876 5896 4883 6012
rect 4996 5967 5003 6114
rect 5056 6080 5063 6083
rect 5053 6067 5067 6080
rect 5096 6047 5103 6083
rect 5156 6067 5163 6414
rect 5176 6287 5183 6393
rect 5196 6387 5203 6414
rect 5236 6327 5243 6383
rect 5276 6307 5283 6383
rect 5436 6347 5443 6372
rect 5496 6287 5503 6372
rect 4836 5567 4843 5853
rect 4856 5807 4863 5863
rect 4896 5747 4903 5863
rect 4936 5787 4943 5953
rect 5013 5943 5027 5953
rect 4996 5940 5027 5943
rect 4996 5936 5023 5940
rect 4996 5903 5003 5936
rect 4976 5896 5003 5903
rect 5013 5900 5027 5913
rect 5016 5896 5023 5900
rect 4956 5667 4963 5893
rect 4976 5847 4983 5896
rect 5036 5807 5043 5852
rect 5076 5807 5083 5863
rect 4816 5507 4823 5552
rect 4636 5376 4663 5383
rect 4696 5376 4703 5433
rect 4636 5107 4643 5376
rect 4716 5340 4723 5343
rect 4676 5307 4683 5332
rect 4713 5327 4727 5340
rect 4776 5303 4783 5374
rect 4796 5327 4803 5393
rect 4756 5296 4783 5303
rect 4656 5076 4663 5213
rect 4696 5087 4703 5173
rect 4680 5043 4693 5047
rect 4676 5036 4693 5043
rect 4680 5033 4693 5036
rect 4696 4907 4703 4953
rect 4673 4860 4687 4873
rect 4676 4856 4683 4860
rect 4596 4636 4623 4643
rect 4576 4547 4583 4573
rect 4596 4527 4603 4613
rect 4616 4567 4623 4636
rect 4636 4607 4643 4773
rect 4656 4747 4663 4823
rect 4716 4627 4723 5113
rect 4736 4827 4743 5293
rect 4756 5187 4763 5296
rect 4756 4987 4763 5173
rect 4796 5167 4803 5292
rect 4816 5167 4823 5493
rect 4836 5283 4843 5532
rect 4856 5467 4863 5633
rect 4873 5607 4887 5613
rect 5016 5596 5023 5773
rect 4896 5507 4903 5553
rect 4976 5523 4983 5563
rect 4976 5516 5003 5523
rect 4896 5376 4903 5493
rect 4856 5307 4863 5332
rect 4836 5276 4863 5283
rect 4796 5076 4803 5153
rect 4776 4863 4783 5013
rect 4816 4967 4823 5032
rect 4856 4927 4863 5276
rect 4756 4856 4783 4863
rect 4813 4860 4827 4873
rect 4816 4856 4823 4860
rect 4653 4560 4667 4573
rect 4696 4568 4703 4593
rect 4656 4556 4663 4560
rect 4533 4407 4547 4413
rect 4533 4400 4553 4407
rect 4536 4396 4553 4400
rect 4540 4393 4553 4396
rect 4516 4336 4523 4393
rect 4576 4363 4583 4473
rect 4547 4356 4583 4363
rect 4596 4267 4603 4334
rect 4516 4036 4523 4153
rect 4536 4047 4543 4173
rect 4616 4103 4623 4513
rect 4636 4287 4643 4491
rect 4736 4467 4743 4593
rect 4676 4300 4683 4303
rect 4716 4300 4723 4303
rect 4656 4207 4663 4293
rect 4673 4287 4687 4300
rect 4713 4287 4727 4300
rect 4756 4267 4763 4856
rect 4840 4823 4853 4827
rect 4836 4813 4853 4823
rect 4796 4727 4803 4791
rect 4596 4096 4623 4103
rect 4456 3967 4463 4003
rect 4496 4000 4503 4003
rect 4493 3987 4507 4000
rect 4496 3947 4503 3973
rect 4513 3967 4527 3973
rect 4456 3816 4463 3853
rect 4496 3816 4503 3893
rect 4536 3847 4543 3933
rect 4556 3786 4563 4013
rect 4336 3667 4343 3733
rect 4216 3576 4243 3583
rect 4156 3440 4163 3443
rect 4153 3427 4167 3440
rect 4016 3296 4063 3303
rect 3856 3280 3863 3283
rect 3853 3267 3867 3280
rect 3956 3276 3983 3283
rect 3876 3223 3883 3273
rect 3856 3216 3883 3223
rect 3636 3116 3663 3123
rect 3656 2967 3663 3116
rect 3576 2927 3583 2963
rect 3696 2943 3703 3033
rect 3676 2936 3703 2943
rect 3476 2788 3483 2833
rect 3576 2776 3583 2833
rect 3416 2736 3443 2743
rect 3396 2446 3403 2593
rect 3136 2256 3163 2263
rect 2896 2200 2903 2203
rect 2893 2187 2907 2200
rect 2676 1956 2703 1963
rect 2633 1927 2647 1933
rect 2616 1916 2633 1923
rect 2507 1896 2523 1903
rect 2320 1443 2333 1447
rect 2316 1436 2333 1443
rect 2320 1433 2333 1436
rect 2356 1407 2363 1573
rect 2516 1527 2523 1896
rect 2536 1716 2543 1893
rect 2556 1726 2563 1853
rect 2256 1347 2263 1393
rect 2236 1186 2243 1253
rect 2076 1156 2103 1163
rect 1936 916 1943 1113
rect 1836 707 1843 773
rect 1856 666 1863 793
rect 1896 667 1903 833
rect 1996 787 2003 1033
rect 2016 847 2023 1092
rect 2076 916 2083 1156
rect 2256 1147 2263 1213
rect 2056 880 2063 883
rect 2053 867 2067 880
rect 2056 807 2063 853
rect 2096 827 2103 883
rect 2136 787 2143 953
rect 2276 916 2283 1373
rect 2376 1303 2383 1434
rect 2396 1327 2403 1473
rect 2436 1436 2443 1513
rect 2516 1487 2523 1513
rect 2476 1436 2483 1473
rect 2556 1423 2563 1673
rect 2576 1487 2583 1683
rect 2516 1403 2523 1423
rect 2556 1416 2583 1423
rect 2496 1396 2523 1403
rect 2496 1307 2503 1396
rect 2376 1296 2403 1303
rect 2376 1228 2383 1273
rect 2396 1227 2403 1296
rect 2316 1107 2323 1183
rect 2396 1067 2403 1173
rect 2176 827 2183 914
rect 2316 887 2323 1053
rect 2216 867 2223 883
rect 2216 787 2223 853
rect 2336 847 2343 1013
rect 1956 696 1963 773
rect 1996 676 2003 713
rect 1796 660 1803 663
rect 1793 647 1807 660
rect 1736 396 1743 633
rect 2036 547 2043 713
rect 2076 683 2083 773
rect 2336 686 2343 733
rect 2056 676 2083 683
rect 2356 676 2363 1033
rect 2416 1027 2423 1214
rect 2456 1107 2463 1293
rect 2516 1247 2523 1273
rect 2513 1220 2527 1233
rect 2516 1216 2523 1220
rect 2496 1167 2503 1183
rect 2556 1167 2563 1333
rect 2496 1156 2513 1167
rect 2500 1153 2513 1156
rect 2576 1147 2583 1416
rect 2616 1223 2623 1916
rect 2696 1827 2703 1956
rect 2736 1787 2743 1993
rect 2796 1956 2823 1963
rect 2816 1847 2823 1956
rect 2836 1947 2843 1993
rect 2856 1907 2863 2033
rect 2896 1947 2903 2073
rect 2956 2007 2963 2153
rect 2956 1956 2963 1993
rect 3016 1988 3023 2173
rect 3096 2167 3103 2223
rect 3096 2127 3103 2153
rect 3156 2107 3163 2256
rect 3176 2226 3183 2373
rect 3196 2268 3203 2443
rect 3436 2367 3443 2736
rect 3556 2527 3563 2743
rect 3616 2707 3623 2774
rect 3556 2487 3563 2513
rect 3233 2268 3247 2273
rect 3433 2260 3447 2273
rect 3436 2256 3443 2260
rect 3476 2256 3483 2353
rect 3516 2287 3523 2413
rect 3636 2327 3643 2853
rect 3676 2803 3683 2936
rect 3656 2796 3683 2803
rect 3656 2587 3663 2796
rect 3693 2780 3707 2793
rect 3736 2788 3743 2933
rect 3756 2927 3763 2963
rect 3796 2956 3823 2963
rect 3816 2887 3823 2956
rect 3836 2947 3843 2994
rect 3696 2776 3703 2780
rect 3716 2607 3723 2743
rect 3776 2687 3783 2793
rect 3796 2727 3803 2833
rect 3816 2827 3823 2873
rect 3856 2867 3863 3216
rect 3956 3127 3963 3276
rect 3956 3116 3973 3127
rect 3960 3113 3973 3116
rect 4016 3107 4023 3243
rect 3876 2966 3883 3013
rect 3996 2966 4003 2993
rect 3856 2740 3863 2743
rect 3816 2627 3823 2733
rect 3853 2727 3867 2740
rect 3796 2616 3813 2623
rect 3653 2480 3667 2493
rect 3656 2476 3663 2480
rect 3716 2476 3743 2483
rect 3676 2407 3683 2443
rect 3736 2307 3743 2476
rect 3756 2407 3763 2473
rect 3776 2367 3783 2573
rect 3796 2446 3803 2616
rect 3820 2603 3833 2607
rect 3816 2600 3833 2603
rect 3813 2593 3833 2600
rect 3813 2587 3827 2593
rect 3896 2587 3903 2793
rect 3916 2787 3923 2931
rect 4016 2867 4023 3053
rect 3916 2667 3923 2773
rect 3836 2507 3843 2553
rect 3833 2480 3847 2493
rect 3836 2476 3843 2480
rect 3593 2260 3607 2273
rect 3596 2256 3603 2260
rect 3376 2226 3383 2253
rect 3256 2187 3263 2223
rect 3307 2216 3323 2223
rect 2936 1920 2943 1923
rect 2933 1907 2947 1920
rect 2976 1887 2983 1923
rect 2976 1767 2983 1813
rect 2693 1720 2707 1733
rect 2696 1716 2703 1720
rect 2676 1627 2683 1714
rect 2736 1687 2743 1733
rect 3076 1727 3083 1974
rect 3316 1827 3323 2216
rect 3416 2187 3423 2223
rect 3616 2187 3623 2223
rect 3696 2207 3703 2293
rect 3756 2256 3763 2313
rect 3736 2127 3743 2223
rect 3776 2220 3783 2223
rect 3773 2207 3787 2220
rect 3356 1847 3363 1943
rect 3376 1887 3383 2053
rect 3396 1936 3423 1943
rect 3396 1863 3403 1936
rect 3436 1907 3443 2093
rect 3536 1943 3543 2073
rect 3516 1936 3543 1943
rect 3636 1936 3643 1993
rect 3456 1887 3463 1934
rect 3776 1867 3783 1973
rect 3396 1856 3453 1863
rect 2876 1587 2883 1723
rect 2976 1716 3003 1723
rect 2756 1416 2763 1533
rect 2936 1487 2943 1573
rect 2976 1567 2983 1716
rect 3136 1716 3163 1723
rect 3156 1567 3163 1716
rect 2856 1327 2863 1454
rect 2956 1427 2963 1553
rect 2976 1407 2983 1532
rect 3076 1436 3083 1533
rect 3156 1407 3163 1473
rect 3196 1467 3203 1533
rect 3236 1487 3243 1593
rect 3256 1527 3263 1672
rect 3253 1440 3267 1453
rect 3256 1436 3263 1440
rect 2596 1216 2623 1223
rect 2636 1216 2643 1313
rect 2416 916 2423 1013
rect 2396 847 2403 883
rect 1676 366 1683 393
rect 1836 366 1843 493
rect 1933 400 1947 413
rect 1936 396 1943 400
rect 1716 327 1723 363
rect 1567 176 1583 183
rect 1556 147 1563 174
rect 1656 156 1663 313
rect 1916 267 1923 363
rect 1956 307 1963 363
rect 1713 160 1727 173
rect 1996 166 2003 253
rect 1716 156 1723 160
rect 2016 156 2023 513
rect 2036 366 2043 433
rect 2053 427 2067 433
rect 2096 408 2103 653
rect 2136 396 2143 433
rect 2116 183 2123 363
rect 2196 347 2203 513
rect 2276 396 2283 533
rect 2116 180 2143 183
rect 2116 176 2147 180
rect 2133 166 2147 176
rect 2156 156 2163 331
rect 2296 267 2303 363
rect 2336 287 2343 352
rect 2376 347 2383 533
rect 2396 263 2403 632
rect 2456 567 2463 953
rect 2476 646 2483 913
rect 2516 827 2523 1093
rect 2536 928 2543 1113
rect 2556 987 2563 1093
rect 2576 967 2583 1133
rect 2596 847 2603 1216
rect 2876 1216 2883 1353
rect 2896 1227 2903 1313
rect 2656 1180 2663 1183
rect 2696 1180 2703 1183
rect 2653 1167 2667 1180
rect 2693 1167 2707 1180
rect 2736 1167 2743 1213
rect 2776 1167 2783 1214
rect 2816 1180 2823 1183
rect 2813 1167 2827 1180
rect 2856 1107 2863 1183
rect 2896 1107 2903 1133
rect 2936 1047 2943 1214
rect 2656 886 2663 953
rect 2816 886 2823 913
rect 2576 696 2583 733
rect 2496 527 2503 694
rect 2656 666 2663 833
rect 2696 827 2703 883
rect 2716 708 2723 793
rect 2736 696 2743 773
rect 2596 567 2603 663
rect 2456 360 2463 363
rect 2453 347 2467 360
rect 2396 256 2423 263
rect 1616 -17 1623 143
rect 2416 126 2423 256
rect 2436 247 2443 333
rect 2516 207 2523 553
rect 2533 487 2547 493
rect 2576 396 2583 513
rect 2596 447 2603 553
rect 2616 408 2623 633
rect 2656 487 2663 652
rect 2756 527 2763 663
rect 2796 427 2803 872
rect 2936 747 2943 1033
rect 2956 1007 2963 1313
rect 2996 1228 3003 1253
rect 3036 1216 3043 1313
rect 3056 1267 3063 1403
rect 3176 1347 3183 1434
rect 3236 1327 3243 1403
rect 3336 1307 3343 1434
rect 3356 1427 3363 1553
rect 3376 1227 3383 1473
rect 3396 1387 3403 1813
rect 3436 1716 3443 1833
rect 3496 1720 3523 1723
rect 3496 1716 3527 1720
rect 3416 1467 3423 1633
rect 3456 1627 3463 1712
rect 3513 1707 3527 1716
rect 3447 1536 3473 1543
rect 3456 1468 3463 1513
rect 3453 1440 3467 1454
rect 3456 1436 3463 1440
rect 3416 1227 3423 1403
rect 3516 1287 3523 1313
rect 3556 1287 3563 1753
rect 3656 1736 3663 1793
rect 3796 1767 3803 1893
rect 3816 1847 3823 1943
rect 3836 1787 3843 2413
rect 3856 2327 3863 2443
rect 3856 2207 3863 2313
rect 3896 2287 3903 2313
rect 3916 2283 3923 2513
rect 3936 2307 3943 2853
rect 3993 2780 4007 2793
rect 3996 2776 4003 2780
rect 4036 2776 4043 3133
rect 4056 3107 4063 3296
rect 4076 3087 4083 3413
rect 4236 3407 4243 3576
rect 4256 3423 4263 3633
rect 4276 3447 4283 3513
rect 4296 3483 4303 3633
rect 4336 3516 4343 3653
rect 4376 3603 4383 3752
rect 4436 3707 4443 3783
rect 4436 3647 4443 3693
rect 4456 3687 4463 3753
rect 4456 3623 4463 3652
rect 4516 3627 4523 3733
rect 4427 3616 4463 3623
rect 4376 3596 4403 3603
rect 4376 3516 4383 3553
rect 4396 3547 4403 3596
rect 4416 3527 4423 3592
rect 4536 3583 4543 3673
rect 4516 3576 4543 3583
rect 4416 3516 4433 3527
rect 4420 3513 4433 3516
rect 4296 3476 4323 3483
rect 4256 3416 4283 3423
rect 4236 3396 4253 3407
rect 4240 3393 4253 3396
rect 4076 2996 4083 3033
rect 4096 3027 4103 3313
rect 4116 2996 4123 3313
rect 4276 3303 4283 3416
rect 4296 3307 4303 3413
rect 4316 3363 4323 3476
rect 4356 3447 4363 3483
rect 4396 3480 4403 3483
rect 4393 3467 4407 3480
rect 4456 3447 4463 3533
rect 4476 3467 4483 3573
rect 4516 3547 4523 3576
rect 4496 3387 4503 3533
rect 4536 3516 4543 3553
rect 4556 3547 4563 3772
rect 4576 3707 4583 4053
rect 4596 4006 4603 4096
rect 4656 4036 4663 4073
rect 4696 4036 4703 4093
rect 4716 4067 4723 4233
rect 4736 4167 4743 4253
rect 4756 4127 4763 4232
rect 4776 4227 4783 4613
rect 4796 4567 4803 4613
rect 4836 4607 4843 4813
rect 4856 4747 4863 4792
rect 4876 4627 4883 5213
rect 4827 4597 4843 4607
rect 4827 4593 4840 4597
rect 4813 4560 4827 4572
rect 4853 4560 4867 4573
rect 4896 4563 4903 5093
rect 4916 5087 4923 5273
rect 4936 5107 4943 5433
rect 4956 5287 4963 5493
rect 4976 5347 4983 5374
rect 4996 5267 5003 5516
rect 5036 5407 5043 5733
rect 5056 5447 5063 5653
rect 5076 5647 5083 5793
rect 5116 5747 5123 5894
rect 5136 5787 5143 5933
rect 5156 5827 5163 6053
rect 5176 5947 5183 6153
rect 5196 5947 5203 6213
rect 5236 6116 5243 6213
rect 5316 6087 5323 6273
rect 5336 6067 5343 6173
rect 5396 6123 5403 6173
rect 5376 6116 5403 6123
rect 5456 6116 5463 6213
rect 5496 6167 5503 6273
rect 5516 6247 5523 6413
rect 5576 6128 5583 6433
rect 5993 6420 6007 6433
rect 5996 6416 6003 6420
rect 6336 6416 6343 6453
rect 6473 6420 6487 6433
rect 6496 6427 6503 6456
rect 6476 6416 6483 6420
rect 5656 6203 5663 6372
rect 5696 6227 5703 6273
rect 5736 6247 5743 6413
rect 5896 6386 5903 6413
rect 5776 6207 5783 6383
rect 5816 6363 5823 6383
rect 5796 6356 5823 6363
rect 5796 6307 5803 6356
rect 5976 6347 5983 6383
rect 5656 6196 5683 6203
rect 5256 5896 5263 5933
rect 5196 5787 5203 5863
rect 5233 5847 5247 5852
rect 5296 5847 5303 5953
rect 5156 5596 5163 5633
rect 5076 5427 5083 5573
rect 5116 5507 5123 5594
rect 5216 5560 5223 5563
rect 5133 5543 5147 5552
rect 5133 5540 5163 5543
rect 5136 5536 5163 5540
rect 5036 5376 5043 5393
rect 5136 5367 5143 5513
rect 5156 5447 5163 5536
rect 5176 5527 5183 5552
rect 5213 5547 5227 5560
rect 5256 5547 5263 5813
rect 5276 5587 5283 5833
rect 5316 5787 5323 5913
rect 5356 5907 5363 6114
rect 5376 6047 5383 6116
rect 5616 6116 5623 6153
rect 5436 6047 5443 6083
rect 5436 5896 5443 6033
rect 5336 5807 5343 5853
rect 5376 5847 5383 5863
rect 5373 5827 5387 5833
rect 5416 5807 5423 5863
rect 5333 5767 5347 5772
rect 5296 5563 5303 5693
rect 5496 5687 5503 6053
rect 5516 5847 5523 6113
rect 5576 5928 5583 5993
rect 5596 5967 5603 6083
rect 5616 5896 5623 6013
rect 5676 5963 5683 6196
rect 5696 6047 5703 6113
rect 5716 6086 5723 6173
rect 5796 6128 5803 6293
rect 5747 6123 5760 6127
rect 5747 6116 5763 6123
rect 5747 6113 5760 6116
rect 5816 6047 5823 6083
rect 5856 6027 5863 6193
rect 5876 5987 5883 6313
rect 5896 6086 5903 6233
rect 6036 6167 6043 6353
rect 5936 6116 5943 6153
rect 6056 6147 6063 6413
rect 6216 6386 6223 6413
rect 6116 6247 6123 6383
rect 6156 6380 6163 6383
rect 6153 6367 6167 6380
rect 6236 6307 6243 6414
rect 6316 6267 6323 6383
rect 6456 6380 6463 6383
rect 6453 6367 6467 6380
rect 6113 6120 6127 6133
rect 6116 6116 6123 6120
rect 5667 5956 5683 5963
rect 5516 5667 5523 5833
rect 5556 5807 5563 5863
rect 5596 5827 5603 5863
rect 5556 5667 5563 5793
rect 5596 5707 5603 5813
rect 5376 5608 5383 5633
rect 5296 5556 5323 5563
rect 4996 5087 5003 5153
rect 5056 5127 5063 5253
rect 5096 5147 5103 5343
rect 4916 4847 4923 4953
rect 4936 4867 4943 4933
rect 4976 4927 4983 5043
rect 5016 4883 5023 5073
rect 5036 5007 5043 5053
rect 5056 4943 5063 5113
rect 5116 5076 5123 5273
rect 5136 5107 5143 5233
rect 5156 5227 5163 5433
rect 5216 5376 5223 5473
rect 5276 5427 5283 5533
rect 5296 5387 5303 5513
rect 5176 5307 5183 5374
rect 5316 5343 5323 5556
rect 5356 5527 5363 5563
rect 5336 5447 5343 5493
rect 5436 5467 5443 5594
rect 5476 5507 5483 5613
rect 5513 5600 5527 5613
rect 5516 5596 5523 5600
rect 5616 5567 5623 5653
rect 5636 5567 5643 5753
rect 5356 5423 5363 5453
rect 5456 5447 5463 5473
rect 5476 5423 5483 5453
rect 5516 5427 5523 5533
rect 5276 5340 5283 5343
rect 5236 5267 5243 5332
rect 5273 5327 5287 5340
rect 5296 5336 5323 5343
rect 5336 5416 5363 5423
rect 5456 5416 5483 5423
rect 5156 5047 5163 5213
rect 4953 4860 4967 4873
rect 4996 4876 5023 4883
rect 5036 4936 5063 4943
rect 4956 4856 4963 4860
rect 4996 4856 5003 4876
rect 5036 4867 5043 4936
rect 5053 4907 5067 4913
rect 5020 4823 5033 4827
rect 5016 4816 5033 4823
rect 5020 4813 5033 4816
rect 4916 4747 4923 4812
rect 4933 4807 4947 4812
rect 5056 4787 5063 4853
rect 5076 4827 5083 5033
rect 4936 4727 4943 4753
rect 4913 4667 4927 4673
rect 4816 4556 4823 4560
rect 4856 4556 4863 4560
rect 4896 4556 4923 4563
rect 4756 4007 4763 4053
rect 4593 3987 4607 3992
rect 4596 3747 4603 3873
rect 4616 3827 4623 3953
rect 4636 3847 4643 3992
rect 4676 3843 4683 4003
rect 4716 4000 4723 4003
rect 4713 3987 4727 4000
rect 4756 3927 4763 3972
rect 4676 3836 4703 3843
rect 4696 3816 4703 3836
rect 4616 3607 4623 3673
rect 4636 3547 4643 3733
rect 4736 3727 4743 3813
rect 4756 3767 4763 3833
rect 4573 3520 4587 3533
rect 4576 3516 4583 3520
rect 4516 3387 4523 3473
rect 4556 3427 4563 3483
rect 4596 3447 4603 3483
rect 4636 3387 4643 3493
rect 4656 3487 4663 3613
rect 4676 3483 4683 3693
rect 4696 3627 4703 3653
rect 4716 3607 4723 3673
rect 4736 3627 4743 3653
rect 4776 3603 4783 4213
rect 4796 4187 4803 4513
rect 4836 4447 4843 4523
rect 4896 4447 4903 4472
rect 4816 4407 4823 4433
rect 4816 4396 4833 4407
rect 4820 4393 4833 4396
rect 4816 4347 4823 4373
rect 4853 4340 4867 4353
rect 4856 4336 4863 4340
rect 4896 4336 4903 4393
rect 4916 4387 4923 4556
rect 4936 4487 4943 4573
rect 4956 4547 4963 4673
rect 4976 4667 4983 4753
rect 4973 4587 4987 4593
rect 5056 4556 5063 4633
rect 5076 4567 5083 4653
rect 4976 4516 5003 4523
rect 4956 4467 4963 4493
rect 4976 4487 4983 4516
rect 5036 4467 5043 4523
rect 4946 4452 4947 4460
rect 4933 4443 4947 4452
rect 4933 4440 4983 4443
rect 4936 4436 4983 4440
rect 4936 4367 4943 4393
rect 4920 4366 4943 4367
rect 4927 4356 4943 4366
rect 4927 4353 4940 4356
rect 4956 4347 4963 4413
rect 4976 4367 4983 4436
rect 4876 4282 4883 4303
rect 4916 4300 4923 4303
rect 4847 4275 4883 4282
rect 4913 4287 4927 4300
rect 4816 4147 4823 4253
rect 4816 4043 4823 4133
rect 4856 4067 4863 4173
rect 4796 4036 4823 4043
rect 4833 4040 4847 4053
rect 4836 4036 4843 4040
rect 4796 3987 4803 4036
rect 4916 4036 4923 4093
rect 4896 4000 4903 4003
rect 4893 3987 4907 4000
rect 4813 3947 4827 3953
rect 4796 3847 4803 3933
rect 4856 3887 4863 3971
rect 4776 3596 4803 3603
rect 4696 3527 4703 3592
rect 4776 3516 4783 3573
rect 4796 3567 4803 3596
rect 4816 3527 4823 3633
rect 4676 3476 4703 3483
rect 4487 3376 4503 3387
rect 4487 3373 4500 3376
rect 4316 3356 4343 3363
rect 4256 3296 4283 3303
rect 4336 3276 4343 3356
rect 4136 3256 4163 3263
rect 4136 3207 4143 3256
rect 4053 2787 4067 2793
rect 3976 2687 3983 2743
rect 4016 2607 4023 2743
rect 3956 2427 3963 2573
rect 4013 2480 4027 2493
rect 4016 2476 4023 2480
rect 4076 2446 4083 2893
rect 4096 2887 4103 2963
rect 4176 2827 4183 3153
rect 4296 3107 4303 3243
rect 4216 2887 4223 3033
rect 4316 3027 4323 3233
rect 4316 2966 4323 2992
rect 4336 2907 4343 3213
rect 4356 3167 4363 3373
rect 4436 3227 4443 3273
rect 4456 3147 4463 3283
rect 4596 3276 4643 3283
rect 4596 3247 4603 3276
rect 4476 3087 4483 3173
rect 4393 3000 4407 3013
rect 4396 2996 4403 3000
rect 4556 3007 4563 3113
rect 4356 2927 4363 2994
rect 4576 2996 4583 3133
rect 4656 3043 4663 3452
rect 4696 3283 4703 3476
rect 4756 3447 4763 3483
rect 4696 3276 4723 3283
rect 4716 3223 4723 3276
rect 4696 3216 4723 3223
rect 4656 3036 4683 3043
rect 4613 3000 4627 3013
rect 4616 2996 4623 3000
rect 4207 2803 4220 2807
rect 4207 2793 4223 2803
rect 4216 2776 4223 2793
rect 4156 2567 4163 2743
rect 4256 2667 4263 2753
rect 4116 2446 4123 2493
rect 3996 2407 4003 2432
rect 3916 2276 3943 2283
rect 3936 2256 3943 2276
rect 3876 2226 3883 2253
rect 4016 2247 4023 2293
rect 4036 2268 4043 2432
rect 4276 2427 4283 2853
rect 4436 2847 4443 2913
rect 4456 2887 4463 2963
rect 4353 2780 4367 2793
rect 4356 2776 4363 2780
rect 4296 2687 4303 2773
rect 4436 2743 4443 2833
rect 4536 2807 4543 2973
rect 4656 2966 4663 3013
rect 4493 2780 4507 2793
rect 4496 2776 4503 2780
rect 4536 2776 4543 2793
rect 4436 2736 4483 2743
rect 4296 2427 4303 2593
rect 4376 2476 4383 2653
rect 4416 2527 4423 2573
rect 4396 2446 4403 2493
rect 3956 2127 3963 2223
rect 3716 1706 3723 1753
rect 3796 1736 3803 1753
rect 3676 1647 3683 1692
rect 3816 1567 3823 1703
rect 3116 1196 3143 1203
rect 2976 1127 2983 1173
rect 3076 1127 3083 1163
rect 3136 1047 3143 1196
rect 3127 1036 3143 1047
rect 3127 1033 3140 1036
rect 3016 916 3023 973
rect 2987 883 3000 887
rect 2987 876 3003 883
rect 2987 873 3000 876
rect 3033 867 3047 872
rect 2876 696 2883 733
rect 2836 647 2843 694
rect 2996 667 3003 853
rect 3056 696 3063 733
rect 3076 727 3083 853
rect 3096 843 3103 913
rect 3136 880 3143 883
rect 3133 867 3147 880
rect 3176 863 3183 883
rect 3156 856 3183 863
rect 3156 843 3163 856
rect 3096 836 3163 843
rect 3116 666 3123 713
rect 3196 696 3203 773
rect 3236 696 3243 1203
rect 3296 883 3303 973
rect 3376 967 3383 1213
rect 3416 1200 3443 1203
rect 3416 1196 3447 1200
rect 3476 1196 3503 1203
rect 3433 1187 3447 1196
rect 3436 1107 3443 1173
rect 3436 947 3443 993
rect 3427 916 3443 923
rect 3296 876 3323 883
rect 3373 843 3387 853
rect 3356 840 3387 843
rect 3356 836 3383 840
rect 3276 696 3283 833
rect 3436 827 3443 916
rect 3456 867 3463 1033
rect 3476 886 3483 933
rect 3396 696 3403 793
rect 3436 696 3443 733
rect 2836 587 2843 633
rect 2536 347 2543 394
rect 2456 156 2463 193
rect 2476 87 2483 154
rect 2616 146 2623 233
rect 2656 176 2663 313
rect 2676 267 2683 394
rect 2696 367 2703 413
rect 2733 400 2747 413
rect 2736 396 2743 400
rect 2696 247 2703 273
rect 2796 87 2803 173
rect 2816 143 2823 313
rect 2836 307 2843 433
rect 2856 227 2863 413
rect 2936 396 2943 493
rect 3036 367 3043 663
rect 3076 507 3083 652
rect 3216 487 3223 663
rect 3256 627 3263 663
rect 3416 647 3423 663
rect 3256 567 3263 613
rect 3056 396 3083 403
rect 2916 327 2923 363
rect 2896 216 2903 253
rect 2956 183 2963 213
rect 3036 203 3043 353
rect 3056 327 3063 396
rect 3176 356 3203 363
rect 3196 267 3203 356
rect 3036 196 3063 203
rect 2936 176 2963 183
rect 3056 176 3063 196
rect 2956 146 2963 176
rect 3156 146 3163 253
rect 3276 207 3283 493
rect 3296 396 3303 433
rect 3376 403 3383 473
rect 3356 396 3383 403
rect 3376 327 3383 396
rect 3416 307 3423 633
rect 3456 607 3463 663
rect 3496 527 3503 1196
rect 3736 1183 3743 1273
rect 3796 1227 3803 1513
rect 3856 1423 3863 1833
rect 3876 1567 3883 1773
rect 3896 1527 3903 2033
rect 3916 1887 3923 1993
rect 3956 1827 3963 2113
rect 3976 1926 3983 2133
rect 4016 2067 4023 2233
rect 4056 2226 4063 2393
rect 4116 2256 4123 2313
rect 4096 2220 4103 2223
rect 4093 2207 4107 2220
rect 4196 2167 4203 2411
rect 4356 2407 4363 2443
rect 4216 2187 4223 2353
rect 4236 2226 4243 2313
rect 4336 2296 4343 2353
rect 4016 1983 4023 2053
rect 4056 1987 4063 2053
rect 4016 1976 4043 1983
rect 4036 1956 4043 1976
rect 4096 1963 4103 2113
rect 4087 1956 4103 1963
rect 3956 1667 3963 1703
rect 3996 1627 4003 1733
rect 3916 1423 3923 1493
rect 3836 1416 3863 1423
rect 3896 1416 3923 1423
rect 3736 1176 3763 1183
rect 3796 1107 3803 1213
rect 3596 916 3603 1073
rect 3696 923 3703 993
rect 3696 916 3723 923
rect 3576 827 3583 883
rect 3596 696 3603 733
rect 3633 700 3647 713
rect 3636 696 3643 700
rect 3576 660 3583 663
rect 3573 647 3587 660
rect 3676 663 3683 914
rect 3836 867 3843 1373
rect 3856 1047 3863 1253
rect 3896 1216 3903 1333
rect 3936 1216 3943 1433
rect 3996 1406 4003 1553
rect 4036 1527 4043 1813
rect 4136 1807 4143 2153
rect 4196 2047 4203 2093
rect 4256 1987 4263 2293
rect 4396 2263 4403 2393
rect 4376 2256 4403 2263
rect 4156 1927 4163 1954
rect 4216 1887 4223 1923
rect 4296 1827 4303 2133
rect 4316 2067 4323 2193
rect 4316 1926 4323 1973
rect 4396 1956 4403 2233
rect 4416 2027 4423 2413
rect 4436 1968 4443 2493
rect 4456 2447 4463 2736
rect 4516 2527 4523 2732
rect 4556 2607 4563 2653
rect 4507 2503 4520 2507
rect 4507 2493 4523 2503
rect 4516 2476 4523 2493
rect 4556 2487 4563 2513
rect 4576 2487 4583 2793
rect 4596 2623 4603 2963
rect 4676 2847 4683 3036
rect 4696 2963 4703 3216
rect 4736 3023 4743 3413
rect 4796 3387 4803 3483
rect 4716 3020 4743 3023
rect 4713 3016 4743 3020
rect 4713 3007 4727 3016
rect 4756 2996 4763 3053
rect 4776 3027 4783 3353
rect 4796 3047 4803 3133
rect 4816 3067 4823 3393
rect 4836 3127 4843 3753
rect 4856 3528 4863 3653
rect 4896 3587 4903 3952
rect 4956 3843 4963 4033
rect 4936 3836 4963 3843
rect 4916 3747 4923 3814
rect 4936 3786 4943 3836
rect 4976 3823 4983 4332
rect 4996 4147 5003 4413
rect 5016 4347 5023 4373
rect 5033 4348 5047 4353
rect 5076 4336 5083 4413
rect 5096 4387 5103 4873
rect 5196 4856 5203 5213
rect 5256 5076 5263 5293
rect 5296 5287 5303 5336
rect 5336 5303 5343 5416
rect 5456 5376 5463 5416
rect 5493 5387 5507 5393
rect 5356 5327 5363 5374
rect 5396 5340 5403 5343
rect 5393 5327 5407 5340
rect 5433 5327 5447 5332
rect 5327 5296 5343 5303
rect 5316 5227 5323 5293
rect 5316 5046 5323 5173
rect 5216 5007 5223 5033
rect 5236 4967 5243 5043
rect 5336 4987 5343 5272
rect 5376 5227 5383 5253
rect 5476 5227 5483 5313
rect 5376 5107 5383 5173
rect 5436 5076 5443 5113
rect 5476 5047 5483 5213
rect 5247 4956 5263 4963
rect 5116 4527 5123 4813
rect 5136 4787 5143 4823
rect 5173 4807 5187 4812
rect 5176 4747 5183 4772
rect 5236 4767 5243 4854
rect 5136 4667 5143 4733
rect 5256 4667 5263 4956
rect 5276 4807 5283 4913
rect 5336 4856 5343 4973
rect 5307 4823 5320 4827
rect 5307 4816 5323 4823
rect 5356 4820 5363 4823
rect 5307 4813 5320 4816
rect 5353 4807 5367 4820
rect 5296 4687 5303 4773
rect 5356 4747 5363 4772
rect 5136 4343 5143 4653
rect 5216 4556 5223 4633
rect 5336 4587 5343 4693
rect 5376 4667 5383 4812
rect 5396 4763 5403 5013
rect 5416 4868 5423 5043
rect 5456 4903 5463 5033
rect 5496 4987 5503 5193
rect 5516 5088 5523 5413
rect 5536 5307 5543 5453
rect 5576 5427 5583 5563
rect 5656 5523 5663 5953
rect 5736 5896 5743 5973
rect 5716 5827 5723 5863
rect 5756 5787 5763 5863
rect 5856 5787 5863 5894
rect 5876 5827 5883 5863
rect 5936 5847 5943 5863
rect 5956 5847 5963 5993
rect 5996 5903 6003 6083
rect 6036 6047 6043 6114
rect 6056 5927 6063 5953
rect 6076 5908 6083 6114
rect 6236 6087 6243 6114
rect 6136 6007 6143 6083
rect 6216 6076 6233 6083
rect 5996 5896 6023 5903
rect 5936 5836 5953 5847
rect 5940 5833 5953 5836
rect 5776 5567 5783 5733
rect 5796 5567 5803 5693
rect 5876 5667 5883 5813
rect 5916 5596 5923 5773
rect 5976 5683 5983 5833
rect 5996 5827 6003 5873
rect 6016 5847 6023 5896
rect 6056 5860 6063 5863
rect 6096 5860 6103 5863
rect 6053 5847 6067 5860
rect 6093 5847 6107 5860
rect 6136 5767 6143 5853
rect 6096 5687 6103 5713
rect 6156 5707 6163 6013
rect 5976 5676 6003 5683
rect 5687 5556 5703 5563
rect 5647 5516 5663 5523
rect 5636 5467 5643 5513
rect 5676 5507 5683 5553
rect 5593 5380 5607 5393
rect 5596 5376 5603 5380
rect 5636 5376 5643 5432
rect 5656 5387 5663 5473
rect 5576 5340 5583 5343
rect 5573 5327 5587 5340
rect 5616 5227 5623 5343
rect 5676 5327 5683 5453
rect 5653 5307 5667 5313
rect 5616 5147 5623 5213
rect 5656 5187 5663 5233
rect 5516 5047 5523 5074
rect 5536 4927 5543 4953
rect 5436 4896 5463 4903
rect 5436 4823 5443 4896
rect 5436 4816 5463 4823
rect 5396 4756 5413 4763
rect 5356 4563 5363 4593
rect 5336 4556 5363 4563
rect 5376 4556 5383 4632
rect 5416 4567 5423 4753
rect 5436 4687 5443 4793
rect 5236 4520 5243 4523
rect 5233 4507 5247 4520
rect 5276 4407 5283 4493
rect 5296 4487 5303 4513
rect 5316 4427 5323 4553
rect 5336 4503 5343 4556
rect 5396 4520 5403 4523
rect 5393 4507 5407 4520
rect 5336 4496 5353 4503
rect 5376 4500 5393 4503
rect 5373 4496 5393 4500
rect 5116 4336 5163 4343
rect 5016 4087 5023 4293
rect 5056 4287 5063 4303
rect 5067 4280 5083 4283
rect 5067 4276 5087 4280
rect 5073 4267 5087 4276
rect 5096 4223 5103 4303
rect 5116 4247 5123 4273
rect 5136 4227 5143 4292
rect 5096 4216 5123 4223
rect 5056 4036 5063 4133
rect 5096 4036 5103 4133
rect 5116 4127 5123 4216
rect 5156 4207 5163 4336
rect 5136 4103 5143 4192
rect 5176 4143 5183 4393
rect 5276 4363 5283 4393
rect 5256 4356 5283 4363
rect 5196 4267 5203 4353
rect 5256 4336 5263 4356
rect 5240 4285 5260 4287
rect 5247 4282 5260 4285
rect 5247 4273 5263 4282
rect 5233 4223 5247 4233
rect 5216 4220 5247 4223
rect 5213 4216 5243 4220
rect 5213 4207 5227 4216
rect 5116 4096 5143 4103
rect 5156 4136 5183 4143
rect 5116 4047 5123 4096
rect 4996 3927 5003 4033
rect 4956 3816 4983 3823
rect 5016 3816 5023 3992
rect 5036 3867 5043 4003
rect 4956 3727 4963 3816
rect 5036 3747 5043 3783
rect 5076 3707 5083 3873
rect 5096 3786 5103 3973
rect 5116 3643 5123 3953
rect 5136 3927 5143 4073
rect 5156 3967 5163 4136
rect 5156 3847 5163 3932
rect 5176 3907 5183 4113
rect 5196 3987 5203 4193
rect 5256 4087 5263 4273
rect 5276 4147 5283 4303
rect 5213 4040 5227 4053
rect 5273 4040 5287 4053
rect 5216 4036 5223 4040
rect 5276 4036 5283 4040
rect 5296 3983 5303 4273
rect 5316 4267 5323 4292
rect 5276 3976 5303 3983
rect 5116 3636 5143 3643
rect 5136 3607 5143 3636
rect 4876 3307 4883 3553
rect 4893 3547 4907 3552
rect 4856 3247 4863 3263
rect 4796 2996 4803 3033
rect 4816 3007 4823 3053
rect 4856 3027 4863 3233
rect 4696 2956 4723 2963
rect 4616 2746 4623 2833
rect 4696 2788 4703 2933
rect 4647 2783 4660 2787
rect 4647 2776 4663 2783
rect 4647 2773 4660 2776
rect 4716 2747 4723 2956
rect 4676 2707 4683 2732
rect 4596 2616 4623 2623
rect 4536 2440 4543 2443
rect 4533 2427 4547 2440
rect 4576 2427 4583 2452
rect 4596 2447 4603 2593
rect 4496 2356 4543 2363
rect 4496 2307 4503 2356
rect 4516 2287 4523 2333
rect 4536 2327 4543 2356
rect 4456 2147 4463 2254
rect 4076 1667 4083 1703
rect 4116 1587 4123 1703
rect 3996 1228 4003 1392
rect 4076 1267 4083 1403
rect 4136 1327 4143 1473
rect 4036 1216 4083 1223
rect 3916 1147 3923 1183
rect 3956 1007 3963 1183
rect 3996 927 4003 973
rect 3936 880 3943 883
rect 3776 840 3783 843
rect 3773 827 3787 840
rect 3856 787 3863 872
rect 3933 867 3947 880
rect 3696 666 3703 713
rect 3816 696 3823 753
rect 3836 707 3843 733
rect 3656 656 3683 663
rect 3656 587 3663 656
rect 3716 567 3723 694
rect 3376 176 3383 292
rect 3436 227 3443 433
rect 3556 403 3563 553
rect 3456 396 3483 403
rect 3536 396 3563 403
rect 3456 247 3463 396
rect 3556 307 3563 396
rect 3513 180 3527 193
rect 3516 176 3523 180
rect 2816 136 2843 143
rect 3076 107 3083 143
rect 3236 107 3243 143
rect 3356 107 3363 143
rect 3536 107 3543 132
rect 3596 127 3603 193
rect 2476 47 2483 73
rect 3616 47 3623 413
rect 3636 366 3643 533
rect 3796 487 3803 663
rect 3856 447 3863 773
rect 3876 547 3883 693
rect 3896 666 3903 853
rect 3956 696 3963 833
rect 3996 707 4003 913
rect 3896 607 3903 652
rect 3976 567 3983 663
rect 4016 647 4023 1133
rect 4036 967 4043 1216
rect 4096 916 4103 1033
rect 4136 916 4143 1053
rect 4156 928 4163 1773
rect 4296 1748 4303 1813
rect 4196 1436 4203 1733
rect 4236 1507 4243 1703
rect 4336 1627 4343 1954
rect 4376 1827 4383 1923
rect 4476 1787 4483 2213
rect 4556 2207 4563 2223
rect 4547 2193 4563 2207
rect 4536 2107 4543 2153
rect 4556 2047 4563 2193
rect 4376 1706 4383 1773
rect 4496 1743 4503 1953
rect 4516 1787 4523 1993
rect 4576 1983 4583 2213
rect 4596 1988 4603 2393
rect 4616 2007 4623 2616
rect 4696 2567 4703 2733
rect 4736 2607 4743 2963
rect 4836 2927 4843 2983
rect 4836 2827 4843 2873
rect 4856 2816 4863 2933
rect 4876 2887 4883 3252
rect 4896 3203 4903 3472
rect 5036 3467 5043 3573
rect 4976 3407 4983 3443
rect 4896 3196 4923 3203
rect 4916 3027 4923 3196
rect 4753 2767 4767 2773
rect 4756 2667 4763 2732
rect 4636 2087 4643 2553
rect 4656 2263 4663 2353
rect 4776 2327 4783 2813
rect 4916 2667 4923 2973
rect 4936 2947 4943 3293
rect 5056 3287 5063 3533
rect 5136 3516 5143 3553
rect 5156 3547 5163 3673
rect 5176 3627 5183 3753
rect 5196 3727 5203 3783
rect 5216 3747 5223 3773
rect 5216 3523 5223 3712
rect 5236 3687 5243 3813
rect 5207 3516 5223 3523
rect 5076 3276 5083 3493
rect 5216 3487 5223 3516
rect 5176 3467 5183 3483
rect 5236 3467 5243 3513
rect 5256 3507 5263 3913
rect 5176 3456 5193 3467
rect 5180 3453 5193 3456
rect 5236 3427 5243 3453
rect 5276 3407 5283 3976
rect 5316 3947 5323 4213
rect 5336 4048 5343 4293
rect 5356 4187 5363 4493
rect 5373 4487 5387 4496
rect 5356 4147 5363 4173
rect 5336 4007 5343 4034
rect 5336 3816 5343 3893
rect 5356 3823 5363 4112
rect 5376 4107 5383 4473
rect 5396 4287 5403 4472
rect 5416 4347 5423 4513
rect 5436 4507 5443 4633
rect 5456 4487 5463 4816
rect 5476 4627 5483 4823
rect 5516 4820 5523 4823
rect 5513 4807 5527 4820
rect 5476 4467 5483 4613
rect 5496 4567 5503 4633
rect 5516 4607 5523 4713
rect 5596 4627 5603 4853
rect 5507 4493 5513 4507
rect 5436 4348 5443 4433
rect 5473 4340 5487 4353
rect 5496 4347 5503 4472
rect 5576 4407 5583 4533
rect 5476 4336 5483 4340
rect 5456 4267 5463 4303
rect 5387 4043 5400 4047
rect 5387 4036 5403 4043
rect 5387 4033 5400 4036
rect 5476 4027 5483 4273
rect 5516 4087 5523 4393
rect 5376 3843 5383 3993
rect 5416 3987 5423 4003
rect 5416 3976 5433 3987
rect 5420 3973 5433 3976
rect 5456 3963 5463 3993
rect 5436 3956 5463 3963
rect 5376 3836 5403 3843
rect 5356 3816 5383 3823
rect 5316 3643 5323 3783
rect 5296 3636 5323 3643
rect 5296 3527 5303 3636
rect 5336 3516 5343 3633
rect 5376 3527 5383 3816
rect 5396 3767 5403 3836
rect 5416 3786 5423 3853
rect 5396 3487 5403 3732
rect 5416 3587 5423 3772
rect 5436 3747 5443 3956
rect 5456 3847 5463 3933
rect 5476 3867 5483 4013
rect 5496 4007 5503 4033
rect 5516 4027 5523 4073
rect 5536 4047 5543 4333
rect 5556 4067 5563 4353
rect 5596 4347 5603 4512
rect 5616 4367 5623 4953
rect 5636 4927 5643 5033
rect 5656 4907 5663 5073
rect 5676 4967 5683 5253
rect 5696 5127 5703 5533
rect 5736 5527 5743 5563
rect 5716 5388 5723 5493
rect 5756 5467 5763 5553
rect 5776 5407 5783 5473
rect 5796 5376 5803 5493
rect 5816 5487 5823 5593
rect 5856 5447 5863 5563
rect 5716 5307 5723 5374
rect 5776 5340 5783 5343
rect 5716 5207 5723 5272
rect 5736 5243 5743 5333
rect 5773 5327 5787 5340
rect 5736 5236 5763 5243
rect 5696 4947 5703 5074
rect 5736 5076 5743 5213
rect 5756 5207 5763 5236
rect 5796 5027 5803 5313
rect 5816 5167 5823 5343
rect 5876 5327 5883 5533
rect 5916 5427 5923 5513
rect 5936 5467 5943 5533
rect 5956 5447 5963 5673
rect 5976 5567 5983 5653
rect 5933 5388 5947 5393
rect 5973 5380 5987 5393
rect 5996 5383 6003 5676
rect 6096 5608 6103 5673
rect 6176 5647 6183 5893
rect 6196 5866 6203 5973
rect 6216 5907 6223 6076
rect 6296 6067 6303 6083
rect 6296 6056 6313 6067
rect 6300 6053 6313 6056
rect 6336 5947 6343 6073
rect 6276 5896 6283 5933
rect 6336 5827 6343 5893
rect 6356 5847 6363 6133
rect 6196 5747 6203 5813
rect 6376 5807 6383 6353
rect 6496 6116 6503 6173
rect 6396 6067 6403 6114
rect 6436 6027 6443 6083
rect 6476 6047 6483 6083
rect 6436 5896 6443 5953
rect 6416 5807 6423 5863
rect 6516 5847 6523 5893
rect 6293 5787 6307 5793
rect 6036 5487 6043 5563
rect 5976 5376 5983 5380
rect 5996 5376 6023 5383
rect 5833 5127 5847 5133
rect 5816 5007 5823 5093
rect 5696 4856 5703 4893
rect 5656 4727 5663 4793
rect 5636 4587 5643 4693
rect 5656 4647 5663 4673
rect 5633 4567 5647 4573
rect 5716 4567 5723 4633
rect 5676 4520 5683 4523
rect 5673 4507 5687 4520
rect 5696 4423 5703 4493
rect 5716 4487 5723 4513
rect 5676 4416 5703 4423
rect 5587 4336 5603 4347
rect 5633 4340 5647 4353
rect 5676 4347 5683 4416
rect 5636 4336 5643 4340
rect 5587 4333 5600 4336
rect 5576 4087 5583 4293
rect 5636 4187 5643 4253
rect 5656 4167 5663 4303
rect 5676 4207 5683 4293
rect 5616 4047 5623 4073
rect 5547 4003 5560 4007
rect 5547 3996 5563 4003
rect 5596 4000 5603 4003
rect 5547 3993 5560 3996
rect 5593 3987 5607 4000
rect 5613 3987 5627 3993
rect 5533 3927 5547 3933
rect 5556 3907 5563 3973
rect 5516 3856 5523 3893
rect 5576 3823 5583 3973
rect 5636 3967 5643 4133
rect 5676 4083 5683 4193
rect 5696 4167 5703 4393
rect 5716 4387 5723 4473
rect 5716 4127 5723 4352
rect 5736 4087 5743 4953
rect 5756 4847 5763 4913
rect 5776 4807 5783 4973
rect 5836 4967 5843 5053
rect 5856 5047 5863 5293
rect 5876 5076 5883 5193
rect 5896 5107 5903 5153
rect 5916 5127 5923 5333
rect 5936 5088 5943 5313
rect 6016 5307 6023 5376
rect 5916 5023 5923 5043
rect 5916 5016 5943 5023
rect 5836 4856 5843 4893
rect 5816 4820 5823 4823
rect 5856 4820 5863 4823
rect 5813 4807 5827 4820
rect 5853 4807 5867 4820
rect 5756 4527 5763 4554
rect 5756 4343 5763 4433
rect 5776 4367 5783 4733
rect 5816 4583 5823 4633
rect 5836 4607 5843 4753
rect 5856 4667 5863 4772
rect 5876 4587 5883 4753
rect 5896 4647 5903 4872
rect 5816 4576 5843 4583
rect 5793 4567 5807 4573
rect 5836 4556 5843 4576
rect 5916 4563 5923 4993
rect 5936 4807 5943 5016
rect 5956 4867 5963 5093
rect 5976 4987 5983 5193
rect 5996 5187 6003 5273
rect 5996 4967 6003 5113
rect 6016 4907 6023 5272
rect 6036 5103 6043 5433
rect 6076 5407 6083 5563
rect 6136 5447 6143 5633
rect 6156 5527 6163 5613
rect 6213 5600 6227 5613
rect 6216 5596 6223 5600
rect 6176 5567 6183 5594
rect 6276 5507 6283 5553
rect 6296 5547 6303 5613
rect 6136 5436 6153 5447
rect 6140 5433 6153 5436
rect 6056 5327 6063 5373
rect 6096 5340 6103 5343
rect 6093 5327 6107 5340
rect 6136 5323 6143 5343
rect 6116 5316 6143 5323
rect 6096 5107 6103 5133
rect 6036 5096 6053 5103
rect 6053 5080 6067 5093
rect 6056 5076 6063 5080
rect 6116 5043 6123 5316
rect 6136 5207 6143 5233
rect 6133 5127 6147 5133
rect 6076 5007 6083 5043
rect 6096 5036 6123 5043
rect 5987 4903 6000 4907
rect 5987 4893 6003 4903
rect 5996 4883 6003 4893
rect 5996 4876 6023 4883
rect 5973 4860 5987 4872
rect 5976 4856 5983 4860
rect 6016 4856 6023 4876
rect 6033 4867 6047 4873
rect 5876 4556 5923 4563
rect 5807 4483 5820 4487
rect 5807 4473 5823 4483
rect 5816 4467 5823 4473
rect 5796 4367 5803 4452
rect 5756 4336 5783 4343
rect 5816 4336 5823 4453
rect 5856 4407 5863 4523
rect 5896 4427 5903 4513
rect 5916 4387 5923 4556
rect 5936 4507 5943 4793
rect 5956 4427 5963 4813
rect 6016 4687 6023 4793
rect 6056 4747 6063 4893
rect 6076 4767 6083 4953
rect 6056 4687 6063 4712
rect 5976 4607 5983 4653
rect 6076 4607 6083 4693
rect 6066 4593 6067 4600
rect 6053 4587 6067 4593
rect 6096 4587 6103 5036
rect 6136 5023 6143 5092
rect 6156 5043 6163 5313
rect 6176 5087 6183 5393
rect 6196 5267 6203 5453
rect 6296 5376 6303 5433
rect 6316 5407 6323 5693
rect 6276 5340 6283 5343
rect 6273 5327 6287 5340
rect 6196 5107 6203 5253
rect 6296 5227 6303 5293
rect 6216 5076 6223 5133
rect 6256 5127 6263 5173
rect 6256 5076 6263 5113
rect 6156 5036 6183 5043
rect 6116 5016 6143 5023
rect 6116 4867 6123 5016
rect 6176 5007 6183 5036
rect 6136 4887 6143 4993
rect 6196 4987 6203 5043
rect 6176 4927 6183 4953
rect 6133 4860 6147 4873
rect 6136 4856 6143 4860
rect 6176 4856 6183 4913
rect 6156 4807 6163 4823
rect 6193 4807 6207 4813
rect 6156 4796 6173 4807
rect 6160 4793 6173 4796
rect 6116 4707 6123 4773
rect 6060 4526 6073 4527
rect 6016 4520 6023 4523
rect 6013 4507 6027 4520
rect 6067 4513 6073 4526
rect 6096 4507 6103 4573
rect 6026 4500 6027 4507
rect 5956 4413 5973 4427
rect 5876 4327 5883 4373
rect 5956 4367 5963 4413
rect 5796 4300 5803 4303
rect 5793 4287 5807 4300
rect 5836 4296 5863 4303
rect 5756 4127 5763 4233
rect 5856 4227 5863 4296
rect 5656 4076 5683 4083
rect 5556 3816 5583 3823
rect 5576 3727 5583 3816
rect 5556 3647 5563 3713
rect 5493 3520 5507 3533
rect 5496 3516 5503 3520
rect 5536 3516 5543 3573
rect 5556 3527 5563 3553
rect 5576 3547 5583 3593
rect 5316 3480 5323 3483
rect 5313 3467 5327 3480
rect 5096 3286 5103 3313
rect 5336 3247 5343 3413
rect 5396 3407 5403 3433
rect 5036 3127 5043 3243
rect 5056 3167 5063 3233
rect 5096 3107 5103 3233
rect 5396 3227 5403 3393
rect 5416 3367 5423 3513
rect 5416 3283 5423 3313
rect 5436 3307 5443 3493
rect 5476 3480 5483 3483
rect 5456 3307 5463 3473
rect 5473 3467 5487 3480
rect 5536 3423 5543 3453
rect 5556 3447 5563 3473
rect 5536 3416 5563 3423
rect 5416 3276 5443 3283
rect 5196 3147 5203 3213
rect 4796 2407 4803 2653
rect 4816 2327 4823 2513
rect 4856 2487 4863 2593
rect 4936 2487 4943 2633
rect 4836 2407 4843 2473
rect 4887 2403 4900 2407
rect 4887 2393 4903 2403
rect 4896 2347 4903 2393
rect 4916 2387 4923 2443
rect 4713 2300 4727 2313
rect 4716 2296 4723 2300
rect 4656 2256 4683 2263
rect 4776 2220 4803 2223
rect 4776 2216 4807 2220
rect 4793 2207 4807 2216
rect 4556 1976 4583 1983
rect 4556 1956 4563 1976
rect 4736 1987 4743 2173
rect 4576 1887 4583 1923
rect 4616 1867 4623 1923
rect 4496 1736 4523 1743
rect 4516 1716 4523 1736
rect 4256 1307 4263 1403
rect 4236 1216 4243 1293
rect 4296 1267 4303 1434
rect 4316 1223 4323 1513
rect 4336 1307 4343 1613
rect 4376 1436 4383 1533
rect 4476 1487 4483 1703
rect 4456 1347 4463 1434
rect 4316 1216 4343 1223
rect 4436 1216 4443 1293
rect 4196 1187 4203 1214
rect 4336 1186 4343 1216
rect 4256 1180 4263 1183
rect 4253 1167 4267 1180
rect 4296 1147 4303 1183
rect 4296 1047 4303 1133
rect 4216 1007 4223 1033
rect 4076 747 4083 883
rect 4116 880 4123 883
rect 4113 867 4127 880
rect 4196 867 4203 952
rect 4216 747 4223 993
rect 4236 787 4243 872
rect 4316 767 4323 843
rect 4036 627 4043 693
rect 4176 666 4183 733
rect 4096 660 4103 663
rect 4093 647 4107 660
rect 3756 356 3783 363
rect 3776 327 3783 356
rect 3716 320 3723 323
rect 3713 307 3727 320
rect 3796 187 3803 394
rect 3856 363 3863 433
rect 3856 356 3883 363
rect 3856 176 3863 293
rect 3916 227 3923 313
rect 4036 307 4043 394
rect 4056 366 4063 453
rect 4116 396 4123 573
rect 4036 267 4043 293
rect 3796 146 3803 173
rect 3676 140 3683 143
rect 3716 140 3723 143
rect 3673 127 3687 140
rect 3713 127 3727 140
rect 3916 143 3923 213
rect 4216 176 4223 652
rect 4376 467 4383 1093
rect 4396 867 4403 1073
rect 4476 967 4483 1473
rect 4496 1047 4503 1693
rect 4536 1436 4543 1533
rect 4556 1467 4563 1773
rect 4576 1716 4583 1833
rect 4656 1827 4663 1973
rect 4673 1947 4687 1953
rect 4696 1887 4703 1973
rect 4727 1963 4740 1967
rect 4727 1956 4743 1963
rect 4773 1960 4787 1973
rect 4776 1956 4783 1960
rect 4727 1953 4740 1956
rect 4756 1827 4763 1923
rect 4796 1887 4803 1923
rect 4836 1827 4843 2313
rect 4916 2287 4923 2373
rect 4936 2367 4943 2433
rect 4887 2283 4900 2287
rect 4887 2273 4903 2283
rect 4856 2127 4863 2273
rect 4896 2256 4903 2273
rect 4936 2256 4943 2353
rect 4956 2343 4963 2873
rect 5016 2776 5023 2853
rect 5096 2827 5103 2873
rect 5176 2847 5183 3093
rect 5236 3087 5243 3113
rect 5236 3016 5243 3073
rect 5276 2987 5283 3113
rect 5116 2803 5123 2833
rect 5053 2788 5067 2793
rect 5096 2796 5123 2803
rect 5096 2746 5103 2796
rect 4996 2627 5003 2733
rect 4976 2367 4983 2533
rect 5036 2507 5043 2743
rect 5116 2727 5123 2773
rect 5056 2687 5063 2713
rect 4996 2446 5003 2493
rect 5013 2487 5027 2493
rect 5053 2480 5067 2493
rect 5096 2487 5103 2673
rect 5136 2547 5143 2793
rect 5153 2783 5167 2793
rect 5153 2780 5183 2783
rect 5156 2776 5183 2780
rect 5216 2776 5223 2933
rect 5236 2807 5243 2953
rect 5273 2943 5287 2952
rect 5256 2940 5287 2943
rect 5256 2936 5283 2940
rect 5256 2907 5263 2936
rect 5296 2923 5303 3093
rect 5276 2916 5303 2923
rect 5056 2476 5063 2480
rect 4956 2336 4983 2343
rect 4976 2263 4983 2336
rect 4996 2287 5003 2432
rect 5076 2407 5083 2443
rect 4976 2256 5003 2263
rect 4956 2220 4963 2223
rect 4953 2207 4967 2220
rect 4616 1527 4623 1813
rect 4856 1667 4863 1912
rect 4876 1887 4883 2073
rect 4940 1983 4953 1987
rect 4936 1973 4953 1983
rect 4936 1956 4943 1973
rect 4976 1967 4983 2153
rect 4956 1887 4963 1923
rect 4916 1680 4923 1683
rect 4913 1667 4927 1680
rect 4613 1440 4627 1453
rect 4616 1436 4623 1440
rect 4756 1436 4763 1513
rect 4836 1447 4843 1573
rect 4956 1567 4963 1713
rect 4556 1347 4563 1403
rect 4596 1400 4603 1403
rect 4593 1387 4607 1400
rect 4556 1216 4563 1253
rect 4516 1147 4523 1214
rect 4576 1167 4583 1183
rect 4516 967 4523 1133
rect 4416 827 4423 914
rect 4436 867 4443 953
rect 4533 947 4547 953
rect 4496 867 4503 883
rect 4487 856 4503 867
rect 4487 853 4500 856
rect 4516 787 4523 853
rect 4556 827 4563 872
rect 4396 708 4403 753
rect 4436 666 4443 773
rect 4536 696 4543 733
rect 4576 707 4583 1153
rect 4656 1107 4663 1433
rect 4696 1407 4703 1434
rect 4836 1406 4843 1433
rect 4676 1186 4683 1213
rect 4676 987 4683 1113
rect 4696 1007 4703 1293
rect 4736 1267 4743 1403
rect 4756 1228 4763 1293
rect 4736 1067 4743 1183
rect 4596 823 4603 953
rect 4616 847 4623 933
rect 4756 923 4763 953
rect 4747 916 4763 923
rect 4776 886 4783 993
rect 4596 816 4643 823
rect 4636 803 4643 816
rect 4636 796 4663 803
rect 4476 643 4483 663
rect 4596 647 4603 693
rect 4616 666 4623 733
rect 4636 707 4643 773
rect 4656 723 4663 796
rect 4656 716 4683 723
rect 4676 696 4683 716
rect 4716 696 4723 813
rect 4753 680 4767 693
rect 4756 676 4763 680
rect 4696 660 4703 663
rect 4693 647 4707 660
rect 4476 636 4503 643
rect 4496 567 4503 636
rect 4473 400 4487 413
rect 4496 407 4503 553
rect 4476 396 4483 400
rect 4236 367 4243 394
rect 4356 327 4363 394
rect 4396 367 4403 394
rect 4516 227 4523 413
rect 4596 327 4603 363
rect 4656 307 4663 433
rect 4076 147 4083 174
rect 3876 136 3923 143
rect 4256 146 4263 193
rect 4373 180 4387 193
rect 4376 176 4383 180
rect 4156 107 4163 143
rect 3707 96 3733 103
rect 4296 87 4303 174
rect 4436 146 4443 173
rect 4476 146 4483 213
rect 4616 187 4623 253
rect 4636 146 4643 193
rect 4656 183 4663 213
rect 4676 207 4683 393
rect 4696 366 4703 573
rect 4796 427 4803 1253
rect 4856 1183 4863 1493
rect 4976 1487 4983 1813
rect 4876 1387 4883 1473
rect 4976 1406 4983 1433
rect 4976 1367 4983 1392
rect 4936 1256 4943 1293
rect 4996 1287 5003 2256
rect 5016 2167 5023 2353
rect 5096 2283 5103 2433
rect 5116 2327 5123 2463
rect 5136 2307 5143 2453
rect 5096 2276 5143 2283
rect 5136 2256 5143 2276
rect 5156 2267 5163 2733
rect 5236 2687 5243 2743
rect 5276 2627 5283 2916
rect 5296 2647 5303 2893
rect 5316 2887 5323 3053
rect 5336 2787 5343 3212
rect 5416 3187 5423 3213
rect 5456 3207 5463 3272
rect 5407 3176 5423 3187
rect 5407 3173 5420 3176
rect 5356 3007 5363 3173
rect 5416 3127 5423 3153
rect 5396 3067 5403 3093
rect 5373 3000 5387 3013
rect 5416 3007 5423 3113
rect 5376 2996 5383 3000
rect 5436 2967 5443 3173
rect 5456 3127 5463 3193
rect 5356 2776 5363 2873
rect 5176 2407 5183 2452
rect 5216 2447 5223 2573
rect 5356 2507 5363 2633
rect 5376 2587 5383 2732
rect 5416 2607 5423 2913
rect 5436 2647 5443 2932
rect 5456 2887 5463 3092
rect 5476 3067 5483 3292
rect 5476 2847 5483 3032
rect 5496 3007 5503 3373
rect 5516 3107 5523 3293
rect 5516 2996 5523 3053
rect 5536 3023 5543 3333
rect 5556 3307 5563 3416
rect 5576 3347 5583 3512
rect 5596 3427 5603 3813
rect 5616 3563 5623 3873
rect 5636 3607 5643 3932
rect 5656 3827 5663 4076
rect 5676 3987 5683 4053
rect 5696 3947 5703 3993
rect 5736 3967 5743 4003
rect 5753 3967 5767 3973
rect 5753 3960 5773 3967
rect 5756 3956 5773 3960
rect 5760 3953 5773 3956
rect 5676 3816 5683 3913
rect 5716 3816 5723 3893
rect 5796 3887 5803 4073
rect 5816 3907 5823 4033
rect 5776 3807 5783 3853
rect 5696 3780 5703 3783
rect 5736 3780 5743 3783
rect 5693 3767 5707 3780
rect 5733 3767 5747 3780
rect 5616 3556 5643 3563
rect 5616 3427 5623 3533
rect 5636 3527 5643 3556
rect 5656 3547 5663 3673
rect 5676 3567 5683 3713
rect 5696 3543 5703 3633
rect 5676 3536 5703 3543
rect 5676 3516 5683 3536
rect 5647 3483 5660 3487
rect 5700 3483 5713 3487
rect 5647 3476 5663 3483
rect 5696 3476 5713 3483
rect 5647 3473 5660 3476
rect 5700 3473 5713 3476
rect 5596 3327 5603 3353
rect 5580 3326 5603 3327
rect 5587 3316 5603 3326
rect 5587 3313 5600 3316
rect 5616 3307 5623 3392
rect 5567 3296 5583 3303
rect 5556 3227 5563 3253
rect 5596 3227 5603 3263
rect 5596 3067 5603 3133
rect 5616 3043 5623 3253
rect 5636 3147 5643 3413
rect 5676 3383 5683 3413
rect 5656 3376 5683 3383
rect 5596 3036 5623 3043
rect 5536 3016 5563 3023
rect 5556 2996 5563 3016
rect 5596 3007 5603 3036
rect 5496 2867 5503 2893
rect 5536 2887 5543 2963
rect 5596 2903 5603 2953
rect 5576 2896 5603 2903
rect 5536 2776 5543 2833
rect 5576 2787 5583 2896
rect 5456 2623 5463 2773
rect 5516 2627 5523 2743
rect 5536 2687 5543 2713
rect 5456 2616 5483 2623
rect 5376 2467 5383 2513
rect 5216 2367 5223 2393
rect 5036 2207 5043 2253
rect 5056 2147 5063 2213
rect 5016 1447 5023 2132
rect 5076 2123 5083 2223
rect 5056 2116 5083 2123
rect 5036 1703 5043 2033
rect 5056 1967 5063 2116
rect 5076 2027 5083 2093
rect 5096 2047 5103 2113
rect 5116 2027 5123 2223
rect 5176 2087 5183 2353
rect 5456 2327 5463 2593
rect 5476 2527 5483 2616
rect 5596 2547 5603 2873
rect 5616 2746 5623 3013
rect 5496 2507 5503 2533
rect 5636 2527 5643 3093
rect 5656 2827 5663 3376
rect 5676 3247 5683 3353
rect 5736 3323 5743 3653
rect 5756 3387 5763 3713
rect 5776 3707 5783 3733
rect 5776 3407 5783 3693
rect 5796 3547 5803 3813
rect 5816 3767 5823 3833
rect 5836 3827 5843 4173
rect 5876 4063 5883 4313
rect 5896 4287 5903 4333
rect 5916 4287 5923 4352
rect 5936 4267 5943 4293
rect 5896 4167 5903 4213
rect 5856 4060 5883 4063
rect 5853 4056 5883 4060
rect 5853 4047 5867 4056
rect 5896 4036 5903 4153
rect 5936 4036 5943 4232
rect 5956 4187 5963 4303
rect 5996 4300 6003 4303
rect 5993 4287 6007 4300
rect 6016 4267 6023 4293
rect 5956 4047 5963 4173
rect 5876 3816 5883 3992
rect 5976 3987 5983 4253
rect 6036 4247 6043 4493
rect 6116 4447 6123 4533
rect 6136 4487 6143 4753
rect 6176 4568 6183 4593
rect 6196 4556 6203 4772
rect 6216 4767 6223 4993
rect 6236 4727 6243 5043
rect 6276 4867 6283 4993
rect 6296 4856 6303 5153
rect 6316 4927 6323 5333
rect 6336 5327 6343 5792
rect 6376 5608 6383 5653
rect 6456 5607 6463 5813
rect 6396 5560 6403 5563
rect 6356 5467 6363 5553
rect 6393 5547 6407 5560
rect 6406 5540 6407 5547
rect 6356 5187 6363 5313
rect 6376 5267 6383 5433
rect 6396 5427 6403 5533
rect 6416 5507 6423 5533
rect 6416 5403 6423 5493
rect 6456 5447 6463 5553
rect 6476 5527 6483 5753
rect 6536 5603 6543 6433
rect 6873 6420 6887 6433
rect 6876 6416 6883 6420
rect 6616 6187 6623 6383
rect 6613 6120 6627 6133
rect 6616 6116 6623 6120
rect 6636 6080 6643 6083
rect 6633 6067 6647 6080
rect 6676 6076 6703 6083
rect 6556 5628 6563 5852
rect 6576 5827 6583 5933
rect 6596 5860 6603 5863
rect 6593 5847 6607 5860
rect 6656 5827 6663 5863
rect 6576 5627 6583 5653
rect 6516 5596 6543 5603
rect 6496 5567 6503 5593
rect 6396 5400 6423 5403
rect 6393 5396 6423 5400
rect 6393 5387 6407 5396
rect 6456 5376 6463 5412
rect 6476 5327 6483 5343
rect 6416 5087 6423 5213
rect 6436 5147 6443 5293
rect 6476 5207 6483 5313
rect 6516 5227 6523 5596
rect 6536 5387 6543 5553
rect 6576 5527 6583 5563
rect 6556 5346 6563 5393
rect 6616 5376 6623 5553
rect 6636 5407 6643 5673
rect 6656 5487 6663 5792
rect 6656 5387 6663 5473
rect 6636 5340 6643 5343
rect 6633 5327 6647 5340
rect 6533 5287 6547 5293
rect 6456 5147 6463 5173
rect 6396 5007 6403 5043
rect 6336 4856 6343 4893
rect 6256 4787 6263 4853
rect 6273 4807 6287 4812
rect 6236 4587 6243 4653
rect 6316 4567 6323 4633
rect 5913 3820 5927 3833
rect 5936 3827 5943 3973
rect 5956 3827 5963 3953
rect 5996 3927 6003 4233
rect 6056 4143 6063 4333
rect 6076 4247 6083 4373
rect 6116 4367 6123 4393
rect 6107 4343 6120 4347
rect 6107 4336 6123 4343
rect 6153 4340 6167 4353
rect 6156 4336 6163 4340
rect 6107 4333 6120 4336
rect 6076 4207 6083 4233
rect 6056 4136 6073 4143
rect 6016 4007 6023 4113
rect 6076 4036 6083 4133
rect 6096 4067 6103 4293
rect 6136 4287 6143 4303
rect 6136 4273 6153 4287
rect 6116 4087 6123 4193
rect 6136 4167 6143 4273
rect 5916 3816 5923 3820
rect 5836 3776 5863 3783
rect 5816 3607 5823 3693
rect 5816 3516 5823 3553
rect 5836 3547 5843 3776
rect 5956 3767 5963 3792
rect 5856 3667 5863 3753
rect 5956 3727 5963 3753
rect 5856 3516 5863 3573
rect 5873 3463 5887 3472
rect 5856 3460 5887 3463
rect 5856 3456 5883 3460
rect 5716 3316 5743 3323
rect 5716 3296 5723 3316
rect 5836 3276 5843 3413
rect 5696 3207 5703 3253
rect 5676 2803 5683 3133
rect 5696 3027 5703 3113
rect 5716 3067 5723 3193
rect 5736 3127 5743 3263
rect 5776 3127 5783 3173
rect 5736 3047 5743 3073
rect 5796 3043 5803 3243
rect 5856 3227 5863 3456
rect 5896 3427 5903 3633
rect 5916 3567 5923 3613
rect 5936 3447 5943 3553
rect 5956 3523 5963 3593
rect 5976 3547 5983 3893
rect 6056 3867 6063 3992
rect 6096 3983 6103 4003
rect 6096 3976 6133 3983
rect 6116 3887 6123 3953
rect 5996 3747 6003 3853
rect 6093 3820 6107 3833
rect 6096 3816 6103 3820
rect 6136 3787 6143 3913
rect 6036 3780 6043 3783
rect 6076 3780 6083 3783
rect 6033 3767 6047 3780
rect 6073 3767 6087 3780
rect 5996 3667 6003 3712
rect 6096 3707 6103 3753
rect 6116 3727 6123 3773
rect 6156 3767 6163 4233
rect 6176 4047 6183 4253
rect 6196 4187 6203 4473
rect 6216 4467 6223 4493
rect 6236 4447 6243 4523
rect 6296 4463 6303 4512
rect 6316 4487 6323 4513
rect 6296 4456 6323 4463
rect 6276 4407 6283 4453
rect 6316 4407 6323 4456
rect 6213 4347 6227 4353
rect 6216 4307 6223 4333
rect 6216 4127 6223 4272
rect 6236 4207 6243 4393
rect 6296 4336 6303 4373
rect 6336 4347 6343 4693
rect 6356 4607 6363 4812
rect 6356 4507 6363 4554
rect 6376 4526 6383 4673
rect 6356 4307 6363 4472
rect 6276 4300 6283 4303
rect 6273 4287 6287 4300
rect 6313 4287 6327 4292
rect 6196 4116 6213 4123
rect 6176 3987 6183 4012
rect 6176 3927 6183 3973
rect 6176 3847 6183 3873
rect 6196 3827 6203 4116
rect 6316 4103 6323 4252
rect 6296 4096 6323 4103
rect 6233 4063 6247 4073
rect 6233 4060 6283 4063
rect 6236 4056 6283 4060
rect 6276 4036 6283 4056
rect 6296 4047 6303 4096
rect 6216 3847 6223 3993
rect 6256 3967 6263 4003
rect 6236 3936 6273 3943
rect 6236 3887 6243 3936
rect 6256 3863 6263 3913
rect 6236 3856 6263 3863
rect 6236 3816 6243 3856
rect 6276 3816 6283 3873
rect 6296 3827 6303 3993
rect 6176 3687 6183 3812
rect 6216 3780 6223 3783
rect 6196 3687 6203 3773
rect 6213 3767 6227 3780
rect 6213 3727 6227 3732
rect 6076 3567 6083 3593
rect 5956 3516 5983 3523
rect 6076 3487 6083 3514
rect 6036 3387 6043 3483
rect 6096 3427 6103 3653
rect 6136 3563 6143 3673
rect 6116 3556 6143 3563
rect 6096 3307 6103 3373
rect 6116 3347 6123 3556
rect 6156 3543 6163 3593
rect 6216 3587 6223 3613
rect 6236 3563 6243 3753
rect 6256 3587 6263 3772
rect 6236 3556 6263 3563
rect 6156 3536 6183 3543
rect 6133 3527 6147 3533
rect 6176 3516 6183 3536
rect 6213 3520 6227 3533
rect 6216 3516 6223 3520
rect 6136 3327 6143 3473
rect 5956 3187 5963 3283
rect 6096 3223 6103 3272
rect 6096 3216 6123 3223
rect 5787 3036 5803 3043
rect 5736 2996 5743 3033
rect 5773 3020 5787 3033
rect 5776 3016 5783 3020
rect 5696 2927 5703 2963
rect 5796 2887 5803 2973
rect 5816 2847 5823 2983
rect 5656 2796 5683 2803
rect 5656 2727 5663 2796
rect 5753 2780 5767 2793
rect 5756 2776 5763 2780
rect 5676 2740 5683 2743
rect 5673 2727 5687 2740
rect 5736 2603 5743 2743
rect 5816 2687 5823 2812
rect 5836 2667 5843 3173
rect 6096 3147 6103 3193
rect 5936 3023 5943 3093
rect 6116 3087 6123 3216
rect 6136 3167 6143 3213
rect 6156 3143 6163 3433
rect 6187 3283 6200 3287
rect 6187 3276 6203 3283
rect 6187 3273 6200 3276
rect 6173 3223 6187 3233
rect 6173 3220 6203 3223
rect 6176 3216 6203 3220
rect 6196 3147 6203 3216
rect 6156 3136 6183 3143
rect 6136 3087 6143 3113
rect 5916 3016 5943 3023
rect 5916 2987 5923 3016
rect 6076 2986 6083 3073
rect 6176 3043 6183 3136
rect 6176 3036 6203 3043
rect 5856 2707 5863 2833
rect 5896 2776 5903 2873
rect 5956 2776 5963 2813
rect 5976 2747 5983 2873
rect 6076 2847 6083 2913
rect 6136 2867 6143 3033
rect 6176 2947 6183 2983
rect 6196 2923 6203 3036
rect 6167 2916 6203 2923
rect 6196 2843 6203 2893
rect 6176 2836 6203 2843
rect 5876 2727 5883 2743
rect 5876 2607 5883 2713
rect 5736 2596 5763 2603
rect 5476 2456 5503 2463
rect 5196 2027 5203 2254
rect 5336 2263 5343 2293
rect 5476 2287 5483 2433
rect 5496 2367 5503 2456
rect 5336 2256 5363 2263
rect 5216 2226 5223 2253
rect 5356 2226 5363 2256
rect 5073 1968 5087 1973
rect 5113 1960 5127 1973
rect 5116 1956 5123 1960
rect 5056 1827 5063 1913
rect 5116 1776 5123 1893
rect 5156 1807 5163 1993
rect 5176 1947 5183 1973
rect 5176 1907 5183 1933
rect 5196 1903 5203 2013
rect 5216 1923 5223 1953
rect 5216 1916 5243 1923
rect 5196 1896 5223 1903
rect 5036 1696 5063 1703
rect 5116 1436 5123 1533
rect 5176 1467 5183 1813
rect 5196 1423 5203 1833
rect 5216 1707 5223 1896
rect 5236 1543 5243 1733
rect 5336 1587 5343 1793
rect 5356 1547 5363 2133
rect 5376 2007 5383 2253
rect 5396 1987 5403 2033
rect 5376 1667 5383 1793
rect 5416 1787 5423 2273
rect 5496 2263 5503 2313
rect 5476 2256 5503 2263
rect 5436 2003 5443 2212
rect 5496 2167 5503 2256
rect 5516 2227 5523 2413
rect 5536 2327 5543 2353
rect 5516 2107 5523 2173
rect 5536 2107 5543 2313
rect 5556 2147 5563 2453
rect 5616 2443 5623 2463
rect 5636 2447 5643 2492
rect 5716 2467 5723 2513
rect 5736 2507 5743 2573
rect 5756 2567 5763 2596
rect 5876 2468 5883 2553
rect 5936 2463 5943 2653
rect 5956 2627 5963 2653
rect 6016 2587 6023 2693
rect 5993 2463 6007 2473
rect 5596 2436 5623 2443
rect 5596 2327 5603 2436
rect 5916 2407 5923 2463
rect 5936 2456 5963 2463
rect 5976 2460 6007 2463
rect 5976 2456 6003 2460
rect 5896 2396 5913 2403
rect 5636 2347 5643 2393
rect 5633 2283 5647 2293
rect 5616 2280 5647 2283
rect 5616 2276 5643 2280
rect 5616 2256 5623 2276
rect 5576 2127 5583 2153
rect 5596 2067 5603 2223
rect 5636 2220 5643 2223
rect 5633 2207 5647 2220
rect 5696 2167 5703 2353
rect 5716 2187 5723 2333
rect 5736 2207 5743 2253
rect 5796 2220 5803 2223
rect 5616 2087 5623 2113
rect 5736 2027 5743 2093
rect 5756 2087 5763 2213
rect 5793 2207 5807 2220
rect 5836 2167 5843 2223
rect 5436 2000 5463 2003
rect 5436 1996 5467 2000
rect 5453 1988 5467 1996
rect 5467 1976 5483 1983
rect 5436 1847 5443 1943
rect 5476 1807 5483 1976
rect 5613 1940 5627 1953
rect 5616 1936 5623 1940
rect 5716 1867 5723 1953
rect 5456 1748 5463 1773
rect 5536 1716 5563 1723
rect 5396 1627 5403 1693
rect 5436 1607 5443 1703
rect 5496 1680 5503 1683
rect 5493 1667 5507 1680
rect 5236 1536 5263 1543
rect 5256 1426 5263 1536
rect 5196 1416 5223 1423
rect 5396 1416 5403 1573
rect 5496 1468 5503 1653
rect 5516 1487 5523 1673
rect 5556 1547 5563 1716
rect 5796 1683 5803 1893
rect 5816 1728 5823 2093
rect 5836 1716 5843 2053
rect 5856 1907 5863 2213
rect 5876 2107 5883 2313
rect 5896 2067 5903 2396
rect 5936 2287 5943 2433
rect 5956 2256 5963 2456
rect 5980 2423 5993 2427
rect 5976 2413 5993 2423
rect 5976 2387 5983 2413
rect 5996 2347 6003 2392
rect 6016 2283 6023 2473
rect 6036 2307 6043 2833
rect 6176 2807 6183 2836
rect 6196 2767 6203 2813
rect 6056 2683 6063 2753
rect 6176 2736 6203 2743
rect 6196 2707 6203 2736
rect 6056 2676 6083 2683
rect 6056 2403 6063 2593
rect 6076 2587 6083 2676
rect 6076 2427 6083 2533
rect 6096 2487 6103 2633
rect 6136 2527 6143 2673
rect 6156 2488 6163 2593
rect 6216 2567 6223 3413
rect 6236 3287 6243 3313
rect 6256 3307 6263 3556
rect 6236 3167 6243 3233
rect 6056 2396 6083 2403
rect 6016 2280 6043 2283
rect 6016 2276 6047 2280
rect 6033 2267 6047 2276
rect 5916 2187 5923 2253
rect 5887 2036 5903 2043
rect 5873 2027 5887 2033
rect 5876 1883 5883 1973
rect 5896 1967 5903 2036
rect 5936 1987 5943 2013
rect 5956 1987 5963 2193
rect 5976 2127 5983 2223
rect 5933 1960 5947 1973
rect 5973 1960 5987 1973
rect 5996 1967 6003 2193
rect 6016 2187 6023 2223
rect 6056 2007 6063 2273
rect 6076 2147 6083 2396
rect 6136 2387 6143 2432
rect 6176 2307 6183 2473
rect 6116 2267 6123 2293
rect 6196 2287 6203 2473
rect 6216 2263 6223 2513
rect 6236 2487 6243 3053
rect 6256 2488 6263 3293
rect 6276 3247 6283 3693
rect 6296 3547 6303 3673
rect 6316 3667 6323 4073
rect 6336 3548 6343 4173
rect 6356 4007 6363 4272
rect 6376 4267 6383 4512
rect 6376 4047 6383 4193
rect 6396 4087 6403 4873
rect 6416 4727 6423 5033
rect 6436 4647 6443 5073
rect 6456 5067 6463 5093
rect 6456 4987 6463 5032
rect 6476 4888 6483 5193
rect 6496 5088 6503 5113
rect 6513 5080 6527 5093
rect 6516 5076 6523 5080
rect 6496 4887 6503 5033
rect 6516 4867 6523 4913
rect 6536 4907 6543 5043
rect 6576 5007 6583 5033
rect 6556 4887 6563 4953
rect 6416 4347 6423 4513
rect 6476 4507 6483 4523
rect 6516 4507 6523 4713
rect 6436 4367 6443 4473
rect 6476 4467 6483 4493
rect 6427 4343 6440 4347
rect 6427 4336 6443 4343
rect 6427 4333 6440 4336
rect 6496 4347 6503 4433
rect 6516 4407 6523 4472
rect 6456 4287 6463 4303
rect 6456 4276 6473 4287
rect 6460 4273 6473 4276
rect 6416 4207 6423 4273
rect 6436 4227 6443 4273
rect 6496 4267 6503 4293
rect 6413 4040 6427 4053
rect 6436 4047 6443 4073
rect 6416 4036 6423 4040
rect 6376 3907 6383 3993
rect 6353 3863 6367 3873
rect 6353 3860 6383 3863
rect 6356 3856 6383 3860
rect 6356 3747 6363 3833
rect 6376 3827 6383 3856
rect 6396 3816 6403 3933
rect 6436 3867 6443 3993
rect 6456 3847 6463 4253
rect 6496 4147 6503 4213
rect 6476 3967 6483 4113
rect 6496 4067 6503 4093
rect 6516 4067 6523 4393
rect 6536 4347 6543 4872
rect 6556 4487 6563 4852
rect 6576 4567 6583 4933
rect 6596 4867 6603 5213
rect 6616 5027 6623 5233
rect 6636 4887 6643 5153
rect 6656 5087 6663 5333
rect 6676 5247 6683 6053
rect 6696 5987 6703 6076
rect 6696 5867 6703 5894
rect 6716 5703 6723 6153
rect 6736 6047 6743 6372
rect 6756 6327 6763 6414
rect 6756 6086 6763 6313
rect 6856 6167 6863 6383
rect 6836 6047 6843 6083
rect 6796 5896 6803 6033
rect 6816 5860 6823 5863
rect 6696 5696 6723 5703
rect 6696 5607 6703 5696
rect 6716 5596 6723 5673
rect 6753 5600 6767 5613
rect 6776 5607 6783 5852
rect 6813 5847 6827 5860
rect 6756 5596 6763 5600
rect 6696 5407 6703 5553
rect 6696 5227 6703 5372
rect 6716 5107 6723 5513
rect 6796 5427 6803 5633
rect 6816 5507 6823 5733
rect 6896 5647 6903 6383
rect 6736 5387 6743 5413
rect 6836 5387 6843 5594
rect 6896 5523 6903 5563
rect 6936 5527 6943 5563
rect 6876 5516 6903 5523
rect 6747 5343 6760 5347
rect 6856 5343 6863 5374
rect 6747 5336 6763 5343
rect 6747 5333 6760 5336
rect 6736 5287 6743 5333
rect 6767 5323 6780 5327
rect 6767 5313 6783 5323
rect 6656 5036 6683 5043
rect 6716 5040 6723 5043
rect 6613 4860 6627 4873
rect 6656 4868 6663 5036
rect 6713 5027 6727 5040
rect 6726 5020 6727 5027
rect 6616 4856 6623 4860
rect 6636 4820 6643 4823
rect 6596 4607 6603 4813
rect 6633 4807 6647 4820
rect 6536 4107 6543 4312
rect 6556 4087 6563 4413
rect 6576 4343 6583 4513
rect 6596 4487 6603 4523
rect 6636 4447 6643 4523
rect 6636 4348 6643 4393
rect 6576 4336 6603 4343
rect 6576 4067 6583 4293
rect 6616 4247 6623 4303
rect 6516 4043 6523 4053
rect 6496 4036 6523 4043
rect 6456 3836 6473 3847
rect 6460 3833 6473 3836
rect 6433 3820 6447 3832
rect 6436 3816 6443 3820
rect 6376 3667 6383 3773
rect 6496 3786 6503 4036
rect 6516 3996 6533 4003
rect 6516 3947 6523 3996
rect 6576 3967 6583 4003
rect 6413 3727 6427 3733
rect 6376 3516 6383 3573
rect 6416 3527 6423 3653
rect 6296 3427 6303 3512
rect 6407 3476 6423 3483
rect 6276 2787 6283 3193
rect 6296 2947 6303 3373
rect 6376 3307 6383 3453
rect 6316 3187 6323 3253
rect 6316 3107 6323 3173
rect 6336 3127 6343 3263
rect 6396 3087 6403 3393
rect 6416 3347 6423 3476
rect 6436 3447 6443 3733
rect 6456 3567 6463 3751
rect 6476 3707 6483 3773
rect 6516 3747 6523 3893
rect 6536 3767 6543 3853
rect 6556 3827 6563 3933
rect 6576 3867 6583 3953
rect 6636 3887 6643 4053
rect 6656 4047 6663 4293
rect 6676 4067 6683 4593
rect 6696 4527 6703 4853
rect 6696 4283 6703 4453
rect 6716 4307 6723 4973
rect 6736 4567 6743 5013
rect 6756 4987 6763 5033
rect 6776 5007 6783 5313
rect 6796 5107 6803 5343
rect 6836 5336 6863 5343
rect 6796 4856 6803 5072
rect 6816 5027 6823 5313
rect 6816 4923 6823 4992
rect 6836 4947 6843 5336
rect 6856 5076 6863 5113
rect 6876 5107 6883 5516
rect 6896 5387 6903 5493
rect 6936 5376 6943 5473
rect 6956 5387 6963 5553
rect 6907 5343 6920 5347
rect 6907 5336 6923 5343
rect 6907 5333 6920 5336
rect 6896 5167 6903 5333
rect 6916 5076 6923 5133
rect 6816 4916 6843 4923
rect 6836 4867 6843 4916
rect 6776 4820 6783 4823
rect 6816 4820 6823 4823
rect 6773 4807 6787 4820
rect 6813 4807 6827 4820
rect 6836 4567 6843 4633
rect 6776 4336 6783 4493
rect 6796 4467 6803 4523
rect 6696 4276 6723 4283
rect 6716 4036 6723 4276
rect 6756 4247 6763 4303
rect 6756 4087 6763 4193
rect 6796 4147 6803 4303
rect 6776 4136 6793 4143
rect 6656 4006 6663 4033
rect 6736 3983 6743 4003
rect 6776 3987 6783 4136
rect 6836 4143 6843 4513
rect 6816 4136 6843 4143
rect 6796 4007 6803 4053
rect 6696 3976 6743 3983
rect 6636 3827 6643 3852
rect 6513 3727 6527 3733
rect 6476 3543 6483 3672
rect 6456 3536 6483 3543
rect 6416 3067 6423 3293
rect 6436 3287 6443 3333
rect 6456 3307 6463 3536
rect 6496 3527 6503 3553
rect 6516 3547 6523 3653
rect 6516 3538 6533 3547
rect 6520 3534 6533 3538
rect 6556 3547 6563 3633
rect 6576 3587 6583 3772
rect 6656 3687 6663 3933
rect 6676 3687 6683 3873
rect 6696 3787 6703 3976
rect 6736 3887 6743 3953
rect 6756 3843 6763 3893
rect 6736 3836 6763 3843
rect 6736 3816 6743 3836
rect 6520 3533 6540 3534
rect 6573 3520 6587 3533
rect 6576 3516 6583 3520
rect 6476 3347 6483 3513
rect 6496 3387 6503 3473
rect 6516 3427 6523 3483
rect 6496 3323 6503 3373
rect 6556 3367 6563 3483
rect 6596 3407 6603 3473
rect 6616 3383 6623 3573
rect 6596 3376 6623 3383
rect 6496 3316 6523 3323
rect 6473 3300 6487 3312
rect 6476 3296 6483 3300
rect 6516 3296 6523 3316
rect 6436 3047 6443 3133
rect 6456 3103 6463 3253
rect 6496 3207 6503 3263
rect 6556 3227 6563 3332
rect 6476 3127 6483 3153
rect 6456 3096 6483 3103
rect 6456 3008 6463 3073
rect 6296 2847 6303 2933
rect 6356 2807 6363 2923
rect 6416 2887 6423 2933
rect 6396 2747 6403 2833
rect 6436 2807 6443 2952
rect 6453 2887 6467 2893
rect 6476 2867 6483 3096
rect 6433 2780 6447 2793
rect 6476 2788 6483 2813
rect 6436 2776 6443 2780
rect 6496 2787 6503 3153
rect 6516 2907 6523 3213
rect 6556 3067 6563 3173
rect 6576 3067 6583 3313
rect 6596 3167 6603 3376
rect 6616 3307 6623 3353
rect 6636 3327 6643 3673
rect 6656 3443 6663 3533
rect 6676 3527 6683 3652
rect 6716 3567 6723 3773
rect 6713 3520 6727 3532
rect 6716 3516 6723 3520
rect 6756 3516 6763 3713
rect 6696 3447 6703 3483
rect 6656 3436 6683 3443
rect 6656 3296 6663 3413
rect 6676 3387 6683 3436
rect 6736 3266 6743 3433
rect 6616 3107 6623 3253
rect 6636 3207 6643 3263
rect 6687 3203 6700 3207
rect 6687 3200 6703 3203
rect 6687 3193 6707 3200
rect 6636 3147 6643 3193
rect 6693 3187 6707 3193
rect 6756 3187 6763 3453
rect 6776 3427 6783 3473
rect 6776 3147 6783 3373
rect 6796 3303 6803 3773
rect 6816 3387 6823 4136
rect 6856 4036 6863 5013
rect 6876 4363 6883 4873
rect 6896 4867 6903 5043
rect 6896 4407 6903 4832
rect 6876 4356 6903 4363
rect 6896 4047 6903 4356
rect 6916 4147 6923 4973
rect 6936 4568 6943 5213
rect 6956 5127 6963 5333
rect 6956 4807 6963 5092
rect 6876 4000 6883 4003
rect 6836 3667 6843 3993
rect 6873 3987 6887 4000
rect 6896 3947 6903 3993
rect 6916 3867 6923 4073
rect 6936 3987 6943 4554
rect 6956 3907 6963 4133
rect 6936 3827 6943 3873
rect 6856 3603 6863 3813
rect 6836 3596 6863 3603
rect 6836 3467 6843 3596
rect 6876 3583 6883 3773
rect 6896 3647 6903 3783
rect 6936 3663 6943 3773
rect 6916 3656 6943 3663
rect 6856 3576 6883 3583
rect 6856 3527 6863 3576
rect 6876 3516 6883 3553
rect 6916 3516 6923 3656
rect 6956 3643 6963 3893
rect 6936 3636 6963 3643
rect 6936 3527 6943 3636
rect 6956 3527 6963 3613
rect 6796 3296 6813 3303
rect 6856 3307 6863 3473
rect 6956 3447 6963 3492
rect 6636 2996 6663 3003
rect 6576 2920 6583 2923
rect 6573 2907 6587 2920
rect 6656 2907 6663 2996
rect 6340 2743 6353 2747
rect 6276 2503 6283 2733
rect 6296 2667 6303 2743
rect 6336 2736 6353 2743
rect 6340 2733 6353 2736
rect 6376 2707 6383 2733
rect 6296 2627 6303 2653
rect 6276 2496 6303 2503
rect 6296 2476 6303 2496
rect 6336 2487 6343 2653
rect 6216 2256 6243 2263
rect 6096 2167 6103 2253
rect 6116 2027 6123 2133
rect 6136 2067 6143 2093
rect 6156 2087 6163 2223
rect 6196 2220 6203 2223
rect 6193 2207 6207 2220
rect 5936 1956 5943 1960
rect 5976 1956 5983 1960
rect 5916 1920 5923 1923
rect 5913 1907 5927 1920
rect 5856 1876 5883 1883
rect 5856 1687 5863 1876
rect 5956 1867 5963 1923
rect 5796 1676 5823 1683
rect 5656 1607 5663 1673
rect 5593 1547 5607 1553
rect 5556 1456 5563 1533
rect 5496 1423 5503 1454
rect 5496 1416 5523 1423
rect 5016 1387 5023 1412
rect 5056 1327 5063 1403
rect 5096 1400 5103 1403
rect 5093 1387 5107 1400
rect 4856 1176 4883 1183
rect 4856 987 4863 1176
rect 4916 916 4923 1033
rect 4816 847 4823 914
rect 4816 676 4823 793
rect 4796 396 4803 413
rect 4856 408 4863 813
rect 4896 787 4903 883
rect 5016 827 5023 1313
rect 5056 916 5063 1273
rect 5076 1223 5083 1353
rect 5076 1216 5103 1223
rect 5136 1216 5143 1253
rect 5116 1107 5123 1183
rect 5196 923 5203 1053
rect 5176 916 5203 923
rect 5196 807 5203 916
rect 5236 827 5243 1393
rect 5596 1307 5603 1473
rect 5636 1387 5643 1533
rect 5656 1387 5663 1553
rect 5716 1436 5723 1493
rect 5696 1400 5703 1403
rect 5693 1387 5707 1400
rect 5796 1387 5803 1423
rect 5816 1307 5823 1676
rect 5916 1448 5923 1733
rect 5956 1587 5963 1773
rect 6016 1747 6023 1993
rect 6060 1986 6080 1987
rect 6036 1736 6043 1973
rect 6067 1983 6080 1986
rect 6067 1980 6083 1983
rect 6067 1973 6087 1980
rect 6056 1787 6063 1972
rect 6073 1967 6087 1973
rect 6116 1956 6123 2013
rect 6156 1956 6163 1993
rect 6096 1763 6103 1912
rect 6136 1767 6143 1923
rect 6176 1827 6183 1893
rect 6096 1756 6123 1763
rect 6116 1743 6123 1756
rect 6116 1736 6143 1743
rect 5996 1667 6003 1713
rect 6096 1700 6103 1703
rect 6093 1687 6107 1700
rect 6107 1676 6123 1683
rect 5956 1547 5963 1573
rect 6096 1420 6103 1423
rect 5456 1216 5463 1293
rect 5336 1207 5343 1213
rect 5336 1194 5353 1207
rect 5336 1193 5360 1194
rect 5316 916 5323 973
rect 5336 943 5343 1193
rect 5376 1127 5383 1214
rect 5536 1196 5563 1203
rect 5436 1147 5443 1183
rect 5536 1067 5543 1196
rect 5596 1187 5603 1253
rect 5736 1200 5743 1203
rect 5733 1187 5747 1200
rect 5836 1196 5863 1203
rect 5336 936 5363 943
rect 5356 916 5363 936
rect 5096 707 5103 773
rect 5096 676 5123 683
rect 5096 527 5103 676
rect 5156 640 5163 643
rect 5153 627 5167 640
rect 5087 516 5103 527
rect 5087 513 5100 516
rect 4656 176 4683 183
rect 4713 180 4727 193
rect 4716 176 4723 180
rect 4396 107 4403 143
rect 4776 107 4783 363
rect 4796 146 4803 173
rect 4816 143 4823 293
rect 4876 287 4883 453
rect 4913 400 4927 413
rect 4916 396 4923 400
rect 4936 307 4943 363
rect 4816 136 4853 143
rect 4873 107 4887 113
rect 4867 100 4887 107
rect 4867 96 4883 100
rect 4867 93 4880 96
rect 4896 47 4903 143
rect 4936 127 4943 213
rect 5016 188 5023 493
rect 5036 366 5043 393
rect 5056 307 5063 433
rect 5196 383 5203 793
rect 5236 727 5243 773
rect 5236 666 5243 713
rect 5316 696 5323 853
rect 5336 807 5343 883
rect 5396 867 5403 914
rect 5416 887 5423 953
rect 5476 928 5483 993
rect 5513 920 5527 933
rect 5516 916 5523 920
rect 5416 747 5423 833
rect 5536 807 5543 883
rect 5576 823 5583 1033
rect 5593 927 5607 933
rect 5756 916 5783 923
rect 5556 816 5583 823
rect 5496 696 5503 773
rect 5256 547 5263 694
rect 5296 547 5303 663
rect 5156 380 5163 383
rect 5153 367 5167 380
rect 5196 376 5223 383
rect 5216 247 5223 376
rect 5256 367 5263 533
rect 5556 447 5563 816
rect 5596 803 5603 913
rect 5776 887 5783 916
rect 5636 876 5663 883
rect 5636 807 5643 876
rect 5796 823 5803 1053
rect 5836 1047 5843 1196
rect 5956 1187 5963 1293
rect 6056 1216 6063 1293
rect 6076 1227 6083 1413
rect 6093 1407 6107 1420
rect 6096 1243 6103 1273
rect 6116 1267 6123 1676
rect 6136 1487 6143 1736
rect 6196 1743 6203 2033
rect 6216 1767 6223 2213
rect 6236 2107 6243 2256
rect 6256 2127 6263 2273
rect 6276 2207 6283 2333
rect 6296 2267 6303 2413
rect 6316 2307 6323 2443
rect 6336 2287 6343 2393
rect 6356 2347 6363 2473
rect 6376 2327 6383 2553
rect 6396 2427 6403 2613
rect 6416 2487 6423 2673
rect 6456 2527 6463 2743
rect 6476 2503 6483 2553
rect 6456 2496 6483 2503
rect 6456 2476 6463 2496
rect 6496 2476 6503 2713
rect 6516 2647 6523 2893
rect 6536 2547 6543 2773
rect 6596 2740 6603 2743
rect 6593 2727 6607 2740
rect 6636 2707 6643 2743
rect 6516 2487 6523 2513
rect 6596 2507 6603 2573
rect 6536 2447 6543 2493
rect 6593 2487 6607 2493
rect 6616 2488 6623 2633
rect 6676 2507 6683 3053
rect 6436 2427 6443 2432
rect 6556 2427 6563 2473
rect 6436 2416 6453 2427
rect 6440 2413 6453 2416
rect 6380 2283 6393 2287
rect 6376 2273 6393 2283
rect 6336 2256 6343 2273
rect 6376 2256 6383 2273
rect 6236 1926 6243 2093
rect 6296 2067 6303 2213
rect 6256 1887 6263 2053
rect 6316 2047 6323 2223
rect 6356 2220 6363 2223
rect 6353 2207 6367 2220
rect 6336 1880 6343 1883
rect 6176 1736 6203 1743
rect 6236 1736 6243 1793
rect 6156 1567 6163 1734
rect 6096 1236 6123 1243
rect 6116 1216 6123 1236
rect 6027 1183 6040 1187
rect 6027 1176 6043 1183
rect 6027 1173 6040 1176
rect 5816 847 5823 913
rect 5787 816 5803 823
rect 5576 796 5603 803
rect 5576 667 5583 796
rect 5616 527 5623 663
rect 5676 646 5683 733
rect 5776 708 5783 813
rect 5836 747 5843 953
rect 5876 916 5883 993
rect 5896 967 5903 1163
rect 5956 1147 5963 1173
rect 5916 916 5923 973
rect 6056 916 6063 973
rect 6036 847 6043 883
rect 6096 807 6103 1033
rect 6116 886 6123 973
rect 6136 807 6143 1393
rect 6156 928 6163 1253
rect 6176 1047 6183 1736
rect 6196 1147 6203 1693
rect 6216 1667 6223 1703
rect 6256 1507 6263 1703
rect 6296 1507 6303 1873
rect 6333 1867 6347 1880
rect 6396 1847 6403 2013
rect 6416 1943 6423 2313
rect 6436 2067 6443 2273
rect 6456 2027 6463 2373
rect 6493 2268 6507 2273
rect 6536 2256 6543 2293
rect 6416 1936 6443 1943
rect 6416 1887 6423 1913
rect 6316 1706 6323 1753
rect 6196 987 6203 1133
rect 6216 1087 6223 1473
rect 6296 1436 6303 1493
rect 6336 1468 6343 1832
rect 6373 1740 6387 1753
rect 6416 1748 6423 1852
rect 6436 1827 6443 1936
rect 6456 1907 6463 1992
rect 6476 1968 6483 2093
rect 6516 1956 6523 2133
rect 6536 2007 6543 2053
rect 6576 2027 6583 2474
rect 6653 2480 6667 2493
rect 6696 2487 6703 3133
rect 6836 3127 6843 3263
rect 6796 3027 6803 3073
rect 6793 3000 6807 3013
rect 6836 3007 6843 3073
rect 6796 2996 6803 3000
rect 6716 2947 6723 2994
rect 6656 2476 6663 2480
rect 6676 2407 6683 2443
rect 6696 2387 6703 2433
rect 6596 2227 6603 2353
rect 6716 2347 6723 2853
rect 6756 2776 6763 2933
rect 6776 2907 6783 2963
rect 6856 2966 6863 3033
rect 6836 2787 6843 2953
rect 6736 2447 6743 2693
rect 6776 2647 6783 2732
rect 6816 2707 6823 2743
rect 6836 2627 6843 2733
rect 6756 2367 6763 2513
rect 6793 2480 6807 2493
rect 6796 2476 6803 2480
rect 6836 2476 6843 2513
rect 6856 2507 6863 2952
rect 6876 2687 6883 3373
rect 6896 2467 6903 3093
rect 6916 3087 6923 3293
rect 6916 2567 6923 3013
rect 6956 2667 6963 3433
rect 6560 1963 6573 1967
rect 6556 1956 6573 1963
rect 6560 1953 6573 1956
rect 6496 1920 6503 1923
rect 6493 1907 6507 1920
rect 6536 1887 6543 1923
rect 6476 1847 6483 1873
rect 6556 1827 6563 1893
rect 6436 1767 6443 1813
rect 6376 1736 6383 1740
rect 6476 1706 6483 1793
rect 6396 1700 6403 1703
rect 6356 1467 6363 1693
rect 6393 1687 6407 1700
rect 6496 1687 6503 1813
rect 6596 1807 6603 2113
rect 6616 2047 6623 2333
rect 6756 2267 6763 2293
rect 6756 2107 6763 2253
rect 6736 2047 6743 2073
rect 6776 2047 6783 2393
rect 6273 1260 6287 1273
rect 6316 1267 6323 1403
rect 6356 1367 6363 1403
rect 6396 1367 6403 1453
rect 6376 1356 6393 1363
rect 6276 1256 6283 1260
rect 6296 967 6303 1033
rect 5876 708 5883 733
rect 5916 676 5923 793
rect 6176 707 6183 793
rect 6216 723 6223 843
rect 6196 716 6223 723
rect 6036 680 6043 683
rect 6033 667 6047 680
rect 5396 376 5403 433
rect 5496 327 5503 433
rect 5556 416 5563 433
rect 5676 428 5683 632
rect 5756 607 5763 663
rect 5816 507 5823 663
rect 6176 627 6183 693
rect 6196 687 6203 716
rect 6213 680 6227 693
rect 6216 676 6223 680
rect 5676 386 5683 414
rect 5656 327 5663 383
rect 5776 376 5783 493
rect 6036 383 6043 513
rect 5256 216 5263 313
rect 5056 176 5063 213
rect 5296 176 5323 183
rect 5036 47 5043 143
rect 5176 143 5183 173
rect 5316 163 5323 176
rect 5316 160 5343 163
rect 5313 156 5343 160
rect 5396 156 5403 233
rect 5313 147 5327 156
rect 5176 136 5203 143
rect 5576 107 5583 163
rect 5676 127 5683 372
rect 5876 176 5883 253
rect 5956 247 5963 383
rect 6016 376 6043 383
rect 6116 367 6123 533
rect 6236 487 6243 713
rect 6276 676 6283 853
rect 6173 400 6187 413
rect 6176 396 6183 400
rect 6216 396 6223 433
rect 6236 427 6243 473
rect 6156 360 6163 363
rect 6153 347 6167 360
rect 5996 156 6023 163
rect 5836 87 5843 153
rect 5916 140 5923 143
rect 5913 126 5927 140
rect 6016 87 6023 156
rect 6256 127 6263 393
rect 6276 243 6283 613
rect 6296 527 6303 913
rect 6316 607 6323 893
rect 6296 347 6303 413
rect 6316 408 6323 593
rect 6336 507 6343 993
rect 6356 886 6363 953
rect 6376 927 6383 1356
rect 6396 987 6403 1253
rect 6416 1007 6423 1433
rect 6436 1406 6443 1453
rect 6496 1436 6503 1473
rect 6516 1447 6523 1793
rect 6533 1743 6547 1753
rect 6533 1740 6563 1743
rect 6536 1736 6563 1740
rect 6576 1700 6583 1703
rect 6573 1687 6587 1700
rect 6616 1647 6623 2012
rect 6667 1963 6680 1967
rect 6736 1963 6743 2033
rect 6667 1956 6683 1963
rect 6736 1956 6763 1963
rect 6667 1953 6680 1956
rect 6656 1907 6663 1953
rect 6636 1687 6643 1833
rect 6656 1706 6663 1773
rect 6756 1768 6763 1956
rect 6776 1767 6783 1993
rect 6796 1706 6803 2353
rect 6896 2227 6903 2432
rect 6916 2307 6923 2553
rect 6936 2243 6943 2453
rect 6916 2236 6943 2243
rect 6916 2127 6923 2236
rect 6856 1956 6863 2033
rect 6816 1923 6823 1954
rect 6816 1916 6833 1923
rect 6456 1216 6463 1253
rect 6536 1127 6543 1633
rect 6656 1587 6663 1692
rect 6556 1267 6563 1433
rect 6576 1406 6583 1573
rect 6676 1448 6683 1693
rect 6816 1607 6823 1753
rect 6836 1747 6843 1912
rect 6876 1887 6883 1923
rect 6893 1740 6907 1753
rect 6936 1748 6943 2213
rect 6896 1736 6903 1740
rect 6956 1747 6963 2653
rect 6836 1687 6843 1733
rect 6867 1703 6880 1707
rect 6867 1696 6883 1703
rect 6867 1693 6880 1696
rect 6556 1187 6563 1214
rect 6416 916 6423 993
rect 6336 396 6343 433
rect 6356 427 6363 872
rect 6456 727 6463 953
rect 6516 883 6523 1053
rect 6576 967 6583 1392
rect 6616 1327 6623 1403
rect 6656 1247 6663 1333
rect 6633 1220 6647 1233
rect 6636 1216 6643 1220
rect 6676 1207 6683 1253
rect 6696 1247 6703 1593
rect 6716 1407 6723 1553
rect 6776 1436 6783 1473
rect 6856 1327 6863 1693
rect 6876 1303 6883 1673
rect 6856 1296 6883 1303
rect 6696 1186 6703 1233
rect 6716 1147 6723 1214
rect 6856 1183 6863 1296
rect 6836 1176 6863 1183
rect 6516 876 6543 883
rect 6576 708 6583 843
rect 6656 696 6663 933
rect 6676 887 6683 1113
rect 6836 1107 6843 1176
rect 6396 656 6423 663
rect 6396 547 6403 656
rect 6576 647 6583 694
rect 6356 307 6363 363
rect 6376 267 6383 333
rect 6276 236 6293 243
rect 6296 156 6303 233
rect 6356 156 6363 213
rect 6396 167 6403 363
rect 6436 307 6443 393
rect 6416 147 6423 173
rect 6456 87 6463 513
rect 6476 227 6483 493
rect 6496 367 6503 433
rect 6576 396 6583 533
rect 6636 408 6643 663
rect 6676 660 6683 663
rect 6673 647 6687 660
rect 6716 627 6723 1093
rect 6756 916 6763 973
rect 6793 920 6807 933
rect 6796 916 6803 920
rect 6816 847 6823 883
rect 6816 696 6823 833
rect 6796 547 6803 663
rect 6696 396 6703 533
rect 6556 327 6563 363
rect 6636 327 6643 394
rect 6556 188 6563 253
rect 6716 216 6723 313
rect 6776 207 6783 433
rect 6796 143 6803 473
rect 6816 287 6823 613
rect 6856 396 6863 1073
rect 6876 847 6883 1213
rect 6896 447 6903 1573
rect 6916 423 6923 1692
rect 6936 1347 6943 1673
rect 6896 416 6923 423
rect 6896 396 6903 416
rect 6536 140 6543 143
rect 6533 127 6547 140
rect 6776 136 6803 143
rect 6836 127 6843 193
rect 6876 183 6883 363
rect 6916 327 6923 363
rect 6956 327 6963 1693
rect 6856 176 6883 183
rect 6916 176 6923 273
rect 6856 146 6863 176
rect 6896 140 6903 143
rect 6893 127 6907 140
rect 1116 -24 1143 -17
rect 1296 -24 1323 -17
rect 1596 -24 1623 -17
<< m3contact >>
rect 293 6513 307 6527
rect 333 6513 347 6527
rect 153 6414 167 6428
rect 273 6414 287 6428
rect 113 6372 127 6386
rect 433 6433 447 6447
rect 413 6414 427 6428
rect 353 6313 367 6327
rect 13 6113 27 6127
rect 173 6114 187 6128
rect 13 6072 27 6086
rect 133 6072 147 6086
rect 153 5894 167 5908
rect 253 6114 267 6128
rect 253 6072 267 6086
rect 313 6072 327 6086
rect 2713 6453 2727 6467
rect 2973 6453 2987 6467
rect 3013 6453 3027 6467
rect 3153 6453 3167 6467
rect 3273 6453 3287 6467
rect 4133 6453 4147 6467
rect 4213 6453 4227 6467
rect 4433 6453 4447 6467
rect 4913 6453 4927 6467
rect 4953 6453 4967 6467
rect 5113 6453 5127 6467
rect 6333 6453 6347 6467
rect 6453 6453 6467 6467
rect 2393 6433 2407 6447
rect 2493 6433 2507 6447
rect 813 6413 827 6427
rect 913 6413 927 6427
rect 493 6393 507 6407
rect 473 6372 487 6386
rect 473 6333 487 6347
rect 573 6313 587 6327
rect 573 6273 587 6287
rect 673 6233 687 6247
rect 713 6233 727 6247
rect 533 6114 547 6128
rect 653 6114 667 6128
rect 1373 6413 1387 6427
rect 1733 6413 1747 6427
rect 933 6393 947 6407
rect 1013 6394 1027 6408
rect 873 6333 887 6347
rect 913 6333 927 6347
rect 813 6213 827 6227
rect 833 6133 847 6147
rect 893 6133 907 6147
rect 793 6114 807 6128
rect 413 6053 427 6067
rect 493 6053 507 6067
rect 253 5894 267 5908
rect 113 5832 127 5846
rect 193 5832 207 5846
rect 53 5713 67 5727
rect 193 5713 207 5727
rect 113 5594 127 5608
rect 153 5493 167 5507
rect 353 5773 367 5787
rect 353 5613 367 5627
rect 533 5973 547 5987
rect 593 5874 607 5888
rect 593 5572 607 5586
rect 513 5493 527 5507
rect 253 5473 267 5487
rect 393 5473 407 5487
rect 233 5453 247 5467
rect 333 5453 347 5467
rect 13 5353 27 5367
rect 53 5353 67 5367
rect 12 5313 26 5327
rect 33 5312 47 5326
rect 13 5273 27 5287
rect 53 5273 67 5287
rect 33 4673 47 4687
rect 13 4293 27 4307
rect 13 3913 27 3927
rect 193 5293 207 5307
rect 373 5354 387 5368
rect 473 5413 487 5427
rect 393 5273 407 5287
rect 433 5273 447 5287
rect 253 5193 267 5207
rect 333 5193 347 5207
rect 113 5074 127 5088
rect 173 5074 187 5088
rect 153 5032 167 5046
rect 233 4993 247 5007
rect 113 4812 127 4826
rect 73 4753 87 4767
rect 193 4673 207 4687
rect 233 4593 247 4607
rect 113 4554 127 4568
rect 353 5113 367 5127
rect 293 5074 307 5088
rect 333 4993 347 5007
rect 273 4854 287 4868
rect 313 4673 327 4687
rect 333 4593 347 4607
rect 393 4993 407 5007
rect 493 5354 507 5368
rect 473 5293 487 5307
rect 453 5153 467 5167
rect 433 4854 447 4868
rect 713 6073 727 6087
rect 813 6072 827 6086
rect 893 5993 907 6007
rect 973 6273 987 6287
rect 933 6213 947 6227
rect 973 6193 987 6207
rect 1073 6193 1087 6207
rect 1013 6153 1027 6167
rect 933 6114 947 6128
rect 973 6114 987 6128
rect 1333 6394 1347 6408
rect 1333 6333 1347 6347
rect 1373 6333 1387 6347
rect 1233 6173 1247 6187
rect 1133 6133 1147 6147
rect 993 6072 1007 6086
rect 1053 6053 1067 6067
rect 933 6033 947 6047
rect 993 6033 1007 6047
rect 1033 6033 1047 6047
rect 913 5973 927 5987
rect 853 5953 867 5967
rect 773 5894 787 5908
rect 933 5894 947 5908
rect 673 5853 687 5867
rect 733 5852 747 5866
rect 673 5773 687 5787
rect 633 5473 647 5487
rect 593 5413 607 5427
rect 533 5393 547 5407
rect 533 5332 547 5346
rect 573 5332 587 5346
rect 613 5332 627 5346
rect 613 5113 627 5127
rect 553 5074 567 5088
rect 813 5853 827 5867
rect 753 5613 767 5627
rect 793 5613 807 5627
rect 773 5552 787 5566
rect 733 5513 747 5527
rect 693 5373 707 5387
rect 773 5433 787 5447
rect 753 5393 767 5407
rect 993 5813 1007 5827
rect 1093 6033 1107 6047
rect 1052 5993 1066 6007
rect 1073 5993 1087 6007
rect 1073 5953 1087 5967
rect 1433 6273 1447 6287
rect 1433 6213 1447 6227
rect 1513 6173 1527 6187
rect 1493 6153 1507 6167
rect 1433 6133 1447 6147
rect 1373 6033 1387 6047
rect 1413 6033 1427 6047
rect 1113 5953 1127 5967
rect 1193 5953 1207 5967
rect 1073 5852 1087 5866
rect 1093 5813 1107 5827
rect 1033 5773 1047 5787
rect 1093 5773 1107 5787
rect 973 5713 987 5727
rect 953 5673 967 5687
rect 833 5593 847 5607
rect 913 5594 927 5608
rect 833 5552 847 5566
rect 893 5552 907 5566
rect 933 5552 947 5566
rect 853 5513 867 5527
rect 893 5513 907 5527
rect 873 5493 887 5507
rect 853 5433 867 5447
rect 693 5332 707 5346
rect 693 5133 707 5147
rect 653 5032 667 5046
rect 693 5032 707 5046
rect 653 4993 667 5007
rect 493 4793 507 4807
rect 473 4773 487 4787
rect 613 4793 627 4807
rect 653 4793 667 4807
rect 593 4753 607 4767
rect 553 4653 567 4667
rect 493 4593 507 4607
rect 353 4553 367 4567
rect 153 4512 167 4526
rect 213 4512 227 4526
rect 113 4334 127 4348
rect 153 4334 167 4348
rect 193 4334 207 4348
rect 73 4293 87 4307
rect 133 4292 147 4306
rect 173 4093 187 4107
rect 113 4034 127 4048
rect 133 3814 147 3828
rect 233 4493 247 4507
rect 253 4433 267 4447
rect 373 4433 387 4447
rect 233 4393 247 4407
rect 313 4393 327 4407
rect 273 4334 287 4348
rect 253 4292 267 4306
rect 293 4292 307 4306
rect 233 4253 247 4267
rect 213 4093 227 4107
rect 333 4253 347 4267
rect 533 4513 547 4527
rect 493 4333 507 4347
rect 473 4292 487 4306
rect 533 4293 547 4307
rect 433 4253 447 4267
rect 633 4773 647 4787
rect 613 4513 627 4527
rect 593 4473 607 4487
rect 793 5374 807 5388
rect 733 5333 747 5347
rect 813 5332 827 5346
rect 933 5433 947 5447
rect 933 5374 947 5388
rect 1013 5633 1027 5647
rect 993 5613 1007 5627
rect 1053 5594 1067 5608
rect 1133 5713 1147 5727
rect 1173 5693 1187 5707
rect 1153 5633 1167 5647
rect 1153 5594 1167 5608
rect 993 5553 1007 5567
rect 973 5373 987 5387
rect 873 5353 887 5367
rect 1033 5552 1047 5566
rect 1053 5473 1067 5487
rect 1113 5552 1127 5566
rect 1253 5594 1267 5608
rect 1473 6092 1487 6106
rect 1473 6033 1487 6047
rect 1473 5953 1487 5967
rect 1433 5813 1447 5827
rect 1313 5773 1327 5787
rect 1293 5593 1307 5607
rect 1173 5552 1187 5566
rect 1273 5552 1287 5566
rect 1513 6073 1527 6087
rect 1773 6394 1787 6408
rect 1853 6273 1867 6287
rect 1793 6253 1807 6267
rect 1733 6193 1747 6207
rect 1633 6133 1647 6147
rect 1713 6133 1727 6147
rect 1653 6072 1667 6086
rect 2033 6393 2047 6407
rect 2093 6273 2107 6287
rect 2193 6273 2207 6287
rect 1893 6213 1907 6227
rect 1833 6153 1847 6167
rect 1993 6153 2007 6167
rect 1793 6114 1807 6128
rect 2033 6133 2047 6147
rect 1733 6073 1747 6087
rect 1813 6072 1827 6086
rect 1853 6072 1867 6086
rect 1973 6072 1987 6086
rect 2013 6072 2027 6086
rect 1713 6013 1727 6027
rect 1613 5993 1627 6007
rect 1573 5973 1587 5987
rect 1713 5973 1727 5987
rect 1673 5933 1687 5947
rect 1613 5894 1627 5908
rect 1673 5894 1687 5908
rect 1773 5893 1787 5907
rect 1893 5894 1907 5908
rect 1613 5853 1627 5867
rect 1493 5733 1507 5747
rect 1413 5633 1427 5647
rect 1333 5593 1347 5607
rect 1453 5594 1467 5608
rect 1333 5552 1347 5566
rect 1313 5533 1327 5547
rect 1233 5513 1247 5527
rect 1333 5493 1347 5507
rect 1153 5473 1167 5487
rect 1293 5473 1307 5487
rect 1033 5413 1047 5427
rect 1033 5373 1047 5387
rect 773 5213 787 5227
rect 893 5313 907 5327
rect 813 5193 827 5207
rect 873 5133 887 5147
rect 733 5093 747 5107
rect 713 5013 727 5027
rect 753 5074 767 5088
rect 813 5074 827 5088
rect 833 5032 847 5046
rect 773 4993 787 5007
rect 753 4913 767 4927
rect 993 5312 1007 5326
rect 1013 5293 1027 5307
rect 953 5273 967 5287
rect 913 5213 927 5227
rect 893 5113 907 5127
rect 893 5032 907 5046
rect 833 4854 847 4868
rect 713 4793 727 4807
rect 753 4793 767 4807
rect 693 4713 707 4727
rect 753 4554 767 4568
rect 653 4512 667 4526
rect 733 4512 747 4526
rect 773 4512 787 4526
rect 933 5093 947 5107
rect 1133 5353 1147 5367
rect 1133 5293 1147 5307
rect 1053 5273 1067 5287
rect 1053 5233 1067 5247
rect 1433 5533 1447 5547
rect 1393 5413 1407 5427
rect 1433 5373 1447 5387
rect 1293 5233 1307 5247
rect 1073 5193 1087 5207
rect 1153 5193 1167 5207
rect 1233 5193 1247 5207
rect 1093 5153 1107 5167
rect 1073 5073 1087 5087
rect 1013 5032 1027 5046
rect 1053 5032 1067 5046
rect 993 5013 1007 5027
rect 973 4993 987 5007
rect 913 4873 927 4887
rect 893 4854 907 4868
rect 933 4854 947 4868
rect 973 4854 987 4868
rect 913 4812 927 4826
rect 913 4753 927 4767
rect 973 4753 987 4767
rect 913 4593 927 4607
rect 853 4573 867 4587
rect 953 4573 967 4587
rect 853 4512 867 4526
rect 933 4512 947 4526
rect 893 4493 907 4507
rect 833 4473 847 4487
rect 1013 4953 1027 4967
rect 1153 5074 1167 5088
rect 1093 5033 1107 5047
rect 1133 5032 1147 5046
rect 1093 4854 1107 4868
rect 1133 4853 1147 4867
rect 1293 5093 1307 5107
rect 1333 5074 1347 5088
rect 1373 5074 1387 5088
rect 1233 4993 1247 5007
rect 1373 5033 1387 5047
rect 1313 4993 1327 5007
rect 1653 5853 1667 5867
rect 1993 5953 2007 5967
rect 1633 5693 1647 5707
rect 1593 5594 1607 5608
rect 1573 5552 1587 5566
rect 1633 5552 1647 5566
rect 1533 5533 1547 5547
rect 1553 5513 1567 5527
rect 1553 5473 1567 5487
rect 1573 5453 1587 5467
rect 1533 5433 1547 5447
rect 1533 5374 1547 5388
rect 1493 5233 1507 5247
rect 1453 5193 1467 5207
rect 1433 5093 1447 5107
rect 1413 5073 1427 5087
rect 1453 5074 1467 5088
rect 1593 5313 1607 5327
rect 1733 5852 1747 5866
rect 1773 5852 1787 5866
rect 1873 5733 1887 5747
rect 1973 5853 1987 5867
rect 1953 5753 1967 5767
rect 1913 5713 1927 5727
rect 1813 5673 1827 5687
rect 1773 5653 1787 5667
rect 1693 5613 1707 5627
rect 1673 5594 1687 5608
rect 1733 5594 1747 5608
rect 1913 5633 1927 5647
rect 1853 5613 1867 5627
rect 1833 5594 1847 5608
rect 1753 5552 1767 5566
rect 1813 5552 1827 5566
rect 1913 5594 1927 5608
rect 1853 5553 1867 5567
rect 1893 5552 1907 5566
rect 1933 5552 1947 5566
rect 2213 6213 2227 6227
rect 2193 6193 2207 6207
rect 2173 6114 2187 6128
rect 2153 6013 2167 6027
rect 2033 5894 2047 5908
rect 2092 5894 2106 5908
rect 2113 5894 2127 5908
rect 2173 5894 2187 5908
rect 2313 6313 2327 6327
rect 2293 6173 2307 6187
rect 2273 6153 2287 6167
rect 2273 6114 2287 6128
rect 2253 5953 2267 5967
rect 2013 5853 2027 5867
rect 1713 5513 1727 5527
rect 1673 5374 1687 5388
rect 1733 5374 1747 5388
rect 1633 5153 1647 5167
rect 1553 5113 1567 5127
rect 1553 5074 1567 5088
rect 1753 5332 1767 5346
rect 1713 5313 1727 5327
rect 1733 5293 1747 5307
rect 1713 5074 1727 5088
rect 1473 5032 1487 5046
rect 1273 4953 1287 4967
rect 1393 4953 1407 4967
rect 1493 4953 1507 4967
rect 1473 4933 1487 4947
rect 1213 4913 1227 4927
rect 1013 4554 1027 4568
rect 1093 4793 1107 4807
rect 1073 4713 1087 4727
rect 1173 4793 1187 4807
rect 1153 4773 1167 4787
rect 1113 4693 1127 4707
rect 1093 4573 1107 4587
rect 1073 4554 1087 4568
rect 1193 4593 1207 4607
rect 1033 4513 1047 4527
rect 1093 4512 1107 4526
rect 1073 4493 1087 4507
rect 993 4433 1007 4447
rect 573 4333 587 4347
rect 633 4333 647 4347
rect 553 4273 567 4287
rect 593 4273 607 4287
rect 573 4253 587 4267
rect 653 4253 667 4267
rect 533 4193 547 4207
rect 813 4293 827 4307
rect 853 4193 867 4207
rect 713 4153 727 4167
rect 813 4153 827 4167
rect 833 4133 847 4147
rect 793 4113 807 4127
rect 252 4033 266 4047
rect 273 4033 287 4047
rect 433 4053 447 4067
rect 733 4053 747 4067
rect 393 4013 407 4027
rect 533 4014 547 4028
rect 673 4014 687 4028
rect 233 3993 247 4007
rect 293 3992 307 4006
rect 193 3953 207 3967
rect 353 3953 367 3967
rect 333 3833 347 3847
rect 253 3814 267 3828
rect 313 3814 327 3828
rect 433 3973 447 3987
rect 413 3913 427 3927
rect 393 3873 407 3887
rect 393 3833 407 3847
rect 53 3713 67 3727
rect 153 3772 167 3786
rect 193 3772 207 3786
rect 113 3633 127 3647
rect 173 3553 187 3567
rect 33 3534 47 3548
rect 93 3533 107 3547
rect 73 3473 87 3487
rect 293 3772 307 3786
rect 333 3772 347 3786
rect 253 3753 267 3767
rect 333 3751 347 3765
rect 193 3513 207 3527
rect 113 3294 127 3308
rect 173 3294 187 3308
rect 273 3294 287 3308
rect 133 3233 147 3247
rect 173 3193 187 3207
rect 353 3713 367 3727
rect 353 3553 367 3567
rect 353 3493 367 3507
rect 333 3233 347 3247
rect 413 3673 427 3687
rect 713 4012 727 4026
rect 473 3913 487 3927
rect 533 3913 547 3927
rect 673 3913 687 3927
rect 433 3633 447 3647
rect 473 3633 487 3647
rect 453 3613 467 3627
rect 453 3473 467 3487
rect 393 3433 407 3447
rect 433 3433 447 3447
rect 513 3633 527 3647
rect 493 3593 507 3607
rect 493 3553 507 3567
rect 473 3413 487 3427
rect 413 3373 427 3387
rect 373 3333 387 3347
rect 473 3333 487 3347
rect 393 3233 407 3247
rect 193 3113 207 3127
rect 253 3113 267 3127
rect 33 3014 47 3028
rect 93 3013 107 3027
rect 73 2953 87 2967
rect 53 2833 67 2847
rect 433 3113 447 3127
rect 393 3053 407 3067
rect 333 2953 347 2967
rect 373 2913 387 2927
rect 233 2833 247 2847
rect 93 2813 107 2827
rect 193 2813 207 2827
rect 113 2774 127 2788
rect 153 2774 167 2788
rect 113 2713 127 2727
rect 73 2693 87 2707
rect 213 2774 227 2788
rect 133 2693 147 2707
rect 193 2693 207 2707
rect 113 2653 127 2667
rect 173 2653 187 2667
rect 113 2513 127 2527
rect 133 2393 147 2407
rect 173 2393 187 2407
rect 273 2774 287 2788
rect 313 2774 327 2788
rect 493 3173 507 3187
rect 473 3033 487 3047
rect 433 2953 447 2967
rect 413 2833 427 2847
rect 413 2793 427 2807
rect 393 2753 407 2767
rect 253 2733 267 2747
rect 233 2653 247 2667
rect 213 2633 227 2647
rect 273 2713 287 2727
rect 253 2513 267 2527
rect 333 2732 347 2746
rect 613 3873 627 3887
rect 653 3814 667 3828
rect 713 3814 727 3828
rect 633 3753 647 3767
rect 593 3593 607 3607
rect 773 3973 787 3987
rect 813 4073 827 4087
rect 753 3933 767 3947
rect 793 3933 807 3947
rect 733 3752 747 3766
rect 713 3733 727 3747
rect 653 3613 667 3627
rect 793 3814 807 3828
rect 873 4173 887 4187
rect 853 4012 867 4026
rect 853 3913 867 3927
rect 773 3773 787 3787
rect 853 3773 867 3787
rect 853 3733 867 3747
rect 773 3693 787 3707
rect 853 3653 867 3667
rect 693 3593 707 3607
rect 753 3593 767 3607
rect 833 3593 847 3607
rect 673 3573 687 3587
rect 633 3514 647 3528
rect 533 3473 547 3487
rect 573 3472 587 3486
rect 673 3473 687 3487
rect 653 3373 667 3387
rect 553 3294 567 3308
rect 593 3294 607 3308
rect 573 3252 587 3266
rect 653 3252 667 3266
rect 753 3553 767 3567
rect 773 3514 787 3528
rect 753 3453 767 3467
rect 833 3433 847 3447
rect 753 3413 767 3427
rect 733 3294 747 3308
rect 773 3294 787 3308
rect 833 3294 847 3308
rect 613 3233 627 3247
rect 693 3233 707 3247
rect 773 3233 787 3247
rect 833 3253 847 3267
rect 813 3233 827 3247
rect 993 4314 1007 4328
rect 1053 4314 1067 4328
rect 1073 4213 1087 4227
rect 1173 4513 1187 4527
rect 1453 4893 1467 4907
rect 1473 4854 1487 4868
rect 1313 4832 1327 4846
rect 1453 4832 1467 4846
rect 1553 5033 1567 5047
rect 1633 5032 1647 5046
rect 1553 4973 1567 4987
rect 1513 4933 1527 4947
rect 1673 4973 1687 4987
rect 1513 4713 1527 4727
rect 1413 4693 1427 4707
rect 1293 4593 1307 4607
rect 1253 4573 1267 4587
rect 1473 4553 1487 4567
rect 1553 4554 1567 4568
rect 1213 4513 1227 4527
rect 1013 4133 1027 4147
rect 913 4113 927 4127
rect 953 4113 967 4127
rect 953 4073 967 4087
rect 1133 4473 1147 4487
rect 1193 4473 1207 4487
rect 1153 4433 1167 4447
rect 1313 4513 1327 4527
rect 1193 4373 1207 4387
rect 1273 4373 1287 4387
rect 1153 4334 1167 4348
rect 1233 4334 1247 4348
rect 1213 4292 1227 4306
rect 1353 4334 1367 4348
rect 1413 4334 1427 4348
rect 1213 4213 1227 4227
rect 1153 4153 1167 4167
rect 1113 4073 1127 4087
rect 1193 4073 1207 4087
rect 1073 4053 1087 4067
rect 1053 4034 1067 4048
rect 1093 4034 1107 4048
rect 933 3992 947 4006
rect 1033 3993 1047 4007
rect 1073 3933 1087 3947
rect 973 3873 987 3887
rect 1053 3873 1067 3887
rect 913 3833 927 3847
rect 993 3833 1007 3847
rect 1153 3933 1167 3947
rect 1293 4053 1307 4067
rect 1373 4273 1387 4287
rect 1573 4473 1587 4487
rect 1493 4373 1507 4387
rect 1593 4373 1607 4387
rect 1473 4333 1487 4347
rect 1533 4334 1547 4348
rect 1433 4314 1447 4328
rect 1413 4233 1427 4247
rect 1513 4292 1527 4306
rect 1493 4271 1507 4285
rect 1573 4293 1587 4307
rect 1573 4233 1587 4247
rect 1553 4213 1567 4227
rect 1433 4193 1447 4207
rect 1593 4113 1607 4127
rect 1353 4093 1367 4107
rect 1873 5453 1887 5467
rect 1953 5374 1967 5388
rect 1853 5332 1867 5346
rect 1913 5253 1927 5267
rect 1813 5113 1827 5127
rect 1853 5113 1867 5127
rect 1813 5074 1827 5088
rect 1753 5033 1767 5047
rect 1753 4893 1767 4907
rect 1713 4854 1727 4868
rect 1733 4812 1747 4826
rect 1793 4812 1807 4826
rect 1913 4973 1927 4987
rect 2053 5852 2067 5866
rect 2133 5873 2147 5887
rect 2113 5853 2127 5867
rect 2093 5713 2107 5727
rect 2133 5813 2147 5827
rect 2173 5813 2187 5827
rect 2153 5713 2167 5727
rect 2113 5673 2127 5687
rect 2053 5633 2067 5647
rect 2052 5593 2066 5607
rect 2073 5594 2087 5608
rect 2133 5594 2147 5608
rect 2093 5552 2107 5566
rect 2133 5553 2147 5567
rect 2053 5513 2067 5527
rect 2013 5374 2027 5388
rect 2113 5493 2127 5507
rect 1973 5193 1987 5207
rect 1953 4913 1967 4927
rect 1873 4873 1887 4887
rect 1913 4873 1927 4887
rect 1833 4853 1847 4867
rect 1693 4793 1707 4807
rect 1813 4793 1827 4807
rect 1653 4753 1667 4767
rect 1893 4793 1907 4807
rect 1893 4693 1907 4707
rect 1893 4633 1907 4647
rect 1793 4554 1807 4568
rect 1833 4554 1847 4568
rect 1933 4554 1947 4568
rect 2133 5453 2147 5467
rect 2233 5693 2247 5707
rect 2233 5653 2247 5667
rect 2313 6133 2327 6147
rect 2353 6114 2367 6128
rect 2293 6073 2307 6087
rect 2333 6072 2347 6086
rect 2453 6414 2467 6428
rect 2533 6413 2547 6427
rect 2613 6414 2627 6428
rect 2653 6414 2667 6428
rect 2993 6433 3007 6447
rect 2813 6414 2827 6428
rect 2873 6413 2887 6427
rect 2953 6414 2967 6428
rect 2993 6414 3007 6428
rect 3193 6414 3207 6428
rect 3233 6414 3247 6428
rect 2633 6372 2647 6386
rect 2473 6353 2487 6367
rect 2533 6353 2547 6367
rect 2433 6253 2447 6267
rect 2433 6193 2447 6207
rect 2413 6173 2427 6187
rect 2713 6372 2727 6386
rect 2833 6372 2847 6386
rect 2773 6333 2787 6347
rect 2533 6153 2547 6167
rect 2673 6153 2687 6167
rect 2713 6153 2727 6167
rect 2573 6113 2587 6127
rect 2433 6072 2447 6086
rect 2513 6072 2527 6086
rect 2573 6072 2587 6086
rect 2453 6033 2467 6047
rect 2833 6313 2847 6327
rect 2813 6253 2827 6267
rect 2793 6153 2807 6167
rect 2673 6072 2687 6086
rect 2733 6072 2747 6086
rect 2593 6013 2607 6027
rect 2633 5993 2647 6007
rect 2573 5933 2587 5947
rect 2413 5913 2427 5927
rect 2373 5894 2387 5908
rect 2453 5893 2467 5907
rect 2533 5894 2547 5908
rect 2393 5852 2407 5866
rect 2453 5852 2467 5866
rect 2353 5813 2367 5827
rect 2513 5813 2527 5827
rect 2373 5793 2387 5807
rect 2293 5773 2307 5787
rect 2373 5753 2387 5767
rect 2293 5713 2307 5727
rect 2273 5633 2287 5647
rect 2233 5594 2247 5608
rect 2273 5594 2287 5608
rect 2353 5573 2367 5587
rect 2193 5553 2207 5567
rect 2193 5532 2207 5546
rect 2173 5513 2187 5527
rect 2193 5473 2207 5487
rect 2293 5552 2307 5566
rect 2353 5473 2367 5487
rect 2493 5733 2507 5747
rect 2433 5594 2447 5608
rect 2413 5533 2427 5547
rect 2413 5493 2427 5507
rect 2493 5552 2507 5566
rect 2593 5852 2607 5866
rect 2633 5813 2647 5827
rect 2753 5933 2767 5947
rect 2673 5894 2687 5908
rect 2713 5894 2727 5908
rect 2813 5993 2827 6007
rect 2653 5793 2667 5807
rect 2633 5773 2647 5787
rect 2573 5733 2587 5747
rect 2553 5613 2567 5627
rect 2633 5713 2647 5727
rect 2773 5852 2787 5866
rect 2813 5852 2827 5866
rect 2973 6333 2987 6347
rect 2993 6313 3007 6327
rect 2873 6113 2887 6127
rect 2933 6114 2947 6128
rect 2913 6072 2927 6086
rect 2933 6033 2947 6047
rect 2993 6033 3007 6047
rect 2893 6013 2907 6027
rect 3233 6373 3247 6387
rect 3153 6333 3167 6347
rect 3133 6313 3147 6327
rect 3113 6193 3127 6207
rect 3073 6114 3087 6128
rect 3113 6114 3127 6128
rect 3013 6013 3027 6027
rect 2953 5893 2967 5907
rect 2833 5813 2847 5827
rect 2733 5793 2747 5807
rect 2913 5852 2927 5866
rect 2973 5852 2987 5866
rect 3093 6072 3107 6086
rect 3073 6013 3087 6027
rect 3113 5973 3127 5987
rect 3053 5852 3067 5866
rect 3013 5773 3027 5787
rect 2873 5733 2887 5747
rect 2913 5733 2927 5747
rect 2673 5693 2687 5707
rect 2673 5653 2687 5667
rect 2653 5633 2667 5647
rect 2593 5552 2607 5566
rect 2633 5552 2647 5566
rect 2513 5533 2527 5547
rect 2633 5493 2647 5507
rect 2453 5473 2467 5487
rect 2373 5453 2387 5467
rect 2413 5453 2427 5467
rect 2313 5413 2327 5427
rect 2153 5333 2167 5347
rect 2073 5293 2087 5307
rect 2033 5233 2047 5247
rect 2233 5173 2247 5187
rect 2213 5113 2227 5127
rect 2033 4854 2047 4868
rect 2013 4773 2027 4787
rect 2093 4693 2107 4707
rect 2133 4853 2147 4867
rect 2053 4653 2067 4667
rect 2113 4653 2127 4667
rect 1693 4512 1707 4526
rect 1812 4512 1826 4526
rect 1833 4512 1847 4526
rect 1913 4512 1927 4526
rect 1733 4473 1747 4487
rect 1773 4473 1787 4487
rect 1813 4473 1827 4487
rect 1953 4473 1967 4487
rect 1633 4353 1647 4367
rect 1613 4073 1627 4087
rect 1673 4334 1687 4348
rect 1713 4334 1727 4348
rect 1953 4373 1967 4387
rect 1793 4333 1807 4347
rect 1853 4334 1867 4348
rect 1733 4292 1747 4306
rect 1773 4292 1787 4306
rect 1693 4273 1707 4287
rect 1693 4193 1707 4207
rect 1673 4113 1687 4127
rect 1433 4053 1447 4067
rect 1633 4053 1647 4067
rect 1473 4034 1487 4048
rect 1513 4034 1527 4048
rect 1353 3993 1367 4007
rect 1413 3992 1427 4006
rect 1273 3973 1287 3987
rect 1333 3973 1347 3987
rect 1213 3953 1227 3967
rect 1073 3814 1087 3828
rect 1073 3793 1087 3807
rect 973 3772 987 3786
rect 1033 3752 1047 3766
rect 913 3713 927 3727
rect 893 3593 907 3607
rect 1113 3893 1127 3907
rect 1193 3893 1207 3907
rect 1473 3953 1487 3967
rect 1373 3913 1387 3927
rect 1172 3793 1186 3807
rect 1193 3792 1207 3806
rect 1333 3793 1347 3807
rect 1393 3813 1407 3827
rect 1353 3673 1367 3687
rect 1293 3633 1307 3647
rect 1493 3873 1507 3887
rect 1473 3733 1487 3747
rect 1453 3713 1467 3727
rect 1293 3592 1307 3606
rect 1393 3593 1407 3607
rect 1093 3573 1107 3587
rect 1153 3573 1167 3587
rect 873 3553 887 3567
rect 913 3553 927 3567
rect 953 3514 967 3528
rect 993 3514 1007 3528
rect 1093 3514 1107 3528
rect 893 3472 907 3486
rect 933 3413 947 3427
rect 1013 3453 1027 3467
rect 993 3393 1007 3407
rect 933 3294 947 3308
rect 993 3293 1007 3307
rect 913 3252 927 3266
rect 953 3252 967 3266
rect 793 3193 807 3207
rect 773 3053 787 3067
rect 593 2994 607 3008
rect 673 2993 687 3007
rect 733 2994 747 3008
rect 513 2953 527 2967
rect 573 2952 587 2966
rect 473 2913 487 2927
rect 713 2952 727 2966
rect 713 2913 727 2927
rect 673 2793 687 2807
rect 533 2752 547 2766
rect 393 2713 407 2727
rect 433 2713 447 2727
rect 373 2693 387 2707
rect 353 2653 367 2667
rect 293 2613 307 2627
rect 313 2513 327 2527
rect 293 2432 307 2446
rect 353 2432 367 2446
rect 53 2333 67 2347
rect 193 2333 207 2347
rect 253 2333 267 2347
rect 373 2273 387 2287
rect 53 2233 67 2247
rect 33 2192 47 2206
rect 193 2213 207 2227
rect 113 1954 127 1968
rect 153 1954 167 1968
rect 253 1954 267 1968
rect 293 1954 307 1968
rect 333 1954 347 1968
rect 693 2752 707 2766
rect 793 2952 807 2966
rect 753 2893 767 2907
rect 773 2773 787 2787
rect 453 2593 467 2607
rect 693 2573 707 2587
rect 673 2513 687 2527
rect 533 2473 547 2487
rect 433 2393 447 2407
rect 493 2433 507 2447
rect 473 2333 487 2347
rect 473 2113 487 2127
rect 413 2093 427 2107
rect 93 1913 107 1927
rect 173 1912 187 1926
rect 253 1913 267 1927
rect 153 1893 167 1907
rect 93 1773 107 1787
rect 293 1893 307 1907
rect 253 1853 267 1867
rect 113 1734 127 1748
rect 213 1692 227 1706
rect 273 1692 287 1706
rect 353 1912 367 1926
rect 393 1913 407 1927
rect 313 1793 327 1807
rect 393 1793 407 1807
rect 353 1734 367 1748
rect 293 1633 307 1647
rect 273 1593 287 1607
rect 193 1553 207 1567
rect 153 1513 167 1527
rect 113 1434 127 1448
rect 73 1393 87 1407
rect 133 1392 147 1406
rect 133 1273 147 1287
rect 173 1213 187 1227
rect 113 1153 127 1167
rect 233 1473 247 1487
rect 213 1434 227 1448
rect 213 1273 227 1287
rect 193 1153 207 1167
rect 193 953 207 967
rect 133 914 147 928
rect 353 1633 367 1647
rect 333 1473 347 1487
rect 593 2432 607 2446
rect 533 2393 547 2407
rect 433 2033 447 2047
rect 493 2033 507 2047
rect 413 1734 427 1748
rect 513 1993 527 2007
rect 473 1954 487 1968
rect 493 1912 507 1926
rect 493 1773 507 1787
rect 433 1692 447 1706
rect 473 1692 487 1706
rect 433 1553 447 1567
rect 513 1533 527 1547
rect 433 1513 447 1527
rect 473 1493 487 1507
rect 513 1493 527 1507
rect 393 1393 407 1407
rect 253 1253 267 1267
rect 293 1253 307 1267
rect 233 1213 247 1227
rect 453 1293 467 1307
rect 493 1293 507 1307
rect 393 1273 407 1287
rect 353 1213 367 1227
rect 453 1214 467 1228
rect 313 1172 327 1186
rect 353 1172 367 1186
rect 393 1172 407 1186
rect 433 1172 447 1186
rect 473 1172 487 1186
rect 273 1133 287 1147
rect 593 2212 607 2226
rect 693 2433 707 2447
rect 813 2833 827 2847
rect 793 2533 807 2547
rect 953 3233 967 3247
rect 993 3113 1007 3127
rect 973 2994 987 3008
rect 893 2952 907 2966
rect 893 2933 907 2947
rect 873 2833 887 2847
rect 853 2774 867 2788
rect 853 2633 867 2647
rect 833 2513 847 2527
rect 753 2474 767 2488
rect 813 2432 827 2446
rect 733 2273 747 2287
rect 673 2212 687 2226
rect 633 2173 647 2187
rect 713 2153 727 2167
rect 573 2113 587 2127
rect 673 1993 687 2007
rect 593 1954 607 1968
rect 633 1954 647 1968
rect 773 2413 787 2427
rect 773 2353 787 2367
rect 753 2093 767 2107
rect 753 1954 767 1968
rect 693 1912 707 1926
rect 693 1873 707 1887
rect 593 1853 607 1867
rect 653 1853 667 1867
rect 653 1734 667 1748
rect 733 1734 747 1748
rect 713 1693 727 1707
rect 673 1613 687 1627
rect 633 1513 647 1527
rect 613 1473 627 1487
rect 573 1433 587 1447
rect 693 1434 707 1448
rect 593 1392 607 1406
rect 553 1293 567 1307
rect 533 1233 547 1247
rect 513 1033 527 1047
rect 513 953 527 967
rect 213 914 227 928
rect 93 753 107 767
rect 193 872 207 886
rect 153 793 167 807
rect 113 713 127 727
rect 153 713 167 727
rect 153 694 167 708
rect 133 652 147 666
rect 273 914 287 928
rect 353 914 367 928
rect 433 914 447 928
rect 473 914 487 928
rect 693 1313 707 1327
rect 593 1273 607 1287
rect 633 1273 647 1287
rect 633 1214 647 1228
rect 673 1214 687 1228
rect 553 1173 567 1187
rect 673 1172 687 1186
rect 613 1133 627 1147
rect 613 1112 627 1126
rect 533 933 547 947
rect 573 933 587 947
rect 273 873 287 887
rect 333 872 347 886
rect 433 873 447 887
rect 233 753 247 767
rect 213 694 227 708
rect 193 613 207 627
rect 113 533 127 547
rect 293 694 307 708
rect 453 793 467 807
rect 533 793 547 807
rect 553 693 567 707
rect 313 652 327 666
rect 473 652 487 666
rect 233 533 247 547
rect 153 473 167 487
rect 213 473 227 487
rect 273 493 287 507
rect 453 493 467 507
rect 553 413 567 427
rect 133 352 147 366
rect 253 353 267 367
rect 293 333 307 347
rect 153 213 167 227
rect 313 213 327 227
rect 493 394 507 408
rect 513 352 527 366
rect 553 353 567 367
rect 1073 3433 1087 3447
rect 1173 3513 1187 3527
rect 1253 3514 1267 3528
rect 1233 3393 1247 3407
rect 1393 3572 1407 3586
rect 1333 3514 1347 3528
rect 1433 3514 1447 3528
rect 1473 3693 1487 3707
rect 1373 3472 1387 3486
rect 1333 3453 1347 3467
rect 1313 3353 1327 3367
rect 1353 3353 1367 3367
rect 1193 3333 1207 3347
rect 1173 3313 1187 3327
rect 1233 3293 1247 3307
rect 1073 3252 1087 3266
rect 1053 3193 1067 3207
rect 1173 3193 1187 3207
rect 1153 3053 1167 3067
rect 1053 2994 1067 3008
rect 1093 2994 1107 3008
rect 1013 2913 1027 2927
rect 993 2893 1007 2907
rect 933 2813 947 2827
rect 973 2813 987 2827
rect 913 2774 927 2788
rect 993 2774 1007 2788
rect 933 2732 947 2746
rect 973 2733 987 2747
rect 993 2573 1007 2587
rect 953 2553 967 2567
rect 873 2413 887 2427
rect 973 2432 987 2446
rect 1073 2952 1087 2966
rect 1133 2953 1147 2967
rect 1113 2933 1127 2947
rect 1093 2833 1107 2847
rect 1053 2774 1067 2788
rect 1073 2732 1087 2746
rect 1133 2613 1147 2627
rect 1313 3293 1327 3307
rect 1413 3413 1427 3427
rect 1513 3713 1527 3727
rect 1553 4033 1567 4047
rect 1553 3992 1567 4006
rect 1593 3992 1607 4006
rect 1633 3992 1647 4006
rect 1553 3933 1567 3947
rect 1633 3873 1647 3887
rect 1573 3814 1587 3828
rect 1553 3773 1567 3787
rect 1533 3513 1547 3527
rect 1673 3772 1687 3786
rect 1633 3673 1647 3687
rect 1593 3533 1607 3547
rect 1673 3513 1687 3527
rect 1493 3473 1507 3487
rect 1473 3393 1487 3407
rect 1553 3393 1567 3407
rect 1533 3353 1547 3367
rect 1373 3293 1387 3307
rect 1473 3294 1487 3308
rect 1273 3273 1287 3287
rect 1513 3253 1527 3267
rect 1393 3173 1407 3187
rect 1273 3153 1287 3167
rect 1333 3153 1347 3167
rect 1253 3013 1267 3027
rect 1173 2994 1187 3008
rect 1233 2994 1247 3008
rect 1333 3113 1347 3127
rect 1313 3013 1327 3027
rect 1253 2952 1267 2966
rect 1233 2873 1247 2887
rect 1173 2813 1187 2827
rect 1053 2474 1067 2488
rect 1093 2474 1107 2488
rect 953 2413 967 2427
rect 1013 2413 1027 2427
rect 933 2393 947 2407
rect 853 2333 867 2347
rect 913 2313 927 2327
rect 873 2212 887 2226
rect 933 2254 947 2268
rect 933 2213 947 2227
rect 913 2153 927 2167
rect 793 2053 807 2067
rect 833 1954 847 1968
rect 873 1954 887 1968
rect 793 1912 807 1926
rect 773 1873 787 1887
rect 893 1893 907 1907
rect 853 1813 867 1827
rect 773 1753 787 1767
rect 753 1693 767 1707
rect 733 1593 747 1607
rect 793 1734 807 1748
rect 853 1734 867 1748
rect 793 1553 807 1567
rect 773 1533 787 1547
rect 853 1633 867 1647
rect 813 1513 827 1527
rect 833 1473 847 1487
rect 753 1434 767 1448
rect 773 1392 787 1406
rect 833 1393 847 1407
rect 773 1353 787 1367
rect 813 1353 827 1367
rect 733 1153 747 1167
rect 713 1113 727 1127
rect 673 973 687 987
rect 653 914 667 928
rect 673 872 687 886
rect 913 1853 927 1867
rect 893 1633 907 1647
rect 873 1613 887 1627
rect 893 1573 907 1587
rect 873 1513 887 1527
rect 993 2254 1007 2268
rect 1153 2432 1167 2446
rect 1253 2732 1267 2746
rect 1273 2693 1287 2707
rect 1233 2653 1247 2667
rect 1213 2593 1227 2607
rect 1113 2393 1127 2407
rect 1153 2393 1167 2407
rect 1193 2393 1207 2407
rect 1253 2553 1267 2567
rect 1233 2473 1247 2487
rect 1233 2432 1247 2446
rect 1413 3153 1427 3167
rect 1493 3113 1507 3127
rect 1413 3053 1427 3067
rect 1453 2994 1467 3008
rect 1493 2994 1507 3008
rect 1473 2933 1487 2947
rect 1453 2893 1467 2907
rect 1393 2853 1407 2867
rect 1433 2833 1447 2847
rect 1453 2773 1467 2787
rect 1413 2732 1427 2746
rect 1453 2733 1467 2747
rect 1373 2593 1387 2607
rect 1413 2533 1427 2547
rect 1373 2513 1387 2527
rect 1213 2293 1227 2307
rect 1093 2253 1107 2267
rect 1153 2254 1167 2268
rect 1013 2212 1027 2226
rect 1073 2213 1087 2227
rect 1033 2013 1047 2027
rect 1113 2213 1127 2227
rect 1053 1893 1067 1907
rect 1013 1833 1027 1847
rect 993 1753 1007 1767
rect 1033 1734 1047 1748
rect 1093 1734 1107 1748
rect 953 1693 967 1707
rect 1013 1692 1027 1706
rect 1073 1553 1087 1567
rect 993 1533 1007 1547
rect 973 1453 987 1467
rect 893 1433 907 1447
rect 933 1434 947 1448
rect 1053 1473 1067 1487
rect 1013 1434 1027 1448
rect 913 1392 927 1406
rect 873 1353 887 1367
rect 953 1353 967 1367
rect 933 1313 947 1327
rect 853 1153 867 1167
rect 793 1033 807 1047
rect 793 973 807 987
rect 752 873 766 887
rect 773 873 787 887
rect 613 833 627 847
rect 673 833 687 847
rect 633 733 647 747
rect 733 733 747 747
rect 613 652 627 666
rect 633 413 647 427
rect 593 393 607 407
rect 473 333 487 347
rect 573 333 587 347
rect 433 213 447 227
rect 553 193 567 207
rect 693 352 707 366
rect 653 313 667 327
rect 933 1133 947 1147
rect 873 914 887 928
rect 833 872 847 886
rect 893 873 907 887
rect 793 833 807 847
rect 853 853 867 867
rect 933 853 947 867
rect 833 733 847 747
rect 893 694 907 708
rect 933 694 947 708
rect 793 652 807 666
rect 773 453 787 467
rect 913 453 927 467
rect 752 353 766 367
rect 833 394 847 408
rect 773 352 787 366
rect 813 352 827 366
rect 853 333 867 347
rect 753 313 767 327
rect 633 293 647 307
rect 733 293 747 307
rect 733 193 747 207
rect 693 173 707 187
rect 113 132 127 146
rect 353 132 367 146
rect 553 133 567 147
rect 613 132 627 146
rect 653 132 667 146
rect 693 132 707 146
rect 733 132 747 146
rect 793 174 807 188
rect 1173 2212 1187 2226
rect 1333 2293 1347 2307
rect 1253 2254 1267 2268
rect 1293 2254 1307 2268
rect 1493 2772 1507 2786
rect 1493 2473 1507 2487
rect 1493 2373 1507 2387
rect 1473 2313 1487 2327
rect 1533 3073 1547 3087
rect 1613 3313 1627 3327
rect 1573 3294 1587 3308
rect 1633 3294 1647 3308
rect 1753 4113 1767 4127
rect 1913 4292 1927 4306
rect 1953 4292 1967 4306
rect 1873 4273 1887 4287
rect 1893 4073 1907 4087
rect 1793 4033 1807 4047
rect 1873 4034 1887 4048
rect 1713 3992 1727 4006
rect 1773 3992 1787 4006
rect 1813 3893 1827 3907
rect 1813 3833 1827 3847
rect 1853 3833 1867 3847
rect 1753 3772 1767 3786
rect 1793 3772 1807 3786
rect 1873 3814 1887 3828
rect 1853 3673 1867 3687
rect 1733 3633 1747 3647
rect 1713 3613 1727 3627
rect 1753 3573 1767 3587
rect 1713 3533 1727 3547
rect 1733 3433 1747 3447
rect 1813 3473 1827 3487
rect 1813 3393 1827 3407
rect 1773 3353 1787 3367
rect 1693 3312 1707 3326
rect 1773 3294 1787 3308
rect 2093 4554 2107 4568
rect 2193 4812 2207 4826
rect 2253 5093 2267 5107
rect 2373 5374 2387 5388
rect 2453 5413 2467 5427
rect 2493 5393 2507 5407
rect 2553 5393 2567 5407
rect 2393 5332 2407 5346
rect 2453 5332 2467 5346
rect 2353 5253 2367 5267
rect 2313 5074 2327 5088
rect 2293 4953 2307 4967
rect 2373 5093 2387 5107
rect 2353 5074 2367 5088
rect 2373 5032 2387 5046
rect 2353 4973 2367 4987
rect 2353 4933 2367 4947
rect 2273 4893 2287 4907
rect 2333 4893 2347 4907
rect 2253 4854 2267 4868
rect 2173 4653 2187 4667
rect 2153 4613 2167 4627
rect 2153 4553 2167 4567
rect 2113 4512 2127 4526
rect 2073 4393 2087 4407
rect 2133 4393 2147 4407
rect 2033 4334 2047 4348
rect 2093 4292 2107 4306
rect 2053 4273 2067 4287
rect 2073 4233 2087 4247
rect 1993 4073 2007 4087
rect 1933 4034 1947 4048
rect 1973 4034 1987 4048
rect 2033 4033 2047 4047
rect 1953 3973 1967 3987
rect 1953 3814 1967 3828
rect 1933 3772 1947 3786
rect 1933 3713 1947 3727
rect 1853 3533 1867 3547
rect 1893 3533 1907 3547
rect 1973 3653 1987 3667
rect 2193 4553 2207 4567
rect 2253 4733 2267 4747
rect 2313 4854 2327 4868
rect 2433 5313 2447 5327
rect 2433 5253 2447 5267
rect 2413 5233 2427 5247
rect 2593 5393 2607 5407
rect 2613 5373 2627 5387
rect 2533 5332 2547 5346
rect 2573 5332 2587 5346
rect 2493 5173 2507 5187
rect 2533 5153 2547 5167
rect 2433 5032 2447 5046
rect 2473 5032 2487 5046
rect 2433 5013 2447 5027
rect 2453 4953 2467 4967
rect 2413 4873 2427 4887
rect 2393 4853 2407 4867
rect 2333 4812 2347 4826
rect 2373 4812 2387 4826
rect 2373 4773 2387 4787
rect 2333 4693 2347 4707
rect 2313 4613 2327 4627
rect 2273 4573 2287 4587
rect 2253 4554 2267 4568
rect 2353 4573 2367 4587
rect 2233 4512 2247 4526
rect 2273 4512 2287 4526
rect 2333 4512 2347 4526
rect 2233 4413 2247 4427
rect 2193 4373 2207 4387
rect 2233 4334 2247 4348
rect 2273 4334 2287 4348
rect 2173 4292 2187 4306
rect 2213 4292 2227 4306
rect 2293 4293 2307 4307
rect 2253 4273 2267 4287
rect 2173 4213 2187 4227
rect 2293 4233 2307 4247
rect 2213 4173 2227 4187
rect 2173 4153 2187 4167
rect 2073 3992 2087 4006
rect 2153 3992 2167 4006
rect 2113 3973 2127 3987
rect 2313 4093 2327 4107
rect 2373 4553 2387 4567
rect 2433 4853 2447 4867
rect 2433 4812 2447 4826
rect 2953 5673 2967 5687
rect 3053 5653 3067 5667
rect 2953 5633 2967 5647
rect 2733 5594 2747 5608
rect 2673 5493 2687 5507
rect 2813 5594 2827 5608
rect 2853 5594 2867 5608
rect 2793 5493 2807 5507
rect 2673 5433 2687 5447
rect 2713 5433 2727 5447
rect 2653 5392 2667 5406
rect 2653 5332 2667 5346
rect 2733 5413 2747 5427
rect 2773 5374 2787 5388
rect 2873 5533 2887 5547
rect 2833 5513 2847 5527
rect 2713 5332 2727 5346
rect 2813 5333 2827 5347
rect 2753 5313 2767 5327
rect 2693 5293 2707 5307
rect 2673 5273 2687 5287
rect 2673 5233 2687 5247
rect 2553 5133 2567 5147
rect 2633 5133 2647 5147
rect 2533 4873 2547 4887
rect 2513 4854 2527 4868
rect 2593 5113 2607 5127
rect 2653 5074 2667 5088
rect 2573 5032 2587 5046
rect 2613 5013 2627 5027
rect 2593 4993 2607 5007
rect 2573 4973 2587 4987
rect 2533 4793 2547 4807
rect 2493 4753 2507 4767
rect 2453 4693 2467 4707
rect 2513 4613 2527 4627
rect 2453 4554 2467 4568
rect 2433 4512 2447 4526
rect 2473 4512 2487 4526
rect 2433 4433 2447 4447
rect 2393 4334 2407 4348
rect 2673 4953 2687 4967
rect 2593 4933 2607 4947
rect 2593 4853 2607 4867
rect 2713 5273 2727 5287
rect 2753 5273 2767 5287
rect 2593 4733 2607 4747
rect 2613 4693 2627 4707
rect 2673 4793 2687 4807
rect 2673 4733 2687 4747
rect 2653 4573 2667 4587
rect 2693 4573 2707 4587
rect 2673 4553 2687 4567
rect 2553 4512 2567 4526
rect 2593 4512 2607 4526
rect 2533 4433 2547 4447
rect 2533 4393 2547 4407
rect 2512 4333 2526 4347
rect 2533 4333 2547 4347
rect 2573 4334 2587 4348
rect 2493 4173 2507 4187
rect 2553 4292 2567 4306
rect 2593 4292 2607 4306
rect 2673 4353 2687 4367
rect 2653 4333 2667 4347
rect 2633 4153 2647 4167
rect 2513 4133 2527 4147
rect 2533 4093 2547 4107
rect 2633 4093 2647 4107
rect 2513 4053 2527 4067
rect 2413 4034 2427 4048
rect 2453 4034 2467 4048
rect 2553 4073 2567 4087
rect 2333 3992 2347 4006
rect 2393 3992 2407 4006
rect 2493 3992 2507 4006
rect 2533 3992 2547 4006
rect 2293 3933 2307 3947
rect 2413 3893 2427 3907
rect 2213 3873 2227 3887
rect 2273 3814 2287 3828
rect 2352 3813 2366 3827
rect 2373 3814 2387 3828
rect 2453 3853 2467 3867
rect 2493 3814 2507 3828
rect 2173 3793 2187 3807
rect 2053 3773 2067 3787
rect 2033 3732 2047 3746
rect 1993 3533 2007 3547
rect 2213 3772 2227 3786
rect 2213 3733 2227 3747
rect 2173 3653 2187 3667
rect 2133 3573 2147 3587
rect 2113 3514 2127 3528
rect 1873 3473 1887 3487
rect 1853 3313 1867 3327
rect 1613 3252 1627 3266
rect 1693 3252 1707 3266
rect 1653 3193 1667 3207
rect 1613 2994 1627 3008
rect 1653 2994 1667 3008
rect 1573 2813 1587 2827
rect 1673 2953 1687 2967
rect 1653 2853 1667 2867
rect 1613 2833 1627 2847
rect 1553 2793 1567 2807
rect 1533 2773 1547 2787
rect 1553 2732 1567 2746
rect 1593 2732 1607 2746
rect 1553 2653 1567 2667
rect 1753 3253 1767 3267
rect 1733 3213 1747 3227
rect 1713 3133 1727 3147
rect 1713 2994 1727 3008
rect 1793 3252 1807 3266
rect 1793 3193 1807 3207
rect 1953 3413 1967 3427
rect 1973 3313 1987 3327
rect 2033 3313 2047 3327
rect 1873 3193 1887 3207
rect 1853 3173 1867 3187
rect 1933 3294 1947 3308
rect 1953 3213 1967 3227
rect 1953 3192 1967 3206
rect 1793 3013 1807 3027
rect 1893 3013 1907 3027
rect 1753 2993 1767 3007
rect 1893 2992 1907 3006
rect 1993 3173 2007 3187
rect 2053 3293 2067 3307
rect 1773 2952 1787 2966
rect 1713 2933 1727 2947
rect 1773 2873 1787 2887
rect 1713 2853 1727 2867
rect 1813 2853 1827 2867
rect 1693 2833 1707 2847
rect 1693 2812 1707 2826
rect 1733 2813 1747 2827
rect 1673 2733 1687 2747
rect 1773 2774 1787 2788
rect 1753 2732 1767 2746
rect 1693 2693 1707 2707
rect 1673 2633 1687 2647
rect 1553 2593 1567 2607
rect 1653 2593 1667 2607
rect 1553 2553 1567 2567
rect 1673 2533 1687 2547
rect 1573 2493 1587 2507
rect 1533 2473 1547 2487
rect 1613 2474 1627 2488
rect 1673 2474 1687 2488
rect 1653 2453 1667 2467
rect 1533 2433 1547 2447
rect 1553 2413 1567 2427
rect 1553 2373 1567 2387
rect 1533 2293 1547 2307
rect 1513 2273 1527 2287
rect 1553 2253 1567 2267
rect 1633 2433 1647 2447
rect 1673 2413 1687 2427
rect 1653 2353 1667 2367
rect 1213 2093 1227 2107
rect 1193 1954 1207 1968
rect 1233 1954 1247 1968
rect 1173 1912 1187 1926
rect 1173 1873 1187 1887
rect 1213 1853 1227 1867
rect 1433 2213 1447 2227
rect 1313 2133 1327 2147
rect 1313 2093 1327 2107
rect 1273 1753 1287 1767
rect 1213 1734 1227 1748
rect 1253 1734 1267 1748
rect 1373 1954 1387 1968
rect 1413 1953 1427 1967
rect 1333 1873 1347 1887
rect 1413 1853 1427 1867
rect 1393 1793 1407 1807
rect 1193 1692 1207 1706
rect 1173 1673 1187 1687
rect 1113 1513 1127 1527
rect 1113 1453 1127 1467
rect 1073 1433 1087 1447
rect 1293 1733 1307 1747
rect 1353 1734 1367 1748
rect 1413 1733 1427 1747
rect 1293 1692 1307 1706
rect 1333 1673 1347 1687
rect 1253 1633 1267 1647
rect 1313 1573 1327 1587
rect 1253 1553 1267 1567
rect 1193 1434 1207 1448
rect 1313 1513 1327 1527
rect 1333 1453 1347 1467
rect 1293 1434 1307 1448
rect 1053 1392 1067 1406
rect 1093 1392 1107 1406
rect 1173 1393 1187 1407
rect 1133 1313 1147 1327
rect 1153 1273 1167 1287
rect 1093 1233 1107 1247
rect 993 1133 1007 1147
rect 1133 1172 1147 1186
rect 1173 1233 1187 1247
rect 1073 1093 1087 1107
rect 1133 1093 1147 1107
rect 1033 833 1047 847
rect 1113 833 1127 847
rect 973 793 987 807
rect 1273 1392 1287 1406
rect 1213 1213 1227 1227
rect 1273 1214 1287 1228
rect 1213 1153 1227 1167
rect 1253 1132 1267 1146
rect 1193 1073 1207 1087
rect 1293 1093 1307 1107
rect 1313 1073 1327 1087
rect 1053 773 1067 787
rect 1133 773 1147 787
rect 973 733 987 747
rect 973 693 987 707
rect 973 652 987 666
rect 973 613 987 627
rect 953 453 967 467
rect 933 433 947 447
rect 1113 652 1127 666
rect 993 493 1007 507
rect 993 453 1007 467
rect 1233 872 1247 886
rect 1273 872 1287 886
rect 1313 773 1327 787
rect 1253 694 1267 708
rect 1313 694 1327 708
rect 1233 652 1247 666
rect 1273 633 1287 647
rect 1313 633 1327 647
rect 1213 453 1227 467
rect 1133 413 1147 427
rect 1173 413 1187 427
rect 973 394 987 408
rect 933 353 947 367
rect 1413 1533 1427 1547
rect 1473 2173 1487 2187
rect 1513 2193 1527 2207
rect 1493 2133 1507 2147
rect 1473 2093 1487 2107
rect 1513 2053 1527 2067
rect 1473 1993 1487 2007
rect 1553 1993 1567 2007
rect 1453 1793 1467 1807
rect 1613 2254 1627 2268
rect 1833 2774 1847 2788
rect 1833 2733 1847 2747
rect 1833 2693 1847 2707
rect 1773 2673 1787 2687
rect 1813 2673 1827 2687
rect 1773 2513 1787 2527
rect 1813 2513 1827 2527
rect 1733 2474 1747 2488
rect 1813 2453 1827 2467
rect 1773 2413 1787 2427
rect 1833 2413 1847 2427
rect 1753 2313 1767 2327
rect 1733 2293 1747 2307
rect 1593 2213 1607 2227
rect 1633 2212 1647 2226
rect 1673 2212 1687 2226
rect 1653 2173 1667 2187
rect 1593 2113 1607 2127
rect 1633 2053 1647 2067
rect 1573 1973 1587 1987
rect 1613 1973 1627 1987
rect 1553 1954 1567 1968
rect 1493 1913 1507 1927
rect 1493 1873 1507 1887
rect 1573 1893 1587 1907
rect 1533 1833 1547 1847
rect 1513 1793 1527 1807
rect 1553 1733 1567 1747
rect 1533 1692 1547 1706
rect 1593 1753 1607 1767
rect 1493 1633 1507 1647
rect 1453 1473 1467 1487
rect 1513 1473 1527 1487
rect 1433 1453 1447 1467
rect 1373 1353 1387 1367
rect 1413 1313 1427 1327
rect 1493 1333 1507 1347
rect 1433 1233 1447 1247
rect 1453 1214 1467 1228
rect 1433 1172 1447 1186
rect 1493 1173 1507 1187
rect 1473 1153 1487 1167
rect 1413 1093 1427 1107
rect 1493 1093 1507 1107
rect 1353 872 1367 886
rect 1333 533 1347 547
rect 1333 493 1347 507
rect 1453 833 1467 847
rect 1433 773 1447 787
rect 1413 694 1427 708
rect 1493 693 1507 707
rect 1353 453 1367 467
rect 1333 413 1347 427
rect 1433 652 1447 666
rect 1493 652 1507 666
rect 1493 533 1507 547
rect 1353 373 1367 387
rect 993 352 1007 366
rect 1213 352 1227 366
rect 1253 352 1267 366
rect 1293 352 1307 366
rect 1333 352 1347 366
rect 1033 333 1047 347
rect 1113 333 1127 347
rect 973 174 987 188
rect 833 132 847 146
rect 913 132 927 146
rect 953 132 967 146
rect 1353 213 1367 227
rect 1193 173 1207 187
rect 1273 174 1287 188
rect 1393 394 1407 408
rect 1433 394 1447 408
rect 1453 352 1467 366
rect 1413 293 1427 307
rect 1553 1573 1567 1587
rect 1693 2013 1707 2027
rect 1733 2173 1747 2187
rect 1833 2273 1847 2287
rect 1793 2254 1807 2268
rect 1933 2833 1947 2847
rect 1953 2774 1967 2788
rect 1913 2732 1927 2746
rect 1913 2653 1927 2667
rect 1953 2633 1967 2647
rect 1913 2533 1927 2547
rect 1993 2952 2007 2966
rect 1993 2913 2007 2927
rect 1993 2732 2007 2746
rect 1993 2693 2007 2707
rect 2093 3472 2107 3486
rect 2293 3772 2307 3786
rect 2353 3772 2367 3786
rect 2253 3713 2267 3727
rect 2293 3713 2307 3727
rect 2253 3533 2267 3547
rect 2353 3693 2367 3707
rect 2213 3493 2227 3507
rect 2193 3453 2207 3467
rect 2273 3453 2287 3467
rect 2173 3433 2187 3447
rect 2133 3393 2147 3407
rect 2173 3233 2187 3247
rect 2073 3213 2087 3227
rect 2113 3213 2127 3227
rect 2153 3213 2167 3227
rect 2153 2993 2167 3007
rect 2173 2973 2187 2987
rect 2053 2952 2067 2966
rect 2093 2952 2107 2966
rect 2153 2953 2167 2967
rect 2133 2893 2147 2907
rect 2093 2873 2107 2887
rect 2133 2774 2147 2788
rect 2033 2732 2047 2746
rect 2013 2653 2027 2667
rect 2033 2633 2047 2647
rect 2213 3393 2227 3407
rect 2313 3393 2327 3407
rect 2233 3333 2247 3347
rect 2273 3333 2287 3347
rect 2313 3294 2327 3308
rect 2293 3233 2307 3247
rect 2253 3173 2267 3187
rect 2333 3013 2347 3027
rect 2273 2994 2287 3008
rect 2333 2973 2347 2987
rect 2213 2953 2227 2967
rect 2293 2953 2307 2967
rect 2473 3772 2487 3786
rect 2433 3733 2447 3747
rect 2413 3713 2427 3727
rect 2373 3673 2387 3687
rect 2393 3333 2407 3347
rect 2373 3293 2387 3307
rect 2373 3252 2387 3266
rect 2393 3133 2407 3147
rect 2513 3633 2527 3647
rect 2433 3533 2447 3547
rect 2493 3514 2507 3528
rect 2473 3433 2487 3447
rect 2453 3294 2467 3308
rect 2433 3252 2447 3266
rect 2473 3233 2487 3247
rect 2413 3073 2427 3087
rect 2393 3013 2407 3027
rect 2433 2994 2447 3008
rect 2493 3073 2507 3087
rect 2253 2913 2267 2927
rect 2193 2873 2207 2887
rect 2233 2833 2247 2847
rect 2173 2813 2187 2827
rect 2213 2773 2227 2787
rect 2353 2732 2367 2746
rect 2213 2713 2227 2727
rect 2233 2693 2247 2707
rect 2213 2633 2227 2647
rect 2033 2533 2047 2547
rect 2073 2533 2087 2547
rect 2153 2533 2167 2547
rect 1973 2473 1987 2487
rect 1873 2433 1887 2447
rect 1873 2293 1887 2307
rect 1853 2253 1867 2267
rect 1753 2153 1767 2167
rect 1853 2053 1867 2067
rect 1713 1993 1727 2007
rect 1813 1972 1827 1986
rect 1773 1954 1787 1968
rect 1673 1913 1687 1927
rect 1653 1873 1667 1887
rect 1713 1912 1727 1926
rect 1713 1873 1727 1887
rect 1933 2413 1947 2427
rect 1913 2333 1927 2347
rect 1993 2333 2007 2347
rect 1893 2254 1907 2268
rect 1953 2293 1967 2307
rect 2013 2313 2027 2327
rect 2113 2493 2127 2507
rect 2093 2432 2107 2446
rect 2193 2474 2207 2488
rect 2413 2952 2427 2966
rect 2472 2953 2486 2967
rect 2493 2952 2507 2966
rect 2893 5413 2907 5427
rect 2853 5374 2867 5388
rect 3053 5594 3067 5608
rect 3093 5593 3107 5607
rect 2953 5533 2967 5547
rect 3073 5552 3087 5566
rect 3033 5513 3047 5527
rect 2973 5493 2987 5507
rect 2833 5233 2847 5247
rect 2873 5333 2887 5347
rect 2853 5213 2867 5227
rect 2733 5133 2747 5147
rect 2793 5074 2807 5088
rect 2833 5074 2847 5088
rect 2893 5074 2907 5088
rect 2813 5032 2827 5046
rect 2872 5033 2886 5047
rect 2893 5033 2907 5047
rect 2773 4993 2787 5007
rect 2733 4893 2747 4907
rect 2813 4854 2827 4868
rect 2793 4812 2807 4826
rect 2813 4753 2827 4767
rect 2793 4713 2807 4727
rect 2773 4673 2787 4687
rect 2753 4613 2767 4627
rect 2833 4633 2847 4647
rect 2853 4613 2867 4627
rect 2813 4593 2827 4607
rect 2853 4573 2867 4587
rect 2793 4512 2807 4526
rect 2833 4512 2847 4526
rect 2733 4373 2747 4387
rect 2793 4373 2807 4387
rect 2713 4353 2727 4367
rect 2693 4333 2707 4347
rect 2733 4334 2747 4348
rect 2713 4292 2727 4306
rect 2693 4253 2707 4267
rect 2753 4253 2767 4267
rect 2673 4093 2687 4107
rect 2653 4073 2667 4087
rect 2673 4053 2687 4067
rect 2713 4093 2727 4107
rect 2773 4093 2787 4107
rect 2653 3873 2667 3887
rect 2673 3853 2687 3867
rect 2553 3513 2567 3527
rect 2533 3333 2547 3347
rect 2613 3812 2627 3826
rect 2733 4053 2747 4067
rect 2713 3813 2727 3827
rect 2893 4953 2907 4967
rect 2933 5233 2947 5247
rect 3073 5473 3087 5487
rect 3013 5393 3027 5407
rect 3053 5393 3067 5407
rect 2993 5374 3007 5388
rect 2993 5253 3007 5267
rect 3133 5813 3147 5827
rect 3133 5552 3147 5566
rect 3113 5513 3127 5527
rect 3133 5493 3147 5507
rect 3173 6253 3187 6267
rect 3193 6213 3207 6227
rect 3473 6433 3487 6447
rect 3333 6414 3347 6428
rect 3373 6414 3387 6428
rect 3953 6433 3967 6447
rect 3993 6433 4007 6447
rect 3613 6414 3627 6428
rect 3753 6414 3767 6428
rect 3793 6414 3807 6428
rect 3313 6372 3327 6386
rect 3873 6413 3887 6427
rect 3913 6414 3927 6428
rect 3513 6393 3527 6407
rect 3453 6313 3467 6327
rect 3373 6253 3387 6267
rect 3333 6173 3347 6187
rect 3313 6153 3327 6167
rect 3273 6114 3287 6128
rect 3313 6114 3327 6128
rect 3172 6072 3186 6086
rect 3193 6073 3207 6087
rect 3253 6072 3267 6086
rect 3293 6013 3307 6027
rect 3213 5894 3227 5908
rect 3193 5852 3207 5866
rect 3233 5773 3247 5787
rect 3413 6114 3427 6128
rect 3393 5933 3407 5947
rect 3593 6372 3607 6386
rect 3633 6353 3647 6367
rect 3773 6372 3787 6386
rect 3933 6372 3947 6386
rect 4033 6413 4047 6427
rect 4093 6414 4107 6428
rect 3993 6353 4007 6367
rect 3733 6333 3747 6347
rect 3873 6333 3887 6347
rect 3973 6333 3987 6347
rect 3973 6193 3987 6207
rect 3893 6153 3907 6167
rect 3553 6114 3567 6128
rect 3593 6114 3607 6128
rect 3653 6114 3667 6128
rect 3513 5973 3527 5987
rect 3433 5913 3447 5927
rect 3353 5894 3367 5908
rect 3413 5893 3427 5907
rect 3293 5793 3307 5807
rect 3213 5594 3227 5608
rect 3173 5553 3187 5567
rect 3273 5552 3287 5566
rect 3313 5513 3327 5527
rect 3233 5493 3247 5507
rect 3193 5473 3207 5487
rect 3233 5472 3247 5486
rect 3173 5433 3187 5447
rect 3113 5332 3127 5346
rect 3073 5273 3087 5287
rect 3013 5233 3027 5247
rect 3053 5213 3067 5227
rect 2973 5173 2987 5187
rect 3013 5074 3027 5088
rect 2953 5032 2967 5046
rect 2993 4973 3007 4987
rect 2913 4893 2927 4907
rect 3033 4893 3047 4907
rect 2913 4854 2927 4868
rect 2973 4854 2987 4868
rect 2893 4733 2907 4747
rect 2893 4573 2907 4587
rect 2893 4552 2907 4566
rect 3013 4853 3027 4867
rect 2993 4673 3007 4687
rect 2973 4554 2987 4568
rect 3033 4713 3047 4727
rect 2913 4493 2927 4507
rect 2893 4473 2907 4487
rect 2993 4512 3007 4526
rect 2953 4493 2967 4507
rect 2933 4373 2947 4387
rect 2873 4333 2887 4347
rect 2913 4334 2927 4348
rect 2793 4053 2807 4067
rect 2973 4433 2987 4447
rect 2953 4253 2967 4267
rect 2933 4133 2947 4147
rect 2913 4053 2927 4067
rect 2813 3992 2827 4006
rect 2793 3933 2807 3947
rect 2693 3693 2707 3707
rect 2633 3653 2647 3667
rect 2773 3653 2787 3667
rect 2713 3613 2727 3627
rect 2613 3573 2627 3587
rect 2673 3573 2687 3587
rect 2633 3533 2647 3547
rect 2893 3992 2907 4006
rect 3153 5133 3167 5147
rect 3133 5074 3147 5088
rect 3153 5032 3167 5046
rect 3273 5374 3287 5388
rect 3253 5332 3267 5346
rect 3373 5852 3387 5866
rect 3413 5853 3427 5867
rect 3533 5913 3547 5927
rect 3453 5894 3467 5908
rect 3493 5894 3507 5908
rect 3353 5473 3367 5487
rect 3333 5373 3347 5387
rect 3313 5313 3327 5327
rect 3333 5293 3347 5307
rect 3253 5233 3267 5247
rect 3233 5193 3247 5207
rect 3213 5073 3227 5087
rect 3073 4853 3087 4867
rect 3113 4854 3127 4868
rect 3213 4973 3227 4987
rect 3193 4853 3207 4867
rect 3333 5173 3347 5187
rect 3433 5473 3447 5487
rect 3393 5413 3407 5427
rect 3373 5373 3387 5387
rect 3433 5374 3447 5388
rect 3393 5313 3407 5327
rect 3353 5153 3367 5167
rect 3333 5133 3347 5147
rect 3273 5113 3287 5127
rect 3313 5032 3327 5046
rect 3253 4893 3267 4907
rect 3373 4973 3387 4987
rect 3313 4873 3327 4887
rect 3073 4812 3087 4826
rect 3133 4812 3147 4826
rect 3093 4773 3107 4787
rect 3193 4773 3207 4787
rect 3053 4673 3067 4687
rect 3053 4593 3067 4607
rect 3053 4493 3067 4507
rect 3293 4854 3307 4868
rect 3353 4853 3367 4867
rect 3233 4833 3247 4847
rect 3273 4812 3287 4826
rect 3373 4812 3387 4826
rect 3353 4793 3367 4807
rect 3313 4773 3327 4787
rect 3373 4773 3387 4787
rect 3273 4733 3287 4747
rect 3353 4733 3367 4747
rect 3233 4653 3247 4667
rect 3113 4554 3127 4568
rect 3153 4554 3167 4568
rect 3213 4552 3227 4566
rect 3073 4473 3087 4487
rect 3133 4473 3147 4487
rect 3073 4413 3087 4427
rect 3113 4393 3127 4407
rect 3033 4373 3047 4387
rect 3053 4334 3067 4348
rect 3133 4353 3147 4367
rect 3073 4292 3087 4306
rect 3113 4292 3127 4306
rect 3373 4633 3387 4647
rect 3353 4613 3367 4627
rect 3353 4573 3367 4587
rect 3193 4393 3207 4407
rect 3293 4554 3307 4568
rect 3373 4512 3387 4526
rect 3313 4493 3327 4507
rect 3353 4493 3367 4507
rect 3613 6072 3627 6086
rect 3693 6113 3707 6127
rect 3753 6114 3767 6128
rect 3933 6114 3947 6128
rect 3653 6013 3667 6027
rect 3713 6072 3727 6086
rect 3773 6072 3787 6086
rect 3913 6072 3927 6086
rect 3953 6073 3967 6087
rect 3593 5973 3607 5987
rect 3693 5973 3707 5987
rect 3573 5733 3587 5747
rect 3673 5894 3687 5908
rect 3853 5894 3867 5908
rect 3653 5852 3667 5866
rect 3973 6013 3987 6027
rect 4273 6414 4287 6428
rect 4373 6413 4387 6427
rect 4473 6414 4487 6428
rect 4513 6413 4527 6427
rect 4613 6414 4627 6428
rect 4693 6413 4707 6427
rect 4753 6414 4767 6428
rect 5573 6433 5587 6447
rect 5993 6433 6007 6447
rect 4993 6414 5007 6428
rect 5073 6414 5087 6428
rect 5113 6414 5127 6428
rect 5153 6414 5167 6428
rect 5193 6414 5207 6428
rect 5253 6414 5267 6428
rect 5293 6414 5307 6428
rect 5453 6414 5467 6428
rect 4033 6313 4047 6327
rect 4213 6353 4227 6367
rect 4253 6353 4267 6367
rect 4373 6372 4387 6386
rect 4413 6372 4427 6386
rect 4453 6313 4467 6327
rect 4133 6293 4147 6307
rect 4293 6293 4307 6307
rect 4013 6253 4027 6267
rect 4073 6114 4087 6128
rect 4033 6073 4047 6087
rect 4333 6173 4347 6187
rect 4233 6153 4247 6167
rect 4293 6153 4307 6167
rect 4173 6113 4187 6127
rect 4313 6114 4327 6128
rect 4013 6033 4027 6047
rect 3993 5933 4007 5947
rect 4093 6033 4107 6047
rect 4053 5993 4067 6007
rect 4093 5893 4107 5907
rect 3953 5853 3967 5867
rect 4053 5852 4067 5866
rect 4033 5813 4047 5827
rect 3833 5793 3847 5807
rect 3653 5753 3667 5767
rect 3593 5673 3607 5687
rect 3573 5594 3587 5608
rect 3613 5594 3627 5608
rect 3593 5552 3607 5566
rect 3633 5553 3647 5567
rect 3553 5513 3567 5527
rect 3633 5493 3647 5507
rect 3613 5473 3627 5487
rect 3513 5373 3527 5387
rect 3573 5374 3587 5388
rect 3613 5373 3627 5387
rect 3513 5332 3527 5346
rect 3553 5332 3567 5346
rect 3593 5333 3607 5347
rect 3633 5333 3647 5347
rect 3473 5313 3487 5327
rect 3533 5293 3547 5307
rect 3413 5273 3427 5287
rect 3433 5253 3447 5267
rect 3433 5193 3447 5207
rect 3473 5074 3487 5088
rect 3493 4993 3507 5007
rect 3593 5233 3607 5247
rect 3633 5133 3647 5147
rect 3573 5093 3587 5107
rect 3833 5733 3847 5747
rect 3773 5713 3787 5727
rect 3673 5594 3687 5608
rect 3733 5594 3747 5608
rect 3813 5693 3827 5707
rect 3813 5594 3827 5608
rect 3673 5553 3687 5567
rect 3753 5552 3767 5566
rect 3713 5513 3727 5527
rect 3953 5653 3967 5667
rect 3913 5594 3927 5608
rect 3833 5473 3847 5487
rect 3713 5433 3727 5447
rect 3793 5433 3807 5447
rect 3753 5393 3767 5407
rect 3773 5373 3787 5387
rect 3693 5332 3707 5346
rect 3753 5333 3767 5347
rect 3733 5193 3747 5207
rect 3653 5093 3667 5107
rect 3693 5074 3707 5088
rect 3573 5032 3587 5046
rect 3653 5032 3667 5046
rect 3453 4933 3467 4947
rect 3553 4933 3567 4947
rect 3673 4933 3687 4947
rect 3433 4873 3447 4887
rect 3553 4873 3567 4887
rect 3613 4873 3627 4887
rect 3473 4854 3487 4868
rect 3513 4854 3527 4868
rect 3453 4812 3467 4826
rect 3513 4733 3527 4747
rect 3453 4693 3467 4707
rect 3413 4673 3427 4687
rect 3413 4573 3427 4587
rect 3513 4613 3527 4627
rect 3393 4473 3407 4487
rect 3473 4512 3487 4526
rect 3633 4854 3647 4868
rect 3973 5553 3987 5567
rect 4093 5793 4107 5807
rect 4093 5693 4107 5707
rect 4173 6072 4187 6086
rect 4213 6072 4227 6086
rect 4253 6072 4267 6086
rect 4293 6072 4307 6086
rect 4593 6372 4607 6386
rect 4633 6293 4647 6307
rect 4673 6233 4687 6247
rect 4393 6114 4407 6128
rect 4513 6112 4527 6126
rect 4553 6114 4567 6128
rect 4593 6114 4607 6128
rect 4633 6114 4647 6128
rect 4413 6072 4427 6086
rect 4473 6072 4487 6086
rect 4313 6053 4327 6067
rect 4373 6053 4387 6067
rect 4133 5993 4147 6007
rect 4173 5973 4187 5987
rect 4253 5933 4267 5947
rect 4293 5933 4307 5947
rect 4173 5894 4187 5908
rect 4193 5852 4207 5866
rect 4153 5773 4167 5787
rect 4133 5693 4147 5707
rect 4113 5673 4127 5687
rect 4093 5594 4107 5608
rect 3933 5473 3947 5487
rect 3893 5433 3907 5447
rect 3833 5374 3847 5388
rect 3873 5374 3887 5388
rect 3813 5333 3827 5347
rect 3793 5193 3807 5207
rect 3893 5333 3907 5347
rect 3893 5233 3907 5247
rect 3853 5173 3867 5187
rect 3813 5153 3827 5167
rect 3773 5113 3787 5127
rect 3873 5113 3887 5127
rect 3793 5074 3807 5088
rect 3833 5074 3847 5088
rect 3733 5032 3747 5046
rect 3773 5032 3787 5046
rect 3853 4993 3867 5007
rect 3813 4933 3827 4947
rect 3693 4913 3707 4927
rect 3813 4912 3827 4926
rect 3773 4893 3787 4907
rect 3613 4793 3627 4807
rect 3673 4773 3687 4787
rect 3553 4693 3567 4707
rect 3653 4693 3667 4707
rect 3673 4673 3687 4687
rect 3613 4633 3627 4647
rect 3553 4573 3567 4587
rect 3453 4473 3467 4487
rect 3293 4413 3307 4427
rect 3433 4413 3447 4427
rect 3153 4293 3167 4307
rect 3193 4292 3207 4306
rect 3233 4292 3247 4306
rect 3033 4273 3047 4287
rect 3133 4273 3147 4287
rect 2993 4233 3007 4247
rect 3053 4233 3067 4247
rect 2973 4073 2987 4087
rect 2993 4034 3007 4048
rect 3033 4034 3047 4048
rect 2933 3992 2947 4006
rect 2973 3992 2987 4006
rect 2913 3933 2927 3947
rect 2993 3933 3007 3947
rect 2853 3893 2867 3907
rect 2813 3853 2827 3867
rect 2873 3814 2887 3828
rect 2913 3814 2927 3828
rect 2953 3814 2967 3828
rect 2893 3772 2907 3786
rect 3033 3873 3047 3887
rect 3113 4193 3127 4207
rect 3073 4113 3087 4127
rect 3213 4233 3227 4247
rect 3193 4133 3207 4147
rect 3133 4053 3147 4067
rect 3073 3993 3087 4007
rect 3133 3992 3147 4006
rect 3313 4393 3327 4407
rect 3373 4353 3387 4367
rect 3413 4334 3427 4348
rect 3313 4293 3327 4307
rect 3293 4253 3307 4267
rect 3433 4293 3447 4307
rect 3393 4253 3407 4267
rect 3353 4233 3367 4247
rect 3433 4193 3447 4207
rect 3533 4513 3547 4527
rect 3893 5072 3907 5086
rect 3893 5013 3907 5027
rect 3873 4933 3887 4947
rect 3713 4813 3727 4827
rect 3693 4573 3707 4587
rect 3653 4554 3667 4568
rect 3553 4473 3567 4487
rect 3573 4353 3587 4367
rect 3533 4334 3547 4348
rect 3793 4812 3807 4826
rect 3733 4733 3747 4747
rect 3953 5433 3967 5447
rect 4033 5552 4047 5566
rect 4073 5552 4087 5566
rect 3993 5493 4007 5507
rect 4033 5513 4047 5527
rect 4013 5413 4027 5427
rect 3973 5373 3987 5387
rect 4093 5473 4107 5487
rect 4033 5393 4047 5407
rect 4093 5373 4107 5387
rect 4273 5793 4287 5807
rect 4213 5753 4227 5767
rect 4253 5753 4267 5767
rect 4333 5894 4347 5908
rect 4453 6013 4467 6027
rect 4413 5894 4427 5908
rect 4313 5853 4327 5867
rect 4573 6072 4587 6086
rect 4773 6273 4787 6287
rect 4813 6213 4827 6227
rect 4853 6213 4867 6227
rect 4713 6173 4727 6187
rect 4773 6173 4787 6187
rect 4693 6114 4707 6128
rect 4613 6053 4627 6067
rect 4673 6053 4687 6067
rect 4513 6013 4527 6027
rect 4693 5993 4707 6007
rect 4493 5973 4507 5987
rect 4533 5973 4547 5987
rect 4473 5894 4487 5908
rect 4353 5852 4367 5866
rect 4393 5852 4407 5866
rect 4453 5852 4467 5866
rect 4312 5813 4326 5827
rect 4333 5813 4347 5827
rect 4633 5933 4647 5947
rect 4573 5913 4587 5927
rect 4613 5913 4627 5927
rect 4493 5853 4507 5867
rect 4553 5852 4567 5866
rect 4533 5773 4547 5787
rect 4473 5733 4487 5747
rect 4293 5713 4307 5727
rect 4193 5693 4207 5707
rect 4413 5673 4427 5687
rect 4313 5653 4327 5667
rect 4193 5633 4207 5647
rect 4173 5613 4187 5627
rect 4193 5593 4207 5607
rect 4253 5594 4267 5608
rect 4413 5614 4427 5628
rect 4413 5593 4427 5607
rect 4453 5594 4467 5608
rect 4493 5594 4507 5608
rect 4193 5552 4207 5566
rect 4233 5552 4247 5566
rect 4273 5552 4287 5566
rect 4313 5552 4327 5566
rect 4433 5552 4447 5566
rect 4473 5513 4487 5527
rect 4393 5493 4407 5507
rect 4153 5473 4167 5487
rect 4253 5473 4267 5487
rect 4153 5433 4167 5447
rect 4193 5433 4207 5447
rect 3993 5332 4007 5346
rect 4033 5332 4047 5346
rect 4113 5332 4127 5346
rect 3953 5253 3967 5267
rect 4013 5213 4027 5227
rect 3973 5173 3987 5187
rect 3933 5133 3947 5147
rect 3933 5073 3947 5087
rect 3973 5074 3987 5088
rect 4213 5293 4227 5307
rect 4233 5213 4247 5227
rect 4173 5173 4187 5187
rect 4213 5173 4227 5187
rect 4053 5153 4067 5167
rect 3953 5013 3967 5027
rect 4033 5033 4047 5047
rect 4013 5013 4027 5027
rect 3953 4992 3967 5006
rect 3993 4993 4007 5007
rect 3913 4893 3927 4907
rect 4013 4973 4027 4987
rect 4013 4933 4027 4947
rect 4013 4853 4027 4867
rect 3893 4812 3907 4826
rect 4073 5133 4087 5147
rect 4053 4933 4067 4947
rect 3933 4812 3947 4826
rect 3973 4812 3987 4826
rect 4033 4812 4047 4826
rect 4033 4753 4047 4767
rect 3892 4713 3906 4727
rect 3913 4713 3927 4727
rect 3873 4633 3887 4647
rect 3793 4613 3807 4627
rect 3873 4573 3887 4587
rect 3833 4554 3847 4568
rect 3733 4512 3747 4526
rect 3613 4473 3627 4487
rect 3593 4333 3607 4347
rect 3493 4293 3507 4307
rect 3553 4292 3567 4306
rect 3593 4293 3607 4307
rect 3472 4253 3486 4267
rect 3493 4253 3507 4267
rect 3473 4193 3487 4207
rect 3413 4173 3427 4187
rect 3453 4173 3467 4187
rect 3293 4073 3307 4087
rect 3333 4053 3347 4067
rect 3372 4053 3386 4067
rect 3393 4053 3407 4067
rect 3133 3953 3147 3967
rect 3033 3833 3047 3847
rect 3073 3814 3087 3828
rect 3093 3772 3107 3786
rect 3173 3793 3187 3807
rect 3073 3733 3087 3747
rect 2913 3713 2927 3727
rect 2953 3713 2967 3727
rect 3053 3713 3067 3727
rect 3073 3693 3087 3707
rect 2913 3653 2927 3667
rect 2853 3613 2867 3627
rect 2813 3553 2827 3567
rect 2893 3553 2907 3567
rect 2733 3533 2747 3547
rect 2573 3294 2587 3308
rect 2713 3473 2727 3487
rect 2653 3453 2667 3467
rect 2793 3532 2807 3546
rect 2833 3514 2847 3528
rect 2813 3472 2827 3486
rect 2853 3472 2867 3486
rect 2893 3472 2907 3486
rect 2753 3453 2767 3467
rect 2733 3413 2747 3427
rect 2853 3373 2867 3387
rect 2653 3333 2667 3347
rect 2733 3294 2747 3308
rect 2773 3294 2787 3308
rect 2813 3294 2827 3308
rect 2553 3133 2567 3147
rect 2793 3252 2807 3266
rect 2733 3233 2747 3247
rect 2693 3193 2707 3207
rect 2633 3113 2647 3127
rect 2653 3073 2667 3087
rect 2593 2994 2607 3008
rect 2493 2774 2507 2788
rect 2573 2952 2587 2966
rect 2593 2833 2607 2847
rect 2333 2653 2347 2667
rect 2273 2474 2287 2488
rect 2193 2433 2207 2447
rect 2093 2393 2107 2407
rect 2153 2393 2167 2407
rect 2073 2313 2087 2327
rect 2033 2273 2047 2287
rect 2053 2253 2067 2267
rect 1893 2212 1907 2226
rect 1973 2212 1987 2226
rect 1933 2153 1947 2167
rect 1813 1913 1827 1927
rect 1893 1893 1907 1907
rect 1673 1734 1687 1748
rect 1693 1692 1707 1706
rect 1653 1653 1667 1667
rect 1613 1493 1627 1507
rect 1633 1453 1647 1467
rect 1793 1734 1807 1748
rect 1813 1692 1827 1706
rect 1893 1734 1907 1748
rect 1873 1673 1887 1687
rect 1753 1653 1767 1667
rect 1713 1593 1727 1607
rect 1713 1553 1727 1567
rect 1613 1392 1627 1406
rect 1693 1393 1707 1407
rect 1613 1353 1627 1367
rect 1693 1273 1707 1287
rect 1953 1993 1967 2007
rect 2052 2212 2066 2226
rect 2073 2212 2087 2226
rect 2013 2173 2027 2187
rect 2153 2254 2167 2268
rect 2233 2253 2247 2267
rect 2133 2212 2147 2226
rect 2173 2212 2187 2226
rect 2233 2212 2247 2226
rect 2173 2173 2187 2187
rect 2293 2432 2307 2446
rect 2473 2653 2487 2667
rect 2493 2633 2507 2647
rect 2573 2732 2587 2746
rect 2513 2593 2527 2607
rect 2493 2573 2507 2587
rect 2393 2553 2407 2567
rect 2373 2513 2387 2527
rect 2353 2433 2367 2447
rect 2533 2513 2547 2527
rect 2393 2493 2407 2507
rect 2473 2493 2487 2507
rect 2393 2333 2407 2347
rect 2373 2293 2387 2307
rect 2333 2273 2347 2287
rect 2313 2254 2327 2268
rect 2273 2173 2287 2187
rect 2153 2133 2167 2147
rect 2253 2133 2267 2147
rect 2093 2093 2107 2107
rect 2053 1973 2067 1987
rect 2013 1954 2027 1968
rect 2113 1954 2127 1968
rect 1953 1833 1967 1847
rect 2113 1913 2127 1927
rect 2193 2093 2207 2107
rect 2233 1954 2247 1968
rect 2213 1912 2227 1926
rect 2073 1893 2087 1907
rect 2153 1893 2167 1907
rect 2173 1853 2187 1867
rect 2053 1833 2067 1847
rect 2033 1813 2047 1827
rect 1933 1773 1947 1787
rect 2033 1773 2047 1787
rect 1973 1734 1987 1748
rect 2013 1733 2027 1747
rect 1913 1693 1927 1707
rect 1953 1673 1967 1687
rect 1773 1493 1787 1507
rect 1893 1493 1907 1507
rect 2013 1633 2027 1647
rect 2113 1734 2127 1748
rect 2213 1833 2227 1847
rect 2173 1714 2187 1728
rect 2053 1692 2067 1706
rect 2093 1692 2107 1706
rect 2073 1633 2087 1647
rect 1973 1513 1987 1527
rect 2033 1513 2047 1527
rect 1953 1473 1967 1487
rect 1813 1434 1827 1448
rect 1853 1434 1867 1448
rect 1893 1434 1907 1448
rect 1933 1434 1947 1448
rect 2033 1473 2047 1487
rect 1713 1253 1727 1267
rect 1793 1392 1807 1406
rect 1853 1353 1867 1367
rect 1633 1172 1647 1186
rect 1553 1153 1567 1167
rect 1593 1153 1607 1167
rect 1633 1013 1647 1027
rect 1573 953 1587 967
rect 1533 913 1547 927
rect 1553 872 1567 886
rect 1653 953 1667 967
rect 1633 833 1647 847
rect 1573 694 1587 708
rect 1753 1233 1767 1247
rect 1813 1233 1827 1247
rect 1873 1233 1887 1247
rect 1693 1214 1707 1228
rect 1773 1214 1787 1228
rect 1713 1172 1727 1186
rect 1753 1172 1767 1186
rect 1693 1093 1707 1107
rect 1833 1133 1847 1147
rect 1793 1093 1807 1107
rect 1813 973 1827 987
rect 1753 953 1767 967
rect 1713 914 1727 928
rect 1773 872 1787 886
rect 1733 833 1747 847
rect 1793 833 1807 847
rect 1713 813 1727 827
rect 1753 813 1767 827
rect 1793 773 1807 787
rect 1713 733 1727 747
rect 1773 733 1787 747
rect 1593 652 1607 666
rect 1633 652 1647 666
rect 1673 652 1687 666
rect 1673 533 1687 547
rect 1533 513 1547 527
rect 1533 453 1547 467
rect 1593 394 1607 408
rect 1833 914 1847 928
rect 1993 1392 2007 1406
rect 2033 1392 2047 1406
rect 1953 1333 1967 1347
rect 1993 1253 2007 1267
rect 1953 1214 1967 1228
rect 2053 1213 2067 1227
rect 2153 1693 2167 1707
rect 2153 1653 2167 1667
rect 2133 1613 2147 1627
rect 2113 1473 2127 1487
rect 2153 1513 2167 1527
rect 2193 1513 2207 1527
rect 2133 1453 2147 1467
rect 2153 1434 2167 1448
rect 2133 1353 2147 1367
rect 2093 1313 2107 1327
rect 2073 1172 2087 1186
rect 2113 1273 2127 1287
rect 2193 1373 2207 1387
rect 2173 1313 2187 1327
rect 2193 1273 2207 1287
rect 2133 1253 2147 1267
rect 2113 1233 2127 1247
rect 2153 1214 2167 1228
rect 2233 1733 2247 1747
rect 2233 1653 2247 1667
rect 2333 2212 2347 2226
rect 2493 2353 2507 2367
rect 2393 2254 2407 2268
rect 2433 2254 2447 2268
rect 2512 2333 2526 2347
rect 2533 2333 2547 2347
rect 2513 2233 2527 2247
rect 2453 2212 2467 2226
rect 2393 2173 2407 2187
rect 2293 2093 2307 2107
rect 2593 2632 2607 2646
rect 2573 2293 2587 2307
rect 2533 2133 2547 2147
rect 2673 3033 2687 3047
rect 2673 2893 2687 2907
rect 2653 2873 2667 2887
rect 2833 3133 2847 3147
rect 2773 3113 2787 3127
rect 2733 2994 2747 3008
rect 2753 2952 2767 2966
rect 2793 2933 2807 2947
rect 2693 2853 2707 2867
rect 2673 2833 2687 2847
rect 2773 2833 2787 2847
rect 2653 2732 2667 2746
rect 2933 3613 2947 3627
rect 3053 3593 3067 3607
rect 3033 3533 3047 3547
rect 2993 3514 3007 3528
rect 2933 3472 2947 3486
rect 2973 3472 2987 3486
rect 3033 3473 3047 3487
rect 2993 3413 3007 3427
rect 2913 3294 2927 3308
rect 2953 3294 2967 3308
rect 3133 3772 3147 3786
rect 3233 3992 3247 4006
rect 3313 3992 3327 4006
rect 3293 3953 3307 3967
rect 3253 3833 3267 3847
rect 3233 3814 3247 3828
rect 3373 3913 3387 3927
rect 3353 3833 3367 3847
rect 3533 4113 3547 4127
rect 3633 4413 3647 4427
rect 3653 4353 3667 4367
rect 3693 4413 3707 4427
rect 3672 4333 3686 4347
rect 3693 4334 3707 4348
rect 3673 4293 3687 4307
rect 3653 4233 3667 4247
rect 3633 4133 3647 4147
rect 3613 4073 3627 4087
rect 3593 4053 3607 4067
rect 3713 4233 3727 4247
rect 3693 4093 3707 4107
rect 3453 3992 3467 4006
rect 3493 3992 3507 4006
rect 3533 3992 3547 4006
rect 3433 3873 3447 3887
rect 3773 4512 3787 4526
rect 3813 4512 3827 4526
rect 3913 4653 3927 4667
rect 3893 4533 3907 4547
rect 3873 4453 3887 4467
rect 3793 4433 3807 4447
rect 3773 4333 3787 4347
rect 3773 4193 3787 4207
rect 3853 4334 3867 4348
rect 3833 4292 3847 4306
rect 3873 4292 3887 4306
rect 3813 4193 3827 4207
rect 3793 4093 3807 4107
rect 3773 4073 3787 4087
rect 3753 4033 3767 4047
rect 3953 4593 3967 4607
rect 3993 4593 4007 4607
rect 3953 4493 3967 4507
rect 3933 4393 3947 4407
rect 3933 4292 3947 4306
rect 3933 4213 3947 4227
rect 3913 4113 3927 4127
rect 3873 4053 3887 4067
rect 3793 3953 3807 3967
rect 3693 3933 3707 3947
rect 3833 3893 3847 3907
rect 3553 3853 3567 3867
rect 3633 3853 3647 3867
rect 3413 3833 3427 3847
rect 3493 3833 3507 3847
rect 3193 3753 3207 3767
rect 3233 3713 3247 3727
rect 3213 3693 3227 3707
rect 3213 3653 3227 3667
rect 3073 3533 3087 3547
rect 3113 3533 3127 3547
rect 3173 3533 3187 3547
rect 3053 3373 3067 3387
rect 3033 3333 3047 3347
rect 2933 3252 2947 3266
rect 2933 3133 2947 3147
rect 2973 3113 2987 3127
rect 2933 3013 2947 3027
rect 2973 3013 2987 3027
rect 2853 2992 2867 3006
rect 2913 2994 2927 3008
rect 2833 2853 2847 2867
rect 2813 2833 2827 2847
rect 2893 2952 2907 2966
rect 2933 2873 2947 2887
rect 2913 2833 2927 2847
rect 2853 2813 2867 2827
rect 2813 2774 2827 2788
rect 2873 2774 2887 2788
rect 2793 2732 2807 2746
rect 2693 2693 2707 2707
rect 2893 2732 2907 2746
rect 2953 2733 2967 2747
rect 2873 2653 2887 2667
rect 2813 2553 2827 2567
rect 2933 2573 2947 2587
rect 2933 2513 2947 2527
rect 2673 2474 2687 2488
rect 2713 2432 2727 2446
rect 2873 2474 2887 2488
rect 2913 2474 2927 2488
rect 2993 2993 3007 3007
rect 3053 3293 3067 3307
rect 3053 3252 3067 3266
rect 3133 3514 3147 3528
rect 3293 3633 3307 3647
rect 3253 3553 3267 3567
rect 3113 3472 3127 3486
rect 3153 3472 3167 3486
rect 3192 3473 3193 3486
rect 3193 3473 3206 3486
rect 3213 3473 3227 3487
rect 3192 3472 3206 3473
rect 3133 3453 3147 3467
rect 3213 3452 3227 3466
rect 3333 3793 3347 3807
rect 3333 3733 3347 3747
rect 3393 3813 3407 3827
rect 3473 3813 3487 3827
rect 3413 3772 3427 3786
rect 3393 3753 3407 3767
rect 3353 3553 3367 3567
rect 3313 3533 3327 3547
rect 3273 3473 3287 3487
rect 3353 3472 3367 3486
rect 3313 3453 3327 3467
rect 3273 3413 3287 3427
rect 3353 3393 3367 3407
rect 3253 3333 3267 3347
rect 3313 3333 3327 3347
rect 3153 3294 3167 3308
rect 3233 3273 3247 3287
rect 3133 3252 3147 3266
rect 3193 3233 3207 3247
rect 3073 3173 3087 3187
rect 3173 3113 3187 3127
rect 3033 2993 3047 3007
rect 3013 2913 3027 2927
rect 3093 2952 3107 2966
rect 3173 2994 3187 3008
rect 3093 2913 3107 2927
rect 3053 2873 3067 2887
rect 3073 2833 3087 2847
rect 2993 2774 3007 2788
rect 3053 2774 3067 2788
rect 3153 2912 3167 2926
rect 3113 2873 3127 2887
rect 3353 3294 3367 3308
rect 3253 3252 3267 3266
rect 3293 3252 3307 3266
rect 3333 3233 3347 3247
rect 3433 3733 3447 3747
rect 3413 3453 3427 3467
rect 3593 3814 3607 3828
rect 3513 3793 3527 3807
rect 3493 3773 3507 3787
rect 3473 3653 3487 3667
rect 3473 3613 3487 3627
rect 3633 3773 3647 3787
rect 3573 3753 3587 3767
rect 3673 3813 3687 3827
rect 3733 3814 3747 3828
rect 3773 3814 3787 3828
rect 3713 3772 3727 3786
rect 3613 3653 3627 3667
rect 3513 3593 3527 3607
rect 3573 3492 3587 3506
rect 3453 3473 3467 3487
rect 3433 3393 3447 3407
rect 3433 3333 3447 3347
rect 3393 3213 3407 3227
rect 3493 3453 3507 3467
rect 3593 3433 3607 3447
rect 3533 3413 3547 3427
rect 3513 3333 3527 3347
rect 3473 3294 3487 3308
rect 3573 3252 3587 3266
rect 3353 3193 3367 3207
rect 3433 3193 3447 3207
rect 3413 3133 3427 3147
rect 3513 3133 3527 3147
rect 3413 3053 3427 3067
rect 3233 2994 3247 3008
rect 3273 2994 3287 3008
rect 3353 2993 3367 3007
rect 3433 2994 3447 3008
rect 3472 2994 3486 3008
rect 3493 2994 3507 3008
rect 3193 2953 3207 2967
rect 3293 2953 3307 2967
rect 3213 2933 3227 2947
rect 3253 2933 3267 2947
rect 3293 2893 3307 2907
rect 3453 2933 3467 2947
rect 3413 2913 3427 2927
rect 3453 2873 3467 2887
rect 3353 2853 3367 2867
rect 3433 2853 3447 2867
rect 3173 2833 3187 2847
rect 3133 2813 3147 2827
rect 3193 2813 3207 2827
rect 3353 2813 3367 2827
rect 3113 2733 3127 2747
rect 3093 2653 3107 2667
rect 3093 2513 3107 2527
rect 2993 2493 3007 2507
rect 2973 2474 2987 2488
rect 3033 2474 3047 2488
rect 2853 2432 2867 2446
rect 2613 2333 2627 2347
rect 2753 2333 2767 2347
rect 2953 2432 2967 2446
rect 2973 2373 2987 2387
rect 2973 2333 2987 2347
rect 2933 2293 2947 2307
rect 2893 2254 2907 2268
rect 2733 2213 2747 2227
rect 2593 2093 2607 2107
rect 2673 2093 2687 2107
rect 2533 2033 2547 2047
rect 2413 1993 2427 2007
rect 2313 1953 2327 1967
rect 2353 1954 2367 1968
rect 2313 1893 2327 1907
rect 2453 1953 2467 1967
rect 2513 1954 2527 1968
rect 2933 2213 2947 2227
rect 3113 2313 3127 2327
rect 3073 2293 3087 2307
rect 3033 2254 3047 2268
rect 3313 2774 3327 2788
rect 3173 2732 3187 2746
rect 3553 3053 3567 3067
rect 3673 3693 3687 3707
rect 3653 3673 3667 3687
rect 3633 3613 3647 3627
rect 3793 3772 3807 3786
rect 3753 3633 3767 3647
rect 3853 3873 3867 3887
rect 3853 3733 3867 3747
rect 4013 4493 4027 4507
rect 4053 4673 4067 4687
rect 4033 4433 4047 4447
rect 4013 4413 4027 4427
rect 3973 4333 3987 4347
rect 4053 4333 4067 4347
rect 3993 4292 4007 4306
rect 3953 4173 3967 4187
rect 3973 4073 3987 4087
rect 4013 4034 4027 4048
rect 4093 5073 4107 5087
rect 4153 5074 4167 5088
rect 4093 5032 4107 5046
rect 4133 5032 4147 5046
rect 4173 5032 4187 5046
rect 4113 4873 4127 4887
rect 4133 4854 4147 4868
rect 4173 4853 4187 4867
rect 4093 4733 4107 4747
rect 4153 4733 4167 4747
rect 4133 4613 4147 4627
rect 4093 4573 4107 4587
rect 4293 5433 4307 5447
rect 4353 5393 4367 5407
rect 4473 5453 4487 5467
rect 4453 5353 4467 5367
rect 4293 5332 4307 5346
rect 4373 5332 4387 5346
rect 4333 5293 4347 5307
rect 4593 5813 4607 5827
rect 4613 5733 4627 5747
rect 4593 5613 4607 5627
rect 4573 5594 4587 5608
rect 4673 5973 4687 5987
rect 4773 6152 4787 6166
rect 4813 6153 4827 6167
rect 4833 6133 4847 6147
rect 4793 6072 4807 6086
rect 4833 6072 4847 6086
rect 4713 5933 4727 5947
rect 4693 5894 4707 5908
rect 4813 6033 4827 6047
rect 4673 5853 4687 5867
rect 4653 5833 4667 5847
rect 4713 5852 4727 5866
rect 4753 5853 4767 5867
rect 4693 5833 4707 5847
rect 4753 5793 4767 5807
rect 4673 5773 4687 5787
rect 4693 5733 4707 5747
rect 4493 5413 4507 5427
rect 4593 5552 4607 5566
rect 4613 5533 4627 5547
rect 4573 5473 4587 5487
rect 4553 5393 4567 5407
rect 4533 5374 4547 5388
rect 4593 5374 4607 5388
rect 4593 5333 4607 5347
rect 4493 5293 4507 5307
rect 4473 5173 4487 5187
rect 4253 5113 4267 5127
rect 4313 5074 4327 5088
rect 4353 5074 4367 5088
rect 4593 5153 4607 5167
rect 4513 5133 4527 5147
rect 4573 5133 4587 5147
rect 4553 5093 4567 5107
rect 4253 5053 4267 5067
rect 4233 5032 4247 5046
rect 4253 4993 4267 5007
rect 4333 5032 4347 5046
rect 4493 5032 4507 5046
rect 4473 5013 4487 5027
rect 4453 4993 4467 5007
rect 4413 4973 4427 4987
rect 4413 4933 4427 4947
rect 4293 4913 4307 4927
rect 4293 4874 4307 4888
rect 4273 4853 4287 4867
rect 4313 4854 4327 4868
rect 4233 4813 4247 4827
rect 4213 4753 4227 4767
rect 4173 4573 4187 4587
rect 4213 4593 4227 4607
rect 4193 4553 4207 4567
rect 4113 4512 4127 4526
rect 4153 4512 4167 4526
rect 4193 4453 4207 4467
rect 4153 4433 4167 4447
rect 4113 4393 4127 4407
rect 4093 4373 4107 4387
rect 4073 4213 4087 4227
rect 4073 4173 4087 4187
rect 4053 4013 4067 4027
rect 3993 3973 4007 3987
rect 3953 3933 3967 3947
rect 4013 3913 4027 3927
rect 3913 3873 3927 3887
rect 3873 3673 3887 3687
rect 3933 3653 3947 3667
rect 3833 3613 3847 3627
rect 3913 3613 3927 3627
rect 3653 3533 3667 3547
rect 3633 3333 3647 3347
rect 3633 3293 3647 3307
rect 3673 3494 3687 3508
rect 3813 3494 3827 3508
rect 4053 3873 4067 3887
rect 4333 4812 4347 4826
rect 4293 4773 4307 4787
rect 4253 4633 4267 4647
rect 4233 4554 4247 4568
rect 4213 4413 4227 4427
rect 4233 4333 4247 4347
rect 4133 4293 4147 4307
rect 4113 4233 4127 4247
rect 4093 4153 4107 4167
rect 4093 4113 4107 4127
rect 4173 4292 4187 4306
rect 4213 4233 4227 4247
rect 4193 4153 4207 4167
rect 4133 4093 4147 4107
rect 4133 4053 4147 4067
rect 4093 3993 4107 4007
rect 4153 3992 4167 4006
rect 4073 3833 4087 3847
rect 4093 3814 4107 3828
rect 4113 3772 4127 3786
rect 4073 3693 4087 3707
rect 3973 3534 3987 3548
rect 4013 3534 4027 3548
rect 3933 3492 3947 3506
rect 3913 3373 3927 3387
rect 3993 3373 4007 3387
rect 3673 3333 3687 3347
rect 3713 3293 3727 3307
rect 3633 3233 3647 3247
rect 3613 3213 3627 3227
rect 4073 3613 4087 3627
rect 4073 3513 4087 3527
rect 4053 3493 4067 3507
rect 4073 3473 4087 3487
rect 4053 3453 4067 3467
rect 4113 3713 4127 3727
rect 4173 3633 4187 3647
rect 4113 3593 4127 3607
rect 4373 4773 4387 4787
rect 4353 4713 4367 4727
rect 4373 4692 4387 4706
rect 4333 4653 4347 4667
rect 4293 4593 4307 4607
rect 4293 4554 4307 4568
rect 4313 4512 4327 4526
rect 4433 4913 4447 4927
rect 4413 4773 4427 4787
rect 4473 4933 4487 4947
rect 4493 4854 4507 4868
rect 4473 4812 4487 4826
rect 4513 4773 4527 4787
rect 4473 4713 4487 4727
rect 4433 4693 4447 4707
rect 4413 4673 4427 4687
rect 4453 4673 4467 4687
rect 4413 4652 4427 4666
rect 4393 4573 4407 4587
rect 4393 4512 4407 4526
rect 4373 4473 4387 4487
rect 4293 4433 4307 4447
rect 4273 4333 4287 4347
rect 4353 4334 4367 4348
rect 4533 4733 4547 4747
rect 4513 4633 4527 4647
rect 4433 4593 4447 4607
rect 4453 4573 4467 4587
rect 4453 4473 4467 4487
rect 4433 4334 4447 4348
rect 4293 4293 4307 4307
rect 4333 4292 4347 4306
rect 4433 4293 4447 4307
rect 4293 4272 4307 4286
rect 4373 4273 4387 4287
rect 4213 4093 4227 4107
rect 4193 3573 4207 3587
rect 4273 4133 4287 4147
rect 4273 4053 4287 4067
rect 4313 4253 4327 4267
rect 4393 4153 4407 4167
rect 4313 4113 4327 4127
rect 4353 4053 4367 4067
rect 4373 4013 4387 4027
rect 4273 3992 4287 4006
rect 4353 3993 4367 4007
rect 4253 3913 4267 3927
rect 4233 3873 4247 3887
rect 4293 3814 4307 3828
rect 4273 3772 4287 3786
rect 4373 3913 4387 3927
rect 4373 3814 4387 3828
rect 4433 4093 4447 4107
rect 4513 4512 4527 4526
rect 4473 4453 4487 4467
rect 4533 4453 4547 4467
rect 4573 5032 4587 5046
rect 4573 4873 4587 4887
rect 4753 5653 4767 5667
rect 4793 5633 4807 5647
rect 4773 5613 4787 5627
rect 4793 5593 4807 5607
rect 5093 6372 5107 6386
rect 4933 6313 4947 6327
rect 4933 6133 4947 6147
rect 5113 6173 5127 6187
rect 4993 6114 5007 6128
rect 5073 6114 5087 6128
rect 4873 6072 4887 6086
rect 4913 6072 4927 6086
rect 4873 6012 4887 6026
rect 4852 5993 4866 6007
rect 4833 5893 4847 5907
rect 5053 6053 5067 6067
rect 5173 6393 5187 6407
rect 5513 6413 5527 6427
rect 5193 6373 5207 6387
rect 5233 6313 5247 6327
rect 5313 6372 5327 6386
rect 5433 6372 5447 6386
rect 5493 6372 5507 6386
rect 5433 6333 5447 6347
rect 5273 6293 5287 6307
rect 5173 6273 5187 6287
rect 5313 6273 5327 6287
rect 5493 6273 5507 6287
rect 5193 6213 5207 6227
rect 5233 6213 5247 6227
rect 5173 6153 5187 6167
rect 5153 6053 5167 6067
rect 5093 6033 5107 6047
rect 5013 5953 5027 5967
rect 4853 5793 4867 5807
rect 4953 5893 4967 5907
rect 5013 5913 5027 5927
rect 4933 5773 4947 5787
rect 4893 5733 4907 5747
rect 5053 5894 5067 5908
rect 5113 5894 5127 5908
rect 5033 5852 5047 5866
rect 4973 5833 4987 5847
rect 5033 5793 5047 5807
rect 5073 5793 5087 5807
rect 5013 5773 5027 5787
rect 4953 5653 4967 5667
rect 4853 5633 4867 5647
rect 4733 5552 4747 5566
rect 4773 5552 4787 5566
rect 4813 5552 4827 5566
rect 4693 5533 4707 5547
rect 4673 5493 4687 5507
rect 4813 5493 4827 5507
rect 4693 5433 4707 5447
rect 4793 5393 4807 5407
rect 4733 5374 4747 5388
rect 4773 5374 4787 5388
rect 4673 5332 4687 5346
rect 4673 5293 4687 5307
rect 4733 5293 4747 5307
rect 4653 5213 4667 5227
rect 4633 5093 4647 5107
rect 4613 5073 4627 5087
rect 4693 5173 4707 5187
rect 4713 5113 4727 5127
rect 4633 5032 4647 5046
rect 4693 4953 4707 4967
rect 4693 4893 4707 4907
rect 4673 4873 4687 4887
rect 4633 4854 4647 4868
rect 4633 4773 4647 4787
rect 4593 4613 4607 4627
rect 4573 4533 4587 4547
rect 4653 4733 4667 4747
rect 4793 5292 4807 5306
rect 4753 5173 4767 5187
rect 4873 5593 4887 5607
rect 4953 5594 4967 5608
rect 5033 5733 5047 5747
rect 4913 5552 4927 5566
rect 4993 5533 5007 5547
rect 4893 5493 4907 5507
rect 4953 5493 4967 5507
rect 4853 5453 4867 5467
rect 4933 5433 4947 5447
rect 4853 5332 4867 5346
rect 4913 5332 4927 5346
rect 4853 5293 4867 5307
rect 4792 5153 4806 5167
rect 4813 5153 4827 5167
rect 4813 5032 4827 5046
rect 4773 5013 4787 5027
rect 4753 4973 4767 4987
rect 4813 4953 4827 4967
rect 4913 5273 4927 5287
rect 4873 5213 4887 5227
rect 4853 4913 4867 4927
rect 4813 4873 4827 4887
rect 4733 4813 4747 4827
rect 4633 4593 4647 4607
rect 4693 4593 4707 4607
rect 4653 4573 4667 4587
rect 4693 4554 4707 4568
rect 4593 4513 4607 4527
rect 4573 4473 4587 4487
rect 4553 4433 4567 4447
rect 4533 4413 4547 4427
rect 4513 4393 4527 4407
rect 4553 4393 4567 4407
rect 4533 4353 4547 4367
rect 4553 4334 4567 4348
rect 4593 4334 4607 4348
rect 4533 4292 4547 4306
rect 4593 4253 4607 4267
rect 4533 4173 4547 4187
rect 4513 4153 4527 4167
rect 4453 4053 4467 4067
rect 4433 4034 4447 4048
rect 4473 4034 4487 4048
rect 4633 4512 4647 4526
rect 4673 4512 4687 4526
rect 4633 4491 4647 4505
rect 4733 4453 4747 4467
rect 4693 4334 4707 4348
rect 4653 4293 4667 4307
rect 4793 4812 4807 4826
rect 4793 4791 4807 4805
rect 4793 4713 4807 4727
rect 4773 4613 4787 4627
rect 4733 4253 4747 4267
rect 4713 4233 4727 4247
rect 4653 4193 4667 4207
rect 4573 4053 4587 4067
rect 4533 3993 4547 4007
rect 4493 3973 4507 3987
rect 4453 3953 4467 3967
rect 4513 3953 4527 3967
rect 4493 3933 4507 3947
rect 4533 3933 4547 3947
rect 4493 3893 4507 3907
rect 4453 3853 4467 3867
rect 4533 3833 4547 3847
rect 4373 3773 4387 3787
rect 4353 3753 4367 3767
rect 4333 3733 4347 3747
rect 4313 3713 4327 3727
rect 4333 3653 4347 3667
rect 4253 3633 4267 3647
rect 4213 3514 4227 3528
rect 4113 3472 4127 3486
rect 4072 3413 4086 3427
rect 4093 3413 4107 3427
rect 4153 3413 4167 3427
rect 4033 3313 4047 3327
rect 3873 3273 3887 3287
rect 3713 3253 3727 3267
rect 3853 3253 3867 3267
rect 3653 3133 3667 3147
rect 3613 3053 3627 3067
rect 3593 3033 3607 3047
rect 3593 2994 3607 3008
rect 3693 3033 3707 3047
rect 3513 2953 3527 2967
rect 3613 2952 3627 2966
rect 3653 2953 3667 2967
rect 3733 2994 3747 3008
rect 3773 2994 3787 3008
rect 3833 2994 3847 3008
rect 3493 2913 3507 2927
rect 3573 2913 3587 2927
rect 3633 2853 3647 2867
rect 3473 2833 3487 2847
rect 3573 2833 3587 2847
rect 3473 2774 3487 2788
rect 3533 2774 3547 2788
rect 3613 2774 3627 2788
rect 3393 2593 3407 2607
rect 3173 2474 3187 2488
rect 3213 2474 3227 2488
rect 3333 2474 3347 2488
rect 3173 2373 3187 2387
rect 2973 2212 2987 2226
rect 3053 2212 3067 2226
rect 2893 2173 2907 2187
rect 3013 2173 3027 2187
rect 2953 2153 2967 2167
rect 2853 2033 2867 2047
rect 2733 1993 2747 2007
rect 2833 1993 2847 2007
rect 2633 1933 2647 1947
rect 2493 1893 2507 1907
rect 2373 1853 2387 1867
rect 2413 1853 2427 1867
rect 2453 1853 2467 1867
rect 2293 1833 2307 1847
rect 2413 1712 2427 1726
rect 2273 1573 2287 1587
rect 2353 1573 2367 1587
rect 2273 1434 2287 1448
rect 2533 1893 2547 1907
rect 2573 1893 2587 1907
rect 2553 1853 2567 1867
rect 2553 1712 2567 1726
rect 2553 1673 2567 1687
rect 2433 1513 2447 1527
rect 2513 1513 2527 1527
rect 2393 1473 2407 1487
rect 2373 1434 2387 1448
rect 2253 1393 2267 1407
rect 2233 1373 2247 1387
rect 2293 1392 2307 1406
rect 2353 1393 2367 1407
rect 2273 1373 2287 1387
rect 2253 1333 2267 1347
rect 2233 1253 2247 1267
rect 2213 1233 2227 1247
rect 2253 1213 2267 1227
rect 2133 1172 2147 1186
rect 2173 1172 2187 1186
rect 2233 1172 2247 1186
rect 2013 1133 2027 1147
rect 1933 1113 1947 1127
rect 1893 1013 1907 1027
rect 1893 914 1907 928
rect 2013 1092 2027 1106
rect 1993 1033 2007 1047
rect 1853 873 1867 887
rect 1913 872 1927 886
rect 1893 833 1907 847
rect 1853 793 1867 807
rect 1833 773 1847 787
rect 1833 693 1847 707
rect 2253 1133 2267 1147
rect 2133 953 2147 967
rect 2053 853 2067 867
rect 2013 833 2027 847
rect 2093 813 2107 827
rect 2053 793 2067 807
rect 2173 914 2187 928
rect 2233 914 2247 928
rect 2473 1473 2487 1487
rect 2513 1473 2527 1487
rect 2573 1473 2587 1487
rect 2413 1393 2427 1407
rect 2453 1392 2467 1406
rect 2393 1313 2407 1327
rect 2553 1333 2567 1347
rect 2373 1273 2387 1287
rect 2333 1214 2347 1228
rect 2373 1214 2387 1228
rect 2453 1293 2467 1307
rect 2493 1293 2507 1307
rect 2413 1214 2427 1228
rect 2353 1172 2367 1186
rect 2313 1093 2327 1107
rect 2313 1053 2327 1067
rect 2393 1053 2407 1067
rect 2333 1013 2347 1027
rect 2253 872 2267 886
rect 2313 873 2327 887
rect 2213 853 2227 867
rect 2173 813 2187 827
rect 2333 833 2347 847
rect 1953 773 1967 787
rect 1993 773 2007 787
rect 2073 773 2087 787
rect 2133 773 2147 787
rect 2213 773 2227 787
rect 1993 713 2007 727
rect 2033 713 2047 727
rect 1753 652 1767 666
rect 1853 652 1867 666
rect 1893 653 1907 667
rect 1933 652 1947 666
rect 1713 433 1727 447
rect 1673 393 1687 407
rect 2333 733 2347 747
rect 2233 672 2247 686
rect 2333 672 2347 686
rect 2513 1273 2527 1287
rect 2513 1233 2527 1247
rect 2693 1813 2707 1827
rect 2833 1933 2847 1947
rect 2953 1993 2967 2007
rect 3093 2153 3107 2167
rect 3093 2113 3107 2127
rect 3353 2432 3367 2446
rect 3393 2432 3407 2446
rect 3613 2693 3627 2707
rect 3553 2513 3567 2527
rect 3473 2474 3487 2488
rect 3513 2474 3527 2488
rect 3553 2473 3567 2487
rect 3493 2432 3507 2446
rect 3533 2432 3547 2446
rect 3513 2413 3527 2427
rect 3433 2353 3447 2367
rect 3473 2353 3487 2367
rect 3233 2273 3247 2287
rect 3433 2273 3447 2287
rect 3193 2254 3207 2268
rect 3233 2254 3247 2268
rect 3273 2254 3287 2268
rect 3373 2253 3387 2267
rect 3733 2933 3747 2947
rect 3693 2793 3707 2807
rect 3753 2913 3767 2927
rect 3813 2873 3827 2887
rect 3793 2833 3807 2847
rect 3773 2793 3787 2807
rect 3733 2774 3747 2788
rect 3993 3273 4007 3287
rect 4033 3133 4047 3147
rect 4013 3093 4027 3107
rect 4013 3053 4027 3067
rect 3873 3013 3887 3027
rect 3933 2994 3947 3008
rect 3993 2993 4007 3007
rect 3873 2952 3887 2966
rect 3913 2952 3927 2966
rect 3953 2952 3967 2966
rect 3993 2952 4007 2966
rect 3853 2853 3867 2867
rect 3813 2813 3827 2827
rect 3833 2774 3847 2788
rect 3813 2733 3827 2747
rect 3793 2713 3807 2727
rect 3773 2673 3787 2687
rect 3853 2713 3867 2727
rect 3713 2593 3727 2607
rect 3653 2573 3667 2587
rect 3773 2573 3787 2587
rect 3653 2493 3667 2507
rect 3673 2393 3687 2407
rect 3633 2313 3647 2327
rect 3753 2473 3767 2487
rect 3753 2393 3767 2407
rect 3813 2613 3827 2627
rect 3833 2593 3847 2607
rect 3933 2853 3947 2867
rect 4013 2853 4027 2867
rect 3913 2773 3927 2787
rect 3913 2653 3927 2667
rect 3813 2573 3827 2587
rect 3893 2573 3907 2587
rect 3833 2553 3847 2567
rect 3913 2513 3927 2527
rect 3833 2493 3847 2507
rect 3873 2474 3887 2488
rect 3793 2432 3807 2446
rect 3833 2413 3847 2427
rect 3773 2353 3787 2367
rect 3753 2313 3767 2327
rect 3693 2293 3707 2307
rect 3733 2293 3747 2307
rect 3513 2273 3527 2287
rect 3593 2273 3607 2287
rect 3173 2212 3187 2226
rect 3293 2212 3307 2226
rect 3253 2173 3267 2187
rect 3153 2093 3167 2107
rect 3013 1974 3027 1988
rect 3073 1974 3087 1988
rect 2893 1933 2907 1947
rect 3053 1932 3067 1946
rect 2973 1873 2987 1887
rect 2813 1833 2827 1847
rect 2973 1813 2987 1827
rect 2733 1773 2747 1787
rect 2973 1753 2987 1767
rect 2693 1733 2707 1747
rect 2733 1733 2747 1747
rect 2633 1714 2647 1728
rect 2673 1714 2687 1728
rect 3173 1934 3187 1948
rect 3373 2212 3387 2226
rect 3453 2212 3467 2226
rect 3793 2254 3807 2268
rect 3693 2193 3707 2207
rect 3413 2173 3427 2187
rect 3613 2173 3627 2187
rect 3773 2193 3787 2207
rect 3733 2113 3747 2127
rect 3433 2093 3447 2107
rect 3373 2053 3387 2067
rect 3373 1873 3387 1887
rect 3533 2073 3547 2087
rect 3473 1974 3487 1988
rect 3453 1934 3467 1948
rect 3633 1993 3647 2007
rect 3773 1973 3787 1987
rect 3433 1893 3447 1907
rect 3453 1873 3467 1887
rect 3793 1893 3807 1907
rect 3453 1852 3467 1866
rect 3773 1853 3787 1867
rect 3353 1833 3367 1847
rect 3433 1833 3447 1847
rect 3313 1813 3327 1827
rect 3393 1813 3407 1827
rect 2733 1673 2747 1687
rect 2673 1613 2687 1627
rect 2873 1573 2887 1587
rect 2933 1573 2947 1587
rect 2753 1533 2767 1547
rect 3073 1713 3087 1727
rect 3033 1672 3047 1686
rect 3093 1672 3107 1686
rect 3253 1712 3267 1726
rect 3253 1672 3267 1686
rect 3233 1593 3247 1607
rect 2933 1473 2947 1487
rect 2853 1454 2867 1468
rect 2913 1454 2927 1468
rect 2973 1532 2987 1546
rect 3073 1533 3087 1547
rect 3193 1533 3207 1547
rect 2873 1412 2887 1426
rect 2953 1413 2967 1427
rect 3153 1473 3167 1487
rect 3113 1434 3127 1448
rect 3253 1513 3267 1527
rect 3233 1473 3247 1487
rect 3193 1453 3207 1467
rect 3253 1453 3267 1467
rect 3173 1434 3187 1448
rect 3293 1434 3307 1448
rect 3333 1434 3347 1448
rect 2973 1393 2987 1407
rect 2873 1353 2887 1367
rect 2633 1313 2647 1327
rect 2853 1313 2867 1327
rect 2573 1133 2587 1147
rect 2533 1113 2547 1127
rect 2453 1093 2467 1107
rect 2513 1093 2527 1107
rect 2413 1013 2427 1027
rect 2453 953 2467 967
rect 2393 833 2407 847
rect 2093 653 2107 667
rect 2033 533 2047 547
rect 1833 493 1847 507
rect 1512 352 1526 366
rect 1533 353 1547 367
rect 1893 394 1907 408
rect 1573 352 1587 366
rect 1673 352 1687 366
rect 1753 352 1767 366
rect 1833 352 1847 366
rect 1873 352 1887 366
rect 1653 313 1667 327
rect 1713 313 1727 327
rect 1493 293 1507 307
rect 1553 174 1567 188
rect 1953 293 1967 307
rect 1913 253 1927 267
rect 1993 253 2007 267
rect 1713 173 1727 187
rect 1893 152 1907 166
rect 1993 152 2007 166
rect 2032 433 2046 447
rect 2053 433 2067 447
rect 2393 632 2407 646
rect 2273 533 2287 547
rect 2373 533 2387 547
rect 2133 433 2147 447
rect 2093 394 2107 408
rect 2033 352 2047 366
rect 2073 352 2087 366
rect 2153 352 2167 366
rect 2313 394 2327 408
rect 2133 152 2147 166
rect 2333 352 2347 366
rect 2333 273 2347 287
rect 2293 253 2307 267
rect 2473 913 2487 927
rect 2553 1093 2567 1107
rect 2553 973 2567 987
rect 2573 953 2587 967
rect 2533 914 2547 928
rect 2573 872 2587 886
rect 2673 1214 2687 1228
rect 2733 1213 2747 1227
rect 2773 1214 2787 1228
rect 2833 1214 2847 1228
rect 2893 1313 2907 1327
rect 2953 1313 2967 1327
rect 3033 1313 3047 1327
rect 2933 1214 2947 1228
rect 2693 1153 2707 1167
rect 2773 1153 2787 1167
rect 2893 1133 2907 1147
rect 2853 1093 2867 1107
rect 2893 1093 2907 1107
rect 2933 1033 2947 1047
rect 2653 953 2667 967
rect 2713 914 2727 928
rect 2813 913 2827 927
rect 2853 914 2867 928
rect 2653 872 2667 886
rect 2513 813 2527 827
rect 2573 733 2587 747
rect 2493 694 2507 708
rect 2533 694 2547 708
rect 2613 694 2627 708
rect 2473 632 2487 646
rect 2453 553 2467 567
rect 2733 872 2747 886
rect 2792 872 2806 886
rect 2813 872 2827 886
rect 2873 872 2887 886
rect 2693 813 2707 827
rect 2713 793 2727 807
rect 2733 773 2747 787
rect 2713 694 2727 708
rect 2553 652 2567 666
rect 2653 652 2667 666
rect 2613 633 2627 647
rect 2513 553 2527 567
rect 2593 553 2607 567
rect 2493 513 2507 527
rect 2473 473 2487 487
rect 2433 394 2447 408
rect 2453 333 2467 347
rect 2273 152 2287 166
rect 1433 132 1447 146
rect 1553 133 1567 147
rect 1373 73 1387 87
rect 2433 233 2447 247
rect 2573 513 2587 527
rect 2533 493 2547 507
rect 2533 394 2547 408
rect 2593 433 2607 447
rect 2753 513 2767 527
rect 2653 473 2667 487
rect 2993 1253 3007 1267
rect 2993 1214 3007 1228
rect 3093 1392 3107 1406
rect 3153 1393 3167 1407
rect 3173 1333 3187 1347
rect 3273 1392 3287 1406
rect 3233 1313 3247 1327
rect 3373 1473 3387 1487
rect 3353 1413 3367 1427
rect 3333 1293 3347 1307
rect 3053 1253 3067 1267
rect 3653 1793 3667 1807
rect 3553 1753 3567 1767
rect 3453 1712 3467 1726
rect 3413 1633 3427 1647
rect 3513 1693 3527 1707
rect 3453 1613 3467 1627
rect 3433 1533 3447 1547
rect 3473 1533 3487 1547
rect 3453 1513 3467 1527
rect 3413 1453 3427 1467
rect 3453 1454 3467 1468
rect 3493 1454 3507 1468
rect 3533 1412 3547 1426
rect 3393 1373 3407 1387
rect 3513 1313 3527 1327
rect 3813 1833 3827 1847
rect 3853 2313 3867 2327
rect 3893 2313 3907 2327
rect 3893 2273 3907 2287
rect 4053 3093 4067 3107
rect 4273 3513 4287 3527
rect 4473 3772 4487 3786
rect 4513 3772 4527 3786
rect 4553 3772 4567 3786
rect 4453 3753 4467 3767
rect 4433 3693 4447 3707
rect 4513 3733 4527 3747
rect 4453 3673 4467 3687
rect 4453 3652 4467 3666
rect 4433 3633 4447 3647
rect 4413 3613 4427 3627
rect 4513 3613 4527 3627
rect 4373 3553 4387 3567
rect 4413 3592 4427 3606
rect 4393 3533 4407 3547
rect 4473 3573 4487 3587
rect 4273 3433 4287 3447
rect 4253 3393 4267 3407
rect 4213 3333 4227 3347
rect 4113 3313 4127 3327
rect 4073 3073 4087 3087
rect 4073 3033 4087 3047
rect 4093 3013 4107 3027
rect 4293 3413 4307 3427
rect 4393 3453 4407 3467
rect 4533 3553 4547 3567
rect 4493 3533 4507 3547
rect 4473 3453 4487 3467
rect 4353 3433 4367 3447
rect 4453 3433 4467 3447
rect 4693 4093 4707 4107
rect 4653 4073 4667 4087
rect 4753 4232 4767 4246
rect 4733 4153 4747 4167
rect 4853 4733 4867 4747
rect 4893 5093 4907 5107
rect 4873 4613 4887 4627
rect 4973 5374 4987 5388
rect 4973 5333 4987 5347
rect 4953 5273 4967 5287
rect 5053 5653 5067 5667
rect 5273 6114 5287 6128
rect 5453 6213 5467 6227
rect 5333 6173 5347 6187
rect 5393 6173 5407 6187
rect 5253 6072 5267 6086
rect 5313 6073 5327 6087
rect 5353 6114 5367 6128
rect 5513 6233 5527 6247
rect 5633 6414 5647 6428
rect 5733 6413 5747 6427
rect 5793 6414 5807 6428
rect 5893 6413 5907 6427
rect 5953 6414 5967 6428
rect 6053 6413 6067 6427
rect 6133 6414 6147 6428
rect 6212 6413 6226 6427
rect 6233 6414 6247 6428
rect 6293 6414 6307 6428
rect 6473 6433 6487 6447
rect 6533 6433 6547 6447
rect 6873 6433 6887 6447
rect 5613 6372 5627 6386
rect 5653 6372 5667 6386
rect 5693 6273 5707 6287
rect 5733 6233 5747 6247
rect 5693 6213 5707 6227
rect 5893 6372 5907 6386
rect 5933 6372 5947 6386
rect 6033 6353 6047 6367
rect 5973 6333 5987 6347
rect 5873 6313 5887 6327
rect 5793 6293 5807 6307
rect 5333 6053 5347 6067
rect 5293 5953 5307 5967
rect 5193 5933 5207 5947
rect 5253 5933 5267 5947
rect 5213 5894 5227 5908
rect 5153 5813 5167 5827
rect 5233 5852 5247 5866
rect 5313 5913 5327 5927
rect 5253 5813 5267 5827
rect 5133 5773 5147 5787
rect 5193 5773 5207 5787
rect 5113 5733 5127 5747
rect 5073 5633 5087 5647
rect 5153 5633 5167 5647
rect 5113 5594 5127 5608
rect 5193 5594 5207 5608
rect 5073 5573 5087 5587
rect 5053 5433 5067 5447
rect 5133 5552 5147 5566
rect 5173 5552 5187 5566
rect 5133 5513 5147 5527
rect 5113 5493 5127 5507
rect 5073 5413 5087 5427
rect 5033 5393 5047 5407
rect 5073 5374 5087 5388
rect 5513 6113 5527 6127
rect 5573 6114 5587 6128
rect 5493 6053 5507 6067
rect 5373 6033 5387 6047
rect 5433 6033 5447 6047
rect 5353 5893 5367 5907
rect 5393 5894 5407 5908
rect 5333 5853 5347 5867
rect 5373 5813 5387 5827
rect 5333 5793 5347 5807
rect 5413 5793 5427 5807
rect 5292 5773 5293 5787
rect 5293 5773 5306 5787
rect 5313 5773 5327 5787
rect 5333 5753 5347 5767
rect 5293 5693 5307 5707
rect 5273 5573 5287 5587
rect 5573 5993 5587 6007
rect 5633 6072 5647 6086
rect 5613 6013 5627 6027
rect 5593 5953 5607 5967
rect 5573 5914 5587 5928
rect 5573 5893 5587 5907
rect 5653 5953 5667 5967
rect 5773 6193 5787 6207
rect 5713 6173 5727 6187
rect 5853 6193 5867 6207
rect 5793 6114 5807 6128
rect 5713 6072 5727 6086
rect 5773 6072 5787 6086
rect 5693 6033 5707 6047
rect 5813 6033 5827 6047
rect 5853 6013 5867 6027
rect 5893 6233 5907 6247
rect 5933 6153 5947 6167
rect 6033 6153 6047 6167
rect 6213 6372 6227 6386
rect 6153 6353 6167 6367
rect 6273 6372 6287 6386
rect 6233 6293 6247 6307
rect 6373 6353 6387 6367
rect 6313 6253 6327 6267
rect 6113 6233 6127 6247
rect 6353 6133 6367 6147
rect 5973 6114 5987 6128
rect 6033 6114 6047 6128
rect 6073 6114 6087 6128
rect 6153 6114 6167 6128
rect 6233 6114 6247 6128
rect 6273 6114 6287 6128
rect 6313 6114 6327 6128
rect 5893 6072 5907 6086
rect 5953 6072 5967 6086
rect 5953 5993 5967 6007
rect 5733 5973 5747 5987
rect 5873 5973 5887 5987
rect 5513 5833 5527 5847
rect 5493 5673 5507 5687
rect 5593 5813 5607 5827
rect 5553 5793 5567 5807
rect 5633 5753 5647 5767
rect 5593 5693 5607 5707
rect 5513 5653 5527 5667
rect 5553 5653 5567 5667
rect 5613 5653 5627 5667
rect 5373 5633 5387 5647
rect 5473 5613 5487 5627
rect 5513 5613 5527 5627
rect 5333 5594 5347 5608
rect 5373 5594 5387 5608
rect 5433 5594 5447 5608
rect 5213 5533 5227 5547
rect 5252 5533 5266 5547
rect 5273 5533 5287 5547
rect 5173 5513 5187 5527
rect 5213 5473 5227 5487
rect 5153 5433 5167 5447
rect 5133 5353 5147 5367
rect 5053 5332 5067 5346
rect 4993 5253 5007 5267
rect 5053 5253 5067 5267
rect 4993 5153 5007 5167
rect 4933 5093 4947 5107
rect 4913 5073 4927 5087
rect 4953 5074 4967 5088
rect 5113 5273 5127 5287
rect 5093 5133 5107 5147
rect 5053 5113 5067 5127
rect 5013 5073 5027 5087
rect 4933 5032 4947 5046
rect 4913 4953 4927 4967
rect 4933 4933 4947 4947
rect 4973 4913 4987 4927
rect 4953 4873 4967 4887
rect 5033 5053 5047 5067
rect 5033 4993 5047 5007
rect 5133 5233 5147 5247
rect 5173 5374 5187 5388
rect 5293 5513 5307 5527
rect 5273 5413 5287 5427
rect 5253 5374 5267 5388
rect 5233 5332 5247 5346
rect 5393 5552 5407 5566
rect 5353 5513 5367 5527
rect 5333 5493 5347 5507
rect 5553 5594 5567 5608
rect 5533 5552 5547 5566
rect 5513 5533 5527 5547
rect 5473 5493 5487 5507
rect 5453 5473 5467 5487
rect 5353 5453 5367 5467
rect 5433 5453 5447 5467
rect 5333 5433 5347 5447
rect 5473 5453 5487 5467
rect 5453 5433 5467 5447
rect 5533 5453 5547 5467
rect 5173 5293 5187 5307
rect 5273 5313 5287 5327
rect 5253 5293 5267 5307
rect 5233 5253 5247 5267
rect 5153 5213 5167 5227
rect 5193 5213 5207 5227
rect 5133 5093 5147 5107
rect 4933 4853 4947 4867
rect 5053 4893 5067 4907
rect 5053 4853 5067 4867
rect 4912 4812 4926 4826
rect 4933 4812 4947 4826
rect 4973 4812 4987 4826
rect 5093 5032 5107 5046
rect 5153 5033 5167 5047
rect 5113 4913 5127 4927
rect 5093 4873 5107 4887
rect 4933 4753 4947 4767
rect 4973 4753 4987 4767
rect 4913 4733 4927 4747
rect 4933 4713 4947 4727
rect 4913 4673 4927 4687
rect 4953 4673 4967 4687
rect 4933 4573 4947 4587
rect 4773 4213 4787 4227
rect 4753 4113 4767 4127
rect 4593 3992 4607 4006
rect 4633 3992 4647 4006
rect 4593 3873 4607 3887
rect 4633 3833 4647 3847
rect 4713 3973 4727 3987
rect 4753 3913 4767 3927
rect 4613 3813 4627 3827
rect 4653 3814 4667 3828
rect 4753 3833 4767 3847
rect 4733 3813 4747 3827
rect 4633 3772 4647 3786
rect 4673 3772 4687 3786
rect 4593 3733 4607 3747
rect 4633 3733 4647 3747
rect 4573 3693 4587 3707
rect 4753 3753 4767 3767
rect 4733 3713 4747 3727
rect 4673 3693 4687 3707
rect 4653 3613 4667 3627
rect 4553 3533 4567 3547
rect 4633 3493 4647 3507
rect 4593 3433 4607 3447
rect 4553 3413 4567 3427
rect 4653 3473 4667 3487
rect 4713 3673 4727 3687
rect 4693 3653 4707 3667
rect 4693 3613 4707 3627
rect 4733 3653 4747 3667
rect 4733 3613 4747 3627
rect 4713 3593 4727 3607
rect 4873 4512 4887 4526
rect 4893 4493 4907 4507
rect 4812 4433 4826 4447
rect 4833 4433 4847 4447
rect 4893 4433 4907 4447
rect 4833 4393 4847 4407
rect 4893 4393 4907 4407
rect 4813 4373 4827 4387
rect 4853 4353 4867 4367
rect 4813 4333 4827 4347
rect 5073 4653 5087 4667
rect 5053 4633 5067 4647
rect 4973 4593 4987 4607
rect 5013 4554 5027 4568
rect 5073 4553 5087 4567
rect 4953 4533 4967 4547
rect 4933 4473 4947 4487
rect 4932 4452 4946 4466
rect 4953 4453 4967 4467
rect 5033 4453 5047 4467
rect 4953 4413 4967 4427
rect 4933 4393 4947 4407
rect 4913 4373 4927 4387
rect 4913 4352 4927 4366
rect 4993 4413 5007 4427
rect 5073 4413 5087 4427
rect 4973 4353 4987 4367
rect 4953 4333 4967 4347
rect 4833 4292 4847 4306
rect 4793 4173 4807 4187
rect 4853 4173 4867 4187
rect 4813 4133 4827 4147
rect 4913 4093 4927 4107
rect 4833 4053 4847 4067
rect 4873 4034 4887 4048
rect 4953 4033 4967 4047
rect 4813 3993 4827 4006
rect 4813 3992 4827 3993
rect 4853 3992 4867 4006
rect 4793 3973 4807 3987
rect 4893 3973 4907 3987
rect 4792 3933 4806 3947
rect 4813 3933 4827 3947
rect 4893 3952 4907 3966
rect 4853 3873 4867 3887
rect 4793 3833 4807 3847
rect 4833 3814 4847 3828
rect 4813 3772 4827 3786
rect 4873 3772 4887 3786
rect 4833 3753 4847 3767
rect 4773 3573 4787 3587
rect 4693 3513 4707 3527
rect 4733 3514 4747 3528
rect 4793 3553 4807 3567
rect 4793 3532 4807 3546
rect 4813 3513 4827 3527
rect 4653 3452 4667 3466
rect 4353 3373 4367 3387
rect 4473 3373 4487 3387
rect 4513 3373 4527 3387
rect 4633 3373 4647 3387
rect 4293 3293 4307 3307
rect 4133 3193 4147 3207
rect 4173 3153 4187 3167
rect 4073 2893 4087 2907
rect 4053 2773 4067 2787
rect 3973 2673 3987 2687
rect 4013 2593 4027 2607
rect 3953 2573 3967 2587
rect 4013 2493 4027 2507
rect 4133 2952 4147 2966
rect 4093 2873 4107 2887
rect 4313 3233 4327 3247
rect 4293 3093 4307 3107
rect 4213 3033 4227 3047
rect 4333 3213 4347 3227
rect 4273 2994 4287 3008
rect 4313 2992 4327 3006
rect 4253 2952 4267 2966
rect 4313 2952 4327 2966
rect 4433 3273 4447 3287
rect 4433 3213 4447 3227
rect 4353 3153 4367 3167
rect 4593 3233 4607 3247
rect 4473 3173 4487 3187
rect 4453 3133 4467 3147
rect 4573 3133 4587 3147
rect 4553 3113 4567 3127
rect 4473 3073 4487 3087
rect 4353 2994 4367 3008
rect 4433 2994 4447 3008
rect 4713 3472 4727 3486
rect 4753 3433 4767 3447
rect 4733 3413 4747 3427
rect 4613 3013 4627 3027
rect 4653 3013 4667 3027
rect 4413 2952 4427 2966
rect 4353 2913 4367 2927
rect 4433 2913 4447 2927
rect 4333 2893 4347 2907
rect 4213 2873 4227 2887
rect 4273 2853 4287 2867
rect 4173 2813 4187 2827
rect 4173 2774 4187 2788
rect 4253 2753 4267 2767
rect 4193 2732 4207 2746
rect 4253 2653 4267 2667
rect 4153 2553 4167 2567
rect 4113 2493 4127 2507
rect 4173 2474 4187 2488
rect 3993 2432 4007 2446
rect 4033 2432 4047 2446
rect 4073 2432 4087 2446
rect 4113 2432 4127 2446
rect 4153 2432 4167 2446
rect 4193 2432 4207 2446
rect 3953 2413 3967 2427
rect 3993 2393 4007 2407
rect 3933 2293 3947 2307
rect 4013 2293 4027 2307
rect 3873 2253 3887 2267
rect 3973 2254 3987 2268
rect 4453 2873 4467 2887
rect 4433 2833 4447 2847
rect 4353 2793 4367 2807
rect 4293 2773 4307 2787
rect 4333 2732 4347 2746
rect 4493 2793 4507 2807
rect 4533 2793 4547 2807
rect 4573 2793 4587 2807
rect 4293 2673 4307 2687
rect 4373 2653 4387 2667
rect 4293 2593 4307 2607
rect 4313 2474 4327 2488
rect 4413 2573 4427 2587
rect 4413 2513 4427 2527
rect 4433 2493 4447 2507
rect 4273 2413 4287 2427
rect 4053 2393 4067 2407
rect 4033 2254 4047 2268
rect 4013 2233 4027 2247
rect 3873 2212 3887 2226
rect 3913 2212 3927 2226
rect 3853 2193 3867 2207
rect 3973 2133 3987 2147
rect 3953 2113 3967 2127
rect 3913 2073 3927 2087
rect 3893 2033 3907 2047
rect 3873 1932 3887 1946
rect 3853 1833 3867 1847
rect 3633 1692 3647 1706
rect 3673 1692 3687 1706
rect 3713 1692 3727 1706
rect 3673 1633 3687 1647
rect 3813 1553 3827 1567
rect 3793 1513 3807 1527
rect 3653 1414 3667 1428
rect 3513 1273 3527 1287
rect 3553 1273 3567 1287
rect 3733 1273 3747 1287
rect 3373 1213 3387 1227
rect 3413 1213 3427 1227
rect 3013 1172 3027 1186
rect 2973 1113 2987 1127
rect 3073 1113 3087 1127
rect 2953 993 2967 1007
rect 3013 973 3027 987
rect 3093 913 3107 927
rect 3153 914 3167 928
rect 3193 914 3207 928
rect 2973 873 2987 887
rect 3033 872 3047 886
rect 2993 853 3007 867
rect 3033 853 3047 867
rect 3073 853 3087 867
rect 2873 733 2887 747
rect 2933 733 2947 747
rect 2833 694 2847 708
rect 2913 694 2927 708
rect 3053 733 3067 747
rect 3133 853 3147 867
rect 3193 773 3207 787
rect 3073 713 3087 727
rect 3113 713 3127 727
rect 2893 652 2907 666
rect 2993 653 3007 667
rect 3293 973 3307 987
rect 3433 1173 3447 1187
rect 3433 1093 3447 1107
rect 3453 1033 3467 1047
rect 3433 993 3447 1007
rect 3373 953 3387 967
rect 3413 914 3427 928
rect 3373 853 3387 867
rect 3273 833 3287 847
rect 3473 872 3487 886
rect 3453 853 3467 867
rect 3433 813 3447 827
rect 3393 793 3407 807
rect 3433 733 3447 747
rect 2833 633 2847 647
rect 2833 573 2847 587
rect 2933 493 2947 507
rect 2833 433 2847 447
rect 2793 413 2807 427
rect 2613 394 2627 408
rect 2673 394 2687 408
rect 2593 352 2607 366
rect 2533 333 2547 347
rect 2653 313 2667 327
rect 2613 233 2627 247
rect 2453 193 2467 207
rect 2513 193 2527 207
rect 2473 154 2487 168
rect 2513 154 2527 168
rect 2053 112 2067 126
rect 2113 112 2127 126
rect 2413 112 2427 126
rect 2773 394 2787 408
rect 2693 353 2707 367
rect 2753 352 2767 366
rect 2813 313 2827 327
rect 2693 273 2707 287
rect 2673 253 2687 267
rect 2693 233 2707 247
rect 2693 174 2707 188
rect 2793 173 2807 187
rect 2613 132 2627 146
rect 2673 132 2687 146
rect 2713 132 2727 146
rect 2853 413 2867 427
rect 2833 293 2847 307
rect 2893 394 2907 408
rect 3073 652 3087 666
rect 3113 652 3127 666
rect 3073 493 3087 507
rect 3253 613 3267 627
rect 3253 553 3267 567
rect 3273 493 3287 507
rect 3213 473 3227 487
rect 2953 352 2967 366
rect 3033 353 3047 367
rect 2913 313 2927 327
rect 2893 253 2907 267
rect 2853 213 2867 227
rect 2953 213 2967 227
rect 3053 313 3067 327
rect 3133 313 3147 327
rect 3153 253 3167 267
rect 3193 253 3207 267
rect 3373 473 3387 487
rect 3293 433 3307 447
rect 3333 352 3347 366
rect 3373 313 3387 327
rect 3453 593 3467 607
rect 3633 1172 3647 1186
rect 3873 1553 3887 1567
rect 3913 1993 3927 2007
rect 3913 1873 3927 1887
rect 4113 2313 4127 2327
rect 4153 2254 4167 2268
rect 4053 2212 4067 2226
rect 4133 2212 4147 2226
rect 4093 2193 4107 2207
rect 4393 2432 4407 2446
rect 4413 2413 4427 2427
rect 4353 2393 4367 2407
rect 4393 2393 4407 2407
rect 4213 2353 4227 2367
rect 4333 2353 4347 2367
rect 4233 2313 4247 2327
rect 4253 2293 4267 2307
rect 4233 2212 4247 2226
rect 4213 2173 4227 2187
rect 4133 2153 4147 2167
rect 4193 2153 4207 2167
rect 4093 2113 4107 2127
rect 4013 2053 4027 2067
rect 4053 2053 4067 2067
rect 4053 1973 4067 1987
rect 4073 1954 4087 1968
rect 3973 1912 3987 1926
rect 4013 1912 4027 1926
rect 4053 1912 4067 1926
rect 3953 1813 3967 1827
rect 4033 1813 4047 1827
rect 3933 1734 3947 1748
rect 3993 1733 4007 1747
rect 3953 1653 3967 1667
rect 3993 1613 4007 1627
rect 3993 1553 4007 1567
rect 3893 1513 3907 1527
rect 3913 1493 3927 1507
rect 3933 1433 3947 1447
rect 3833 1373 3847 1387
rect 3793 1213 3807 1227
rect 3793 1093 3807 1107
rect 3593 1073 3607 1087
rect 3553 914 3567 928
rect 3693 993 3707 1007
rect 3673 914 3687 928
rect 3533 872 3547 886
rect 3573 813 3587 827
rect 3593 733 3607 747
rect 3633 713 3647 727
rect 3613 652 3627 666
rect 3813 872 3827 886
rect 3893 1333 3907 1347
rect 3853 1253 3867 1267
rect 4193 2093 4207 2107
rect 4193 2033 4207 2047
rect 4393 2233 4407 2247
rect 4273 2212 4287 2226
rect 4313 2193 4327 2207
rect 4293 2133 4307 2147
rect 4253 1973 4267 1987
rect 4153 1954 4167 1968
rect 4193 1954 4207 1968
rect 4233 1954 4247 1968
rect 4153 1913 4167 1927
rect 4253 1912 4267 1926
rect 4213 1873 4227 1887
rect 4313 2053 4327 2067
rect 4313 1973 4327 1987
rect 4333 1954 4347 1968
rect 4413 2013 4427 2027
rect 4513 2732 4527 2746
rect 4553 2653 4567 2667
rect 4553 2593 4567 2607
rect 4513 2513 4527 2527
rect 4553 2513 4567 2527
rect 4653 2952 4667 2966
rect 4813 3393 4827 3407
rect 4793 3373 4807 3387
rect 4773 3353 4787 3367
rect 4753 3053 4767 3067
rect 4793 3133 4807 3147
rect 4853 3653 4867 3667
rect 4913 3814 4927 3828
rect 5013 4373 5027 4387
rect 5033 4353 5047 4367
rect 5033 4334 5047 4348
rect 5153 4854 5167 4868
rect 5353 5374 5367 5388
rect 5413 5374 5427 5388
rect 5513 5413 5527 5427
rect 5493 5373 5507 5387
rect 5353 5313 5367 5327
rect 5433 5332 5447 5346
rect 5293 5273 5307 5287
rect 5333 5272 5347 5286
rect 5313 5213 5327 5227
rect 5313 5173 5327 5187
rect 5213 5033 5227 5047
rect 5213 4993 5227 5007
rect 5273 5032 5287 5046
rect 5313 5032 5327 5046
rect 5373 5253 5387 5267
rect 5373 5213 5387 5227
rect 5473 5213 5487 5227
rect 5373 5173 5387 5187
rect 5433 5113 5447 5127
rect 5373 5093 5387 5107
rect 5393 5074 5407 5088
rect 5493 5193 5507 5207
rect 5393 5013 5407 5027
rect 5333 4973 5347 4987
rect 5233 4953 5247 4967
rect 5233 4854 5247 4868
rect 5173 4812 5187 4826
rect 5173 4793 5187 4807
rect 5213 4773 5227 4787
rect 5233 4753 5247 4767
rect 5133 4733 5147 4747
rect 5173 4733 5187 4747
rect 5213 4733 5227 4747
rect 5273 4913 5287 4927
rect 5293 4853 5307 4867
rect 5373 4812 5387 4826
rect 5273 4793 5287 4807
rect 5353 4793 5367 4807
rect 5273 4733 5287 4747
rect 5353 4772 5367 4786
rect 5353 4733 5367 4747
rect 5333 4693 5347 4707
rect 5293 4673 5307 4687
rect 5133 4653 5147 4667
rect 5253 4653 5267 4667
rect 5113 4513 5127 4527
rect 5093 4373 5107 4387
rect 5213 4633 5227 4647
rect 5173 4554 5187 4568
rect 5473 5033 5487 5047
rect 5613 5553 5627 5567
rect 5633 5513 5647 5527
rect 5853 5894 5867 5908
rect 5913 5894 5927 5908
rect 5713 5813 5727 5827
rect 6033 6033 6047 6047
rect 6053 5953 6067 5967
rect 6053 5913 6067 5927
rect 6173 6072 6187 6086
rect 6153 6013 6167 6027
rect 6133 5993 6147 6007
rect 5993 5873 6007 5887
rect 5973 5833 5987 5847
rect 5873 5813 5887 5827
rect 5753 5773 5767 5787
rect 5853 5773 5867 5787
rect 5773 5733 5787 5747
rect 5713 5594 5727 5608
rect 5793 5693 5807 5707
rect 5913 5773 5927 5787
rect 5873 5653 5887 5667
rect 5813 5593 5827 5607
rect 5873 5594 5887 5608
rect 5953 5673 5967 5687
rect 6073 5894 6087 5908
rect 6113 5894 6127 5908
rect 6013 5833 6027 5847
rect 6133 5853 6147 5867
rect 6093 5833 6107 5847
rect 5993 5813 6007 5827
rect 6133 5753 6147 5767
rect 6093 5713 6107 5727
rect 6193 5973 6207 5987
rect 6173 5893 6187 5907
rect 6153 5693 6167 5707
rect 5693 5533 5707 5547
rect 5673 5493 5687 5507
rect 5653 5473 5667 5487
rect 5633 5453 5647 5467
rect 5633 5432 5647 5446
rect 5573 5413 5587 5427
rect 5673 5453 5687 5467
rect 5653 5373 5667 5387
rect 5533 5293 5547 5307
rect 5673 5313 5687 5327
rect 5653 5293 5667 5307
rect 5673 5253 5687 5267
rect 5653 5233 5667 5247
rect 5613 5213 5627 5227
rect 5653 5173 5667 5187
rect 5613 5133 5627 5147
rect 5513 5074 5527 5088
rect 5573 5074 5587 5088
rect 5613 5074 5627 5088
rect 5553 5032 5567 5046
rect 5593 5032 5607 5046
rect 5633 5033 5647 5047
rect 5493 4973 5507 4987
rect 5533 4953 5547 4967
rect 5613 4953 5627 4967
rect 5533 4913 5547 4927
rect 5413 4854 5427 4868
rect 5493 4854 5507 4868
rect 5533 4854 5547 4868
rect 5593 4853 5607 4867
rect 5433 4793 5447 4807
rect 5413 4753 5427 4767
rect 5373 4653 5387 4667
rect 5373 4632 5387 4646
rect 5353 4593 5367 4607
rect 5233 4573 5247 4587
rect 5333 4573 5347 4587
rect 5253 4554 5267 4568
rect 5433 4673 5447 4687
rect 5433 4633 5447 4647
rect 5193 4512 5207 4526
rect 5293 4513 5307 4527
rect 5273 4493 5287 4507
rect 5293 4473 5307 4487
rect 5413 4553 5427 4567
rect 5413 4513 5427 4527
rect 5313 4413 5327 4427
rect 5173 4393 5187 4407
rect 5273 4393 5287 4407
rect 5013 4293 5027 4307
rect 4993 4133 5007 4147
rect 5073 4253 5087 4267
rect 5133 4292 5147 4306
rect 5113 4233 5127 4247
rect 5053 4133 5067 4147
rect 5093 4133 5107 4147
rect 5013 4073 5027 4087
rect 4993 4033 5007 4047
rect 5133 4213 5147 4227
rect 5153 4193 5167 4207
rect 5113 4113 5127 4127
rect 5193 4353 5207 4367
rect 5293 4334 5307 4348
rect 5233 4292 5247 4306
rect 5193 4253 5207 4267
rect 5233 4233 5247 4247
rect 5193 4193 5207 4207
rect 5133 4073 5147 4087
rect 5113 4033 5127 4047
rect 5013 3992 5027 4006
rect 4993 3913 5007 3927
rect 5073 3992 5087 4006
rect 5073 3873 5087 3887
rect 5033 3853 5047 3867
rect 4933 3772 4947 3786
rect 4913 3733 4927 3747
rect 4993 3772 5007 3786
rect 5033 3733 5047 3747
rect 4953 3713 4967 3727
rect 5093 3772 5107 3786
rect 5073 3693 5087 3707
rect 5173 4113 5187 4127
rect 5153 3932 5167 3946
rect 5133 3913 5147 3927
rect 5313 4292 5327 4306
rect 5293 4273 5307 4287
rect 5273 4133 5287 4147
rect 5253 4073 5267 4087
rect 5213 4053 5227 4067
rect 5273 4053 5287 4067
rect 5253 3992 5267 4006
rect 5313 4253 5327 4267
rect 5313 4213 5327 4227
rect 5253 3913 5267 3927
rect 5173 3893 5187 3907
rect 5153 3833 5167 3847
rect 5173 3814 5187 3828
rect 5233 3813 5247 3827
rect 5153 3772 5167 3786
rect 5173 3753 5187 3767
rect 5153 3673 5167 3687
rect 5133 3593 5147 3607
rect 4893 3573 4907 3587
rect 5033 3573 5047 3587
rect 4872 3553 4886 3567
rect 4853 3514 4867 3528
rect 4893 3552 4907 3566
rect 4913 3514 4927 3528
rect 4893 3472 4907 3486
rect 5013 3472 5027 3486
rect 4873 3293 4887 3307
rect 4873 3252 4887 3266
rect 4853 3233 4867 3247
rect 4833 3113 4847 3127
rect 4813 3053 4827 3067
rect 4793 3033 4807 3047
rect 4773 3013 4787 3027
rect 4853 3013 4867 3027
rect 4813 2993 4827 3007
rect 4613 2833 4627 2847
rect 4673 2833 4687 2847
rect 4633 2773 4647 2787
rect 4693 2774 4707 2788
rect 4613 2732 4627 2746
rect 4673 2732 4687 2746
rect 4713 2733 4727 2747
rect 4673 2693 4687 2707
rect 4593 2593 4607 2607
rect 4552 2473 4566 2487
rect 4573 2473 4587 2487
rect 4573 2452 4587 2466
rect 4453 2433 4467 2447
rect 4493 2432 4507 2446
rect 4533 2413 4547 2427
rect 4573 2413 4587 2427
rect 4513 2333 4527 2347
rect 4493 2293 4507 2307
rect 4533 2313 4547 2327
rect 4513 2273 4527 2287
rect 4453 2254 4467 2268
rect 4493 2254 4507 2268
rect 4533 2254 4547 2268
rect 4473 2213 4487 2227
rect 4453 2133 4467 2147
rect 4433 1954 4447 1968
rect 4313 1912 4327 1926
rect 4293 1813 4307 1827
rect 4133 1793 4147 1807
rect 4153 1773 4167 1787
rect 4093 1734 4107 1748
rect 4073 1653 4087 1667
rect 4113 1573 4127 1587
rect 4033 1513 4047 1527
rect 4133 1473 4147 1487
rect 4053 1434 4067 1448
rect 3993 1392 4007 1406
rect 4033 1392 4047 1406
rect 4133 1313 4147 1327
rect 4073 1253 4087 1267
rect 3993 1214 4007 1228
rect 3913 1133 3927 1147
rect 3853 1033 3867 1047
rect 4013 1133 4027 1147
rect 3953 993 3967 1007
rect 3993 973 4007 987
rect 3953 914 3967 928
rect 3993 913 4007 927
rect 3853 872 3867 886
rect 3773 813 3787 827
rect 3853 773 3867 787
rect 3813 753 3827 767
rect 3693 713 3707 727
rect 3713 694 3727 708
rect 3773 694 3787 708
rect 3833 733 3847 747
rect 3693 652 3707 666
rect 3653 573 3667 587
rect 3833 693 3847 707
rect 3753 652 3767 666
rect 3553 553 3567 567
rect 3713 553 3727 567
rect 3493 513 3507 527
rect 3433 433 3447 447
rect 3273 193 3287 207
rect 3213 174 3227 188
rect 3633 533 3647 547
rect 3613 413 3627 427
rect 3513 352 3527 366
rect 3553 293 3567 307
rect 3453 233 3467 247
rect 3433 213 3447 227
rect 3513 193 3527 207
rect 3593 193 3607 207
rect 2953 132 2967 146
rect 3153 132 3167 146
rect 3193 132 3207 146
rect 3393 132 3407 146
rect 3533 132 3547 146
rect 3593 113 3607 127
rect 3073 93 3087 107
rect 3233 93 3247 107
rect 3353 93 3367 107
rect 3533 93 3547 107
rect 2473 73 2487 87
rect 2793 73 2807 87
rect 3793 473 3807 487
rect 3873 693 3887 707
rect 3953 833 3967 847
rect 3993 693 4007 707
rect 3893 652 3907 666
rect 3933 652 3947 666
rect 3893 593 3907 607
rect 4113 1214 4127 1228
rect 4093 1172 4107 1186
rect 4133 1053 4147 1067
rect 4093 1033 4107 1047
rect 4033 953 4047 967
rect 4193 1733 4207 1747
rect 4253 1734 4267 1748
rect 4293 1734 4307 1748
rect 4273 1692 4287 1706
rect 4413 1912 4427 1926
rect 4373 1813 4387 1827
rect 4513 2212 4527 2226
rect 4573 2213 4587 2227
rect 4533 2193 4547 2207
rect 4533 2153 4547 2167
rect 4533 2093 4547 2107
rect 4553 2033 4567 2047
rect 4513 1993 4527 2007
rect 4493 1953 4507 1967
rect 4373 1773 4387 1787
rect 4473 1773 4487 1787
rect 4413 1734 4427 1748
rect 4453 1734 4467 1748
rect 4773 2952 4787 2966
rect 4853 2933 4867 2947
rect 4833 2913 4847 2927
rect 4833 2873 4847 2887
rect 4773 2813 4787 2827
rect 4833 2813 4847 2827
rect 5133 3553 5147 3567
rect 5053 3533 5067 3547
rect 5033 3453 5047 3467
rect 4973 3393 4987 3407
rect 4933 3293 4947 3307
rect 4913 3013 4927 3027
rect 4892 2972 4906 2986
rect 4913 2973 4927 2987
rect 4873 2873 4887 2887
rect 4753 2773 4767 2787
rect 4753 2732 4767 2746
rect 4753 2653 4767 2667
rect 4733 2593 4747 2607
rect 4633 2553 4647 2567
rect 4693 2553 4707 2567
rect 4753 2474 4767 2488
rect 4653 2432 4667 2446
rect 4693 2393 4707 2407
rect 4653 2353 4667 2367
rect 4893 2774 4907 2788
rect 4793 2732 4807 2746
rect 5213 3773 5227 3787
rect 5213 3733 5227 3747
rect 5192 3713 5206 3727
rect 5213 3712 5227 3726
rect 5173 3613 5187 3627
rect 5153 3533 5167 3547
rect 5193 3514 5207 3528
rect 5233 3673 5247 3687
rect 5073 3493 5087 3507
rect 5053 3273 5067 3287
rect 5233 3513 5247 3527
rect 5253 3493 5267 3507
rect 5233 3453 5247 3467
rect 5233 3413 5247 3427
rect 5373 4473 5387 4487
rect 5353 4173 5367 4187
rect 5353 4133 5367 4147
rect 5353 4112 5367 4126
rect 5333 4034 5347 4048
rect 5333 3993 5347 4007
rect 5313 3933 5327 3947
rect 5333 3893 5347 3907
rect 5433 4493 5447 4507
rect 5513 4713 5527 4727
rect 5493 4633 5507 4647
rect 5473 4613 5487 4627
rect 5593 4613 5607 4627
rect 5513 4593 5527 4607
rect 5492 4553 5506 4567
rect 5513 4554 5527 4568
rect 5533 4512 5547 4526
rect 5513 4493 5527 4507
rect 5493 4472 5507 4486
rect 5473 4453 5487 4467
rect 5433 4433 5447 4447
rect 5433 4334 5447 4348
rect 5593 4512 5607 4526
rect 5513 4393 5527 4407
rect 5573 4393 5587 4407
rect 5393 4273 5407 4287
rect 5473 4273 5487 4287
rect 5453 4253 5467 4267
rect 5373 4093 5387 4107
rect 5433 4034 5447 4048
rect 5533 4333 5547 4347
rect 5513 4073 5527 4087
rect 5493 4033 5507 4047
rect 5473 4013 5487 4027
rect 5453 3993 5467 4007
rect 5413 3853 5427 3867
rect 5333 3633 5347 3647
rect 5293 3513 5307 3527
rect 5413 3772 5427 3786
rect 5393 3753 5407 3767
rect 5373 3513 5387 3527
rect 5633 4913 5647 4927
rect 5773 5553 5787 5567
rect 5733 5513 5747 5527
rect 5713 5493 5727 5507
rect 5793 5493 5807 5507
rect 5773 5473 5787 5487
rect 5753 5453 5767 5467
rect 5773 5393 5787 5407
rect 5713 5374 5727 5388
rect 5753 5374 5767 5388
rect 5813 5473 5827 5487
rect 5893 5552 5907 5566
rect 5873 5533 5887 5547
rect 5933 5533 5947 5547
rect 5853 5433 5867 5447
rect 5853 5393 5867 5407
rect 5733 5333 5747 5347
rect 5713 5293 5727 5307
rect 5713 5272 5727 5286
rect 5793 5313 5807 5327
rect 5733 5213 5747 5227
rect 5713 5193 5727 5207
rect 5693 5113 5707 5127
rect 5692 5074 5706 5088
rect 5673 4953 5687 4967
rect 5713 5073 5727 5087
rect 5753 5193 5767 5207
rect 5773 5113 5787 5127
rect 5753 5032 5767 5046
rect 5913 5513 5927 5527
rect 5933 5453 5947 5467
rect 5973 5653 5987 5667
rect 5973 5553 5987 5567
rect 5953 5433 5967 5447
rect 5913 5413 5927 5427
rect 5933 5374 5947 5388
rect 6093 5673 6107 5687
rect 6233 6073 6247 6087
rect 6333 6073 6347 6087
rect 6273 5933 6287 5947
rect 6333 5933 6347 5947
rect 6212 5893 6226 5907
rect 6233 5894 6247 5908
rect 6333 5893 6347 5907
rect 6193 5852 6207 5866
rect 6253 5852 6267 5866
rect 6293 5852 6307 5866
rect 6353 5833 6367 5847
rect 6193 5813 6207 5827
rect 6493 6173 6507 6187
rect 6393 6114 6407 6128
rect 6453 6114 6467 6128
rect 6473 6033 6487 6047
rect 6433 6013 6447 6027
rect 6433 5953 6447 5967
rect 6473 5894 6487 5908
rect 6513 5893 6527 5907
rect 6453 5852 6467 5866
rect 6333 5792 6347 5806
rect 6373 5793 6387 5807
rect 6413 5793 6427 5807
rect 6293 5773 6307 5787
rect 6193 5733 6207 5747
rect 6313 5693 6327 5707
rect 6133 5633 6147 5647
rect 6173 5633 6187 5647
rect 6053 5594 6067 5608
rect 6093 5594 6107 5608
rect 6033 5473 6047 5487
rect 6033 5433 6047 5447
rect 5913 5333 5927 5347
rect 5853 5293 5867 5307
rect 5813 5153 5827 5167
rect 5833 5133 5847 5147
rect 5813 5093 5827 5107
rect 5793 5013 5807 5027
rect 5833 5053 5847 5067
rect 5813 4993 5827 5007
rect 5773 4973 5787 4987
rect 5733 4953 5747 4967
rect 5693 4933 5707 4947
rect 5653 4893 5667 4907
rect 5693 4893 5707 4907
rect 5653 4854 5667 4868
rect 5673 4812 5687 4826
rect 5653 4793 5667 4807
rect 5653 4713 5667 4727
rect 5633 4693 5647 4707
rect 5653 4673 5667 4687
rect 5653 4633 5667 4647
rect 5713 4633 5727 4647
rect 5633 4573 5647 4587
rect 5653 4554 5667 4568
rect 5693 4554 5707 4568
rect 5673 4493 5687 4507
rect 5613 4353 5627 4367
rect 5573 4333 5587 4347
rect 5693 4393 5707 4407
rect 5613 4292 5627 4306
rect 5633 4253 5647 4267
rect 5633 4173 5647 4187
rect 5673 4193 5687 4207
rect 5653 4153 5667 4167
rect 5633 4133 5647 4147
rect 5573 4073 5587 4087
rect 5613 4073 5627 4087
rect 5553 4053 5567 4067
rect 5533 4033 5547 4047
rect 5573 4034 5587 4048
rect 5513 4013 5527 4027
rect 5573 3973 5587 3987
rect 5613 3973 5627 3987
rect 5533 3913 5547 3927
rect 5513 3893 5527 3907
rect 5553 3893 5567 3907
rect 5473 3853 5487 3867
rect 5453 3833 5467 3847
rect 5713 4352 5727 4366
rect 5693 4153 5707 4167
rect 5713 4113 5727 4127
rect 5753 4913 5767 4927
rect 5753 4833 5767 4847
rect 5873 5193 5887 5207
rect 5893 5153 5907 5167
rect 5953 5332 5967 5346
rect 5913 5113 5927 5127
rect 5893 5093 5907 5107
rect 6013 5293 6027 5307
rect 5992 5273 6006 5287
rect 5973 5193 5987 5207
rect 5953 5093 5967 5107
rect 5933 5074 5947 5088
rect 5853 5033 5867 5047
rect 5913 4993 5927 5007
rect 5833 4953 5847 4967
rect 5833 4893 5847 4907
rect 5893 4893 5907 4907
rect 5773 4793 5787 4807
rect 5813 4793 5827 4807
rect 5853 4772 5867 4786
rect 5833 4753 5847 4767
rect 5773 4733 5787 4747
rect 5753 4554 5767 4568
rect 5753 4513 5767 4527
rect 5753 4433 5767 4447
rect 5813 4633 5827 4647
rect 5793 4573 5807 4587
rect 5873 4753 5887 4767
rect 5853 4653 5867 4667
rect 5893 4633 5907 4647
rect 5873 4573 5887 4587
rect 6013 5272 6027 5286
rect 5993 5173 6007 5187
rect 5993 5113 6007 5127
rect 5973 4973 5987 4987
rect 5993 4953 6007 4967
rect 6213 5613 6227 5627
rect 6293 5613 6307 5627
rect 6173 5594 6187 5608
rect 6253 5594 6267 5608
rect 6173 5553 6187 5567
rect 6233 5552 6247 5566
rect 6273 5553 6287 5567
rect 6153 5513 6167 5527
rect 6293 5533 6307 5547
rect 6273 5493 6287 5507
rect 6193 5453 6207 5467
rect 6153 5433 6167 5447
rect 6173 5393 6187 5407
rect 6053 5373 6067 5387
rect 6113 5374 6127 5388
rect 6053 5313 6067 5327
rect 6093 5313 6107 5327
rect 6093 5133 6107 5147
rect 6053 5093 6067 5107
rect 6093 5093 6107 5107
rect 6153 5313 6167 5327
rect 6133 5233 6147 5247
rect 6133 5193 6147 5207
rect 6133 5133 6147 5147
rect 6133 5092 6147 5106
rect 6073 4993 6087 5007
rect 6073 4953 6087 4967
rect 6013 4893 6027 4907
rect 6053 4893 6067 4907
rect 5953 4853 5967 4867
rect 6033 4853 6047 4867
rect 5953 4813 5967 4827
rect 5813 4512 5827 4526
rect 5792 4452 5806 4466
rect 5813 4453 5827 4467
rect 5773 4353 5787 4367
rect 5893 4513 5907 4527
rect 5893 4413 5907 4427
rect 5853 4393 5867 4407
rect 5933 4493 5947 4507
rect 5993 4812 6007 4826
rect 6073 4753 6087 4767
rect 6053 4733 6067 4747
rect 6053 4712 6067 4726
rect 6073 4693 6087 4707
rect 6013 4673 6027 4687
rect 6053 4673 6067 4687
rect 5973 4653 5987 4667
rect 6052 4593 6066 4607
rect 6073 4593 6087 4607
rect 6293 5433 6307 5447
rect 6253 5374 6267 5388
rect 6313 5393 6327 5407
rect 6233 5332 6247 5346
rect 6313 5333 6327 5347
rect 6293 5293 6307 5307
rect 6193 5253 6207 5267
rect 6293 5213 6307 5227
rect 6253 5173 6267 5187
rect 6213 5133 6227 5147
rect 6193 5093 6207 5107
rect 6173 5073 6187 5087
rect 6293 5153 6307 5167
rect 6253 5113 6267 5127
rect 6173 4993 6187 5007
rect 6213 4993 6227 5007
rect 6193 4973 6207 4987
rect 6173 4953 6187 4967
rect 6173 4913 6187 4927
rect 6113 4853 6127 4867
rect 6133 4793 6147 4807
rect 6193 4793 6207 4807
rect 6113 4773 6127 4787
rect 6133 4753 6147 4767
rect 6113 4693 6127 4707
rect 5993 4554 6007 4568
rect 6033 4554 6047 4568
rect 6053 4512 6067 4526
rect 6113 4533 6127 4547
rect 6012 4493 6026 4507
rect 6033 4493 6047 4507
rect 6093 4493 6107 4507
rect 5973 4413 5987 4427
rect 5913 4352 5927 4366
rect 5953 4353 5967 4367
rect 5893 4333 5907 4347
rect 5873 4313 5887 4327
rect 5753 4233 5767 4247
rect 5833 4173 5847 4187
rect 5753 4113 5767 4127
rect 5633 3953 5647 3967
rect 5613 3873 5627 3887
rect 5453 3772 5467 3786
rect 5552 3713 5566 3727
rect 5573 3713 5587 3727
rect 5553 3633 5567 3647
rect 5573 3593 5587 3607
rect 5413 3573 5427 3587
rect 5533 3573 5547 3587
rect 5493 3533 5507 3547
rect 5413 3513 5427 3527
rect 5553 3553 5567 3567
rect 5552 3513 5566 3527
rect 5293 3473 5307 3486
rect 5293 3472 5307 3473
rect 5353 3472 5367 3486
rect 5313 3453 5327 3467
rect 5393 3433 5407 3447
rect 5333 3413 5347 3427
rect 5273 3393 5287 3407
rect 5093 3313 5107 3327
rect 5093 3272 5107 3286
rect 5193 3272 5207 3286
rect 4973 3252 4987 3266
rect 5393 3393 5407 3407
rect 5373 3274 5387 3288
rect 5053 3233 5067 3247
rect 5093 3233 5107 3247
rect 5333 3233 5347 3247
rect 5053 3153 5067 3167
rect 5033 3113 5047 3127
rect 5573 3512 5587 3526
rect 5433 3493 5447 3507
rect 5413 3353 5427 3367
rect 5413 3313 5427 3327
rect 5513 3472 5527 3486
rect 5553 3473 5567 3487
rect 5473 3453 5487 3467
rect 5553 3433 5567 3447
rect 5493 3373 5507 3387
rect 5473 3313 5487 3327
rect 5433 3293 5447 3307
rect 5453 3272 5467 3286
rect 5193 3213 5207 3227
rect 5333 3212 5347 3226
rect 5392 3213 5406 3227
rect 5413 3213 5427 3227
rect 5193 3133 5207 3147
rect 5233 3113 5247 3127
rect 5093 3093 5107 3107
rect 5173 3093 5187 3107
rect 5073 2974 5087 2988
rect 4933 2933 4947 2947
rect 4953 2873 4967 2887
rect 5093 2873 5107 2887
rect 4793 2653 4807 2667
rect 4913 2653 4927 2667
rect 4933 2633 4947 2647
rect 4853 2593 4867 2607
rect 4813 2513 4827 2527
rect 4833 2473 4847 2487
rect 4893 2474 4907 2488
rect 4933 2473 4947 2487
rect 4873 2432 4887 2446
rect 4833 2393 4847 2407
rect 4853 2373 4867 2387
rect 4913 2373 4927 2387
rect 4893 2333 4907 2347
rect 4713 2313 4727 2327
rect 4773 2313 4787 2327
rect 4833 2313 4847 2327
rect 4873 2313 4887 2327
rect 4793 2273 4807 2287
rect 4793 2193 4807 2207
rect 4733 2173 4747 2187
rect 4633 2073 4647 2087
rect 4613 1993 4627 2007
rect 4693 1973 4707 1987
rect 4733 1973 4747 1987
rect 4773 1973 4787 1987
rect 4593 1953 4607 1967
rect 4573 1873 4587 1887
rect 4613 1853 4627 1867
rect 4573 1833 4587 1847
rect 4513 1773 4527 1787
rect 4553 1773 4567 1787
rect 4373 1692 4387 1706
rect 4433 1692 4447 1706
rect 4333 1613 4347 1627
rect 4313 1513 4327 1527
rect 4233 1493 4247 1507
rect 4233 1434 4247 1448
rect 4293 1434 4307 1448
rect 4213 1392 4227 1406
rect 4232 1293 4246 1307
rect 4253 1293 4267 1307
rect 4193 1214 4207 1228
rect 4293 1253 4307 1267
rect 4273 1214 4287 1228
rect 4373 1533 4387 1547
rect 4493 1693 4507 1707
rect 4473 1473 4487 1487
rect 4413 1434 4427 1448
rect 4453 1434 4467 1448
rect 4393 1392 4407 1406
rect 4453 1333 4467 1347
rect 4333 1293 4347 1307
rect 4433 1293 4447 1307
rect 4193 1173 4207 1187
rect 4253 1153 4267 1167
rect 4333 1172 4347 1186
rect 4413 1172 4427 1186
rect 4293 1133 4307 1147
rect 4373 1093 4387 1107
rect 4213 1033 4227 1047
rect 4293 1033 4307 1047
rect 4213 993 4227 1007
rect 4193 973 4207 987
rect 4193 952 4207 966
rect 4153 914 4167 928
rect 4113 853 4127 867
rect 4193 853 4207 867
rect 4233 973 4247 987
rect 4253 914 4267 928
rect 4233 872 4247 886
rect 4353 872 4367 886
rect 4233 773 4247 787
rect 4313 753 4327 767
rect 4073 733 4087 747
rect 4173 733 4187 747
rect 4213 733 4227 747
rect 4033 693 4047 707
rect 4113 694 4127 708
rect 4313 732 4327 746
rect 4353 694 4367 708
rect 4133 652 4147 666
rect 4173 652 4187 666
rect 4213 652 4227 666
rect 4253 652 4267 666
rect 4033 613 4047 627
rect 4113 573 4127 587
rect 3973 553 3987 567
rect 3873 533 3887 547
rect 4053 453 4067 467
rect 3853 433 3867 447
rect 3653 394 3667 408
rect 3793 394 3807 408
rect 3633 352 3647 366
rect 3773 313 3787 327
rect 3713 293 3727 307
rect 3653 174 3667 188
rect 3693 174 3707 188
rect 3973 394 3987 408
rect 4033 394 4047 408
rect 3913 313 3927 327
rect 3853 293 3867 307
rect 3793 173 3807 187
rect 4153 394 4167 408
rect 4053 352 4067 366
rect 4093 352 4107 366
rect 4133 352 4147 366
rect 4033 293 4047 307
rect 4033 253 4047 267
rect 3913 213 3927 227
rect 3673 113 3687 127
rect 3793 132 3807 146
rect 3833 132 3847 146
rect 3993 174 4007 188
rect 4033 174 4047 188
rect 4073 174 4087 188
rect 4173 174 4187 188
rect 4393 1073 4407 1087
rect 4533 1533 4547 1547
rect 4673 1933 4687 1947
rect 4693 1873 4707 1887
rect 4793 1873 4807 1887
rect 4933 2353 4947 2367
rect 4853 2273 4867 2287
rect 4913 2273 4927 2287
rect 5013 2853 5027 2867
rect 5233 3073 5247 3087
rect 5293 3093 5307 3107
rect 5193 2972 5207 2986
rect 5273 2973 5287 2987
rect 5233 2953 5247 2967
rect 5213 2933 5227 2947
rect 5113 2833 5127 2847
rect 5173 2833 5187 2847
rect 5093 2813 5107 2827
rect 5053 2774 5067 2788
rect 4993 2733 5007 2747
rect 5133 2793 5147 2807
rect 5113 2773 5127 2787
rect 4993 2613 5007 2627
rect 4973 2533 4987 2547
rect 5093 2732 5107 2746
rect 5053 2713 5067 2727
rect 5113 2713 5127 2727
rect 5053 2673 5067 2687
rect 5093 2673 5107 2687
rect 5013 2493 5027 2507
rect 5053 2493 5067 2507
rect 5313 3053 5327 3067
rect 5253 2893 5267 2907
rect 5233 2793 5247 2807
rect 5153 2733 5167 2747
rect 5133 2533 5147 2547
rect 5093 2473 5107 2487
rect 4993 2432 5007 2446
rect 5033 2432 5047 2446
rect 4973 2353 4987 2367
rect 5093 2433 5107 2447
rect 5073 2393 5087 2407
rect 5013 2353 5027 2367
rect 4993 2273 5007 2287
rect 4913 2212 4927 2226
rect 4953 2193 4967 2207
rect 4853 2113 4867 2127
rect 4873 2073 4887 2087
rect 4853 1912 4867 1926
rect 4613 1813 4627 1827
rect 4653 1813 4667 1827
rect 4753 1813 4767 1827
rect 4833 1813 4847 1827
rect 4753 1712 4767 1726
rect 4913 1912 4927 1926
rect 4873 1873 4887 1887
rect 4953 1873 4967 1887
rect 4973 1813 4987 1827
rect 4873 1714 4887 1728
rect 4953 1713 4967 1727
rect 4853 1653 4867 1667
rect 4913 1653 4927 1667
rect 4833 1573 4847 1587
rect 4613 1513 4627 1527
rect 4753 1513 4767 1527
rect 4553 1453 4567 1467
rect 4613 1453 4627 1467
rect 4573 1434 4587 1448
rect 4653 1433 4667 1447
rect 4693 1434 4707 1448
rect 4793 1434 4807 1448
rect 4893 1553 4907 1567
rect 4953 1553 4967 1567
rect 4853 1493 4867 1507
rect 4593 1373 4607 1387
rect 4553 1333 4567 1347
rect 4553 1253 4567 1267
rect 4513 1214 4527 1228
rect 4593 1214 4607 1228
rect 4613 1172 4627 1186
rect 4573 1153 4587 1167
rect 4513 1133 4527 1147
rect 4493 1033 4507 1047
rect 4533 953 4547 967
rect 4413 914 4427 928
rect 4473 914 4487 928
rect 4513 914 4527 928
rect 4553 872 4567 886
rect 4433 853 4447 867
rect 4513 853 4527 867
rect 4413 813 4427 827
rect 4553 813 4567 827
rect 4433 773 4447 787
rect 4513 773 4527 787
rect 4393 753 4407 767
rect 4393 694 4407 708
rect 4533 733 4547 747
rect 4493 694 4507 708
rect 4833 1433 4847 1447
rect 4693 1393 4707 1407
rect 4693 1293 4707 1307
rect 4673 1213 4687 1227
rect 4673 1172 4687 1186
rect 4673 1113 4687 1127
rect 4653 1093 4667 1107
rect 4773 1392 4787 1406
rect 4833 1392 4847 1406
rect 4753 1293 4767 1307
rect 4733 1253 4747 1267
rect 4793 1253 4807 1267
rect 4753 1214 4767 1228
rect 4733 1053 4747 1067
rect 4693 993 4707 1007
rect 4773 993 4787 1007
rect 4673 973 4687 987
rect 4753 953 4767 967
rect 4733 914 4747 928
rect 4633 872 4647 886
rect 4773 872 4787 886
rect 4613 833 4627 847
rect 4673 833 4687 847
rect 4713 813 4727 827
rect 4633 773 4647 787
rect 4613 733 4627 747
rect 4573 693 4587 707
rect 4593 693 4607 707
rect 4433 652 4447 666
rect 4513 652 4527 666
rect 4633 693 4647 707
rect 4753 693 4767 707
rect 4613 652 4627 666
rect 4653 652 4667 666
rect 4693 573 4707 587
rect 4493 553 4507 567
rect 4373 453 4387 467
rect 4233 394 4247 408
rect 4273 394 4287 408
rect 4313 394 4327 408
rect 4353 394 4367 408
rect 4393 394 4407 408
rect 4433 394 4447 408
rect 4653 433 4667 447
rect 4233 353 4247 367
rect 4293 352 4307 366
rect 4493 393 4507 407
rect 4393 353 4407 367
rect 4453 352 4467 366
rect 4353 313 4367 327
rect 4613 394 4627 408
rect 4593 313 4607 327
rect 4673 393 4687 407
rect 4653 293 4667 307
rect 4613 253 4627 267
rect 4473 213 4487 227
rect 4513 213 4527 227
rect 4253 193 4267 207
rect 4373 193 4387 207
rect 4013 132 4027 146
rect 4073 133 4087 147
rect 4293 174 4307 188
rect 4333 174 4347 188
rect 3713 113 3727 127
rect 4193 132 4207 146
rect 4253 132 4267 146
rect 3693 93 3707 107
rect 3733 93 3747 107
rect 4153 93 4167 107
rect 4433 173 4447 187
rect 4533 174 4547 188
rect 4653 213 4667 227
rect 4633 193 4647 207
rect 4613 173 4627 187
rect 4873 1473 4887 1487
rect 4973 1473 4987 1487
rect 4913 1434 4927 1448
rect 4973 1433 4987 1447
rect 4933 1392 4947 1406
rect 4973 1392 4987 1406
rect 4873 1373 4887 1387
rect 4973 1353 4987 1367
rect 4933 1293 4947 1307
rect 5133 2453 5147 2467
rect 5113 2313 5127 2327
rect 5133 2293 5147 2307
rect 5033 2253 5047 2267
rect 5093 2254 5107 2268
rect 5193 2732 5207 2746
rect 5233 2673 5247 2687
rect 5293 2893 5307 2907
rect 5313 2873 5327 2887
rect 5453 3193 5467 3207
rect 5353 3173 5367 3187
rect 5393 3173 5407 3187
rect 5433 3173 5447 3187
rect 5413 3153 5427 3167
rect 5413 3113 5427 3127
rect 5393 3093 5407 3107
rect 5373 3013 5387 3027
rect 5453 3113 5467 3127
rect 5453 3092 5467 3106
rect 5393 2952 5407 2966
rect 5433 2953 5447 2967
rect 5413 2913 5427 2927
rect 5353 2873 5367 2887
rect 5333 2773 5347 2787
rect 5373 2732 5387 2746
rect 5293 2633 5307 2647
rect 5353 2633 5367 2647
rect 5273 2613 5287 2627
rect 5213 2573 5227 2587
rect 5173 2452 5187 2466
rect 5473 3032 5487 3046
rect 5453 2873 5467 2887
rect 5533 3333 5547 3347
rect 5513 3293 5527 3307
rect 5513 3093 5527 3107
rect 5513 3053 5527 3067
rect 5493 2993 5507 3007
rect 5733 4073 5747 4087
rect 5793 4073 5807 4087
rect 5673 4053 5687 4067
rect 5713 4034 5727 4048
rect 5753 4034 5767 4048
rect 5693 3993 5707 4007
rect 5753 3973 5767 3987
rect 5733 3953 5747 3967
rect 5773 3953 5787 3967
rect 5673 3913 5687 3927
rect 5713 3893 5727 3907
rect 5813 3893 5827 3907
rect 5793 3873 5807 3887
rect 5773 3853 5787 3867
rect 5813 3833 5827 3847
rect 5793 3813 5807 3827
rect 5773 3793 5787 3807
rect 5733 3753 5747 3767
rect 5773 3733 5787 3747
rect 5673 3713 5687 3727
rect 5753 3713 5767 3727
rect 5653 3673 5667 3687
rect 5633 3593 5647 3607
rect 5613 3533 5627 3547
rect 5733 3653 5747 3667
rect 5693 3633 5707 3647
rect 5673 3553 5687 3567
rect 5633 3513 5647 3527
rect 5713 3473 5727 3487
rect 5613 3413 5627 3427
rect 5673 3413 5687 3427
rect 5613 3392 5627 3406
rect 5593 3353 5607 3367
rect 5573 3333 5587 3347
rect 5613 3293 5627 3307
rect 5613 3253 5627 3267
rect 5553 3213 5567 3227
rect 5593 3213 5607 3227
rect 5593 3133 5607 3147
rect 5593 3053 5607 3067
rect 5633 3133 5647 3147
rect 5633 3093 5647 3107
rect 5613 3013 5627 3027
rect 5493 2893 5507 2907
rect 5573 2952 5587 2966
rect 5533 2873 5547 2887
rect 5493 2853 5507 2867
rect 5473 2833 5487 2847
rect 5533 2833 5547 2847
rect 5453 2773 5467 2787
rect 5493 2774 5507 2788
rect 5593 2873 5607 2887
rect 5573 2773 5587 2787
rect 5433 2633 5447 2647
rect 5553 2732 5567 2746
rect 5533 2673 5547 2687
rect 5413 2593 5427 2607
rect 5453 2593 5467 2607
rect 5373 2573 5387 2587
rect 5373 2513 5387 2527
rect 5353 2493 5367 2507
rect 5352 2454 5366 2468
rect 5373 2453 5387 2467
rect 5213 2433 5227 2447
rect 5173 2393 5187 2407
rect 5213 2393 5227 2407
rect 5173 2353 5187 2367
rect 5213 2353 5227 2367
rect 5053 2213 5067 2227
rect 5033 2193 5047 2207
rect 5033 2033 5047 2047
rect 5093 2113 5107 2127
rect 5073 2093 5087 2107
rect 5093 2033 5107 2047
rect 5513 2613 5527 2627
rect 5613 2732 5627 2746
rect 5493 2533 5507 2547
rect 5593 2533 5607 2547
rect 5473 2513 5487 2527
rect 5673 3353 5687 3367
rect 5773 3693 5787 3707
rect 5973 4334 5987 4348
rect 5913 4273 5927 4287
rect 5933 4253 5947 4267
rect 5933 4232 5947 4246
rect 5893 4153 5907 4167
rect 5993 4273 6007 4287
rect 5973 4253 5987 4267
rect 6013 4253 6027 4267
rect 5953 4173 5967 4187
rect 5953 4033 5967 4047
rect 5873 3992 5887 4006
rect 5913 3992 5927 4006
rect 5833 3813 5847 3827
rect 6173 4593 6187 4607
rect 6173 4554 6187 4568
rect 6213 4753 6227 4767
rect 6273 4993 6287 5007
rect 6253 4853 6267 4867
rect 6373 5653 6387 5667
rect 6373 5594 6387 5608
rect 6413 5594 6427 5608
rect 6473 5753 6487 5767
rect 6353 5553 6367 5567
rect 6433 5552 6447 5566
rect 6392 5533 6406 5547
rect 6413 5533 6427 5547
rect 6353 5453 6367 5467
rect 6373 5433 6387 5447
rect 6333 5313 6347 5327
rect 6413 5493 6427 5507
rect 6393 5413 6407 5427
rect 6493 5593 6507 5607
rect 6593 6427 6607 6428
rect 6593 6414 6607 6427
rect 6653 6414 6667 6428
rect 6713 6414 6727 6428
rect 6753 6414 6767 6428
rect 6673 6372 6687 6386
rect 6733 6372 6747 6386
rect 6613 6173 6627 6187
rect 6713 6153 6727 6167
rect 6613 6133 6627 6147
rect 6653 6114 6667 6128
rect 6633 6053 6647 6067
rect 6673 6053 6687 6067
rect 6573 5933 6587 5947
rect 6553 5852 6567 5866
rect 6633 5894 6647 5908
rect 6573 5813 6587 5827
rect 6653 5813 6667 5827
rect 6653 5792 6667 5806
rect 6633 5673 6647 5687
rect 6573 5653 6587 5667
rect 6573 5613 6587 5627
rect 6493 5553 6507 5567
rect 6473 5513 6487 5527
rect 6453 5433 6467 5447
rect 6453 5412 6467 5426
rect 6413 5374 6427 5388
rect 6393 5333 6407 5346
rect 6393 5332 6407 5333
rect 6433 5332 6447 5346
rect 6473 5313 6487 5327
rect 6373 5253 6387 5267
rect 6413 5213 6427 5227
rect 6353 5173 6367 5187
rect 6373 5074 6387 5088
rect 6553 5593 6567 5607
rect 6593 5594 6607 5608
rect 6613 5553 6627 5567
rect 6573 5513 6587 5527
rect 6553 5393 6567 5407
rect 6533 5373 6547 5387
rect 6653 5473 6667 5487
rect 6633 5393 6647 5407
rect 6553 5332 6567 5346
rect 6593 5332 6607 5346
rect 6633 5313 6647 5327
rect 6533 5273 6547 5287
rect 6613 5233 6627 5247
rect 6513 5213 6527 5227
rect 6593 5213 6607 5227
rect 6473 5193 6487 5207
rect 6453 5173 6467 5187
rect 6432 5133 6446 5147
rect 6453 5133 6467 5147
rect 6433 5073 6447 5087
rect 6353 5032 6367 5046
rect 6393 4993 6407 5007
rect 6313 4913 6327 4927
rect 6333 4893 6347 4907
rect 6273 4812 6287 4826
rect 6313 4812 6327 4826
rect 6353 4812 6367 4826
rect 6233 4713 6247 4727
rect 6333 4693 6347 4707
rect 6233 4653 6247 4667
rect 6313 4633 6327 4647
rect 6253 4554 6267 4568
rect 6173 4513 6187 4527
rect 6133 4473 6147 4487
rect 6193 4473 6207 4487
rect 6113 4433 6127 4447
rect 6113 4393 6127 4407
rect 6073 4373 6087 4387
rect 6053 4333 6067 4347
rect 6033 4233 6047 4247
rect 5933 3973 5947 3987
rect 5973 3973 5987 3987
rect 5913 3833 5927 3847
rect 5953 3953 5967 3967
rect 6093 4333 6107 4347
rect 6093 4293 6107 4307
rect 6073 4193 6087 4207
rect 6073 4133 6087 4147
rect 6013 4113 6027 4127
rect 6173 4293 6187 4307
rect 6113 4193 6127 4207
rect 6153 4233 6167 4247
rect 6133 4153 6147 4167
rect 6093 4053 6107 4067
rect 6113 4034 6127 4048
rect 6013 3993 6027 4007
rect 6053 3992 6067 4006
rect 5993 3913 6007 3927
rect 5973 3893 5987 3907
rect 5953 3813 5967 3827
rect 5813 3753 5827 3767
rect 5813 3693 5827 3707
rect 5813 3593 5827 3607
rect 5813 3553 5827 3567
rect 5793 3533 5807 3547
rect 5893 3772 5907 3786
rect 5953 3713 5967 3727
rect 5853 3653 5867 3667
rect 5853 3573 5867 3587
rect 5833 3533 5847 3547
rect 5833 3472 5847 3486
rect 5873 3472 5887 3486
rect 5833 3413 5847 3427
rect 5773 3393 5787 3407
rect 5753 3373 5767 3387
rect 5753 3294 5767 3308
rect 5693 3253 5707 3267
rect 5713 3233 5727 3247
rect 5692 3193 5706 3207
rect 5713 3193 5727 3207
rect 5673 3133 5687 3147
rect 5653 2813 5667 2827
rect 5693 3113 5707 3127
rect 5773 3173 5787 3187
rect 5733 3113 5747 3127
rect 5773 3113 5787 3127
rect 5733 3073 5747 3087
rect 5713 3053 5727 3067
rect 5733 3033 5747 3047
rect 5773 3033 5787 3047
rect 5913 3613 5927 3627
rect 5953 3593 5967 3607
rect 5933 3553 5947 3567
rect 6133 3973 6147 3987
rect 6113 3953 6127 3967
rect 6133 3913 6147 3927
rect 6113 3873 6127 3887
rect 5993 3853 6007 3867
rect 6053 3853 6067 3867
rect 6093 3833 6107 3847
rect 6053 3814 6067 3828
rect 6133 3773 6147 3787
rect 6093 3753 6107 3767
rect 5993 3733 6007 3747
rect 5993 3712 6007 3726
rect 6213 4453 6227 4467
rect 6293 4512 6307 4526
rect 6273 4453 6287 4467
rect 6313 4473 6327 4487
rect 6233 4433 6247 4447
rect 6233 4393 6247 4407
rect 6273 4393 6287 4407
rect 6313 4393 6327 4407
rect 6213 4333 6227 4347
rect 6213 4272 6227 4286
rect 6193 4173 6207 4187
rect 6293 4373 6307 4387
rect 6373 4673 6387 4687
rect 6353 4593 6367 4607
rect 6353 4554 6367 4568
rect 6373 4512 6387 4526
rect 6353 4472 6367 4486
rect 6333 4333 6347 4347
rect 6313 4292 6327 4306
rect 6353 4293 6367 4307
rect 6313 4273 6327 4287
rect 6273 4252 6287 4266
rect 6233 4193 6247 4207
rect 6173 4033 6187 4047
rect 6173 4012 6187 4026
rect 6173 3973 6187 3987
rect 6173 3913 6187 3927
rect 6173 3873 6187 3887
rect 6213 4113 6227 4127
rect 6333 4173 6347 4187
rect 6233 4034 6247 4048
rect 6313 4073 6327 4087
rect 6213 3993 6227 4007
rect 6293 3993 6307 4007
rect 6253 3953 6267 3967
rect 6273 3933 6287 3947
rect 6253 3913 6267 3927
rect 6233 3873 6247 3887
rect 6273 3873 6287 3887
rect 6213 3833 6227 3847
rect 6173 3812 6187 3826
rect 6293 3813 6307 3827
rect 6113 3713 6127 3727
rect 6093 3693 6107 3707
rect 6253 3772 6267 3786
rect 6213 3753 6227 3767
rect 6213 3713 6227 3727
rect 6133 3673 6147 3687
rect 6172 3673 6186 3687
rect 6193 3673 6207 3687
rect 5993 3653 6007 3667
rect 6093 3653 6107 3667
rect 6013 3553 6027 3567
rect 6073 3553 6087 3567
rect 5973 3533 5987 3547
rect 6013 3514 6027 3528
rect 6073 3514 6087 3528
rect 5993 3472 6007 3486
rect 5933 3433 5947 3447
rect 5893 3413 5907 3427
rect 6073 3473 6087 3487
rect 6113 3593 6127 3607
rect 6213 3613 6227 3627
rect 6153 3593 6167 3607
rect 6093 3413 6107 3427
rect 6033 3373 6047 3387
rect 6093 3373 6107 3387
rect 6133 3533 6147 3547
rect 6213 3573 6227 3587
rect 6273 3693 6287 3707
rect 6253 3573 6267 3587
rect 6113 3333 6127 3347
rect 6153 3472 6167 3486
rect 6193 3472 6207 3486
rect 6233 3473 6247 3486
rect 6233 3472 6247 3473
rect 6153 3433 6167 3447
rect 6133 3313 6147 3327
rect 6093 3293 6107 3307
rect 5853 3213 5867 3227
rect 6093 3272 6107 3286
rect 6133 3274 6147 3288
rect 6093 3193 6107 3207
rect 5833 3173 5847 3187
rect 5953 3173 5967 3187
rect 5693 3013 5707 3027
rect 5793 2973 5807 2987
rect 5693 2913 5707 2927
rect 5793 2873 5807 2887
rect 5813 2812 5827 2826
rect 5753 2793 5767 2807
rect 5693 2774 5707 2788
rect 5673 2713 5687 2727
rect 5813 2673 5827 2687
rect 6093 3133 6107 3147
rect 5933 3093 5947 3107
rect 6133 3213 6147 3227
rect 6133 3153 6147 3167
rect 6213 3413 6227 3427
rect 6173 3273 6187 3287
rect 6173 3233 6187 3247
rect 6133 3113 6147 3127
rect 6073 3073 6087 3087
rect 6112 3073 6126 3087
rect 6133 3073 6147 3087
rect 5912 2973 5926 2987
rect 5933 2974 5947 2988
rect 6133 3033 6147 3047
rect 6193 3133 6207 3147
rect 6073 2972 6087 2986
rect 6113 2972 6127 2986
rect 6073 2913 6087 2927
rect 5893 2873 5907 2887
rect 5973 2873 5987 2887
rect 5953 2813 5967 2827
rect 6173 2933 6187 2947
rect 6153 2913 6167 2927
rect 6193 2893 6207 2907
rect 6133 2853 6147 2867
rect 6033 2833 6047 2847
rect 6073 2833 6087 2847
rect 5933 2732 5947 2746
rect 5973 2733 5987 2747
rect 5873 2713 5887 2727
rect 5853 2693 5867 2707
rect 5833 2653 5847 2667
rect 6013 2693 6027 2707
rect 5932 2653 5946 2667
rect 5953 2653 5967 2667
rect 5733 2573 5747 2587
rect 5633 2513 5647 2527
rect 5713 2513 5727 2527
rect 5492 2493 5506 2507
rect 5513 2494 5527 2508
rect 5573 2494 5587 2508
rect 5633 2492 5647 2506
rect 5473 2433 5487 2447
rect 5453 2313 5467 2327
rect 5333 2293 5347 2307
rect 5193 2254 5207 2268
rect 5173 2073 5187 2087
rect 5253 2254 5267 2268
rect 5293 2254 5307 2268
rect 5553 2453 5567 2467
rect 5513 2413 5527 2427
rect 5493 2353 5507 2367
rect 5493 2313 5507 2327
rect 5413 2273 5427 2287
rect 5473 2273 5487 2287
rect 5373 2253 5387 2267
rect 5213 2212 5227 2226
rect 5273 2212 5287 2226
rect 5313 2212 5327 2226
rect 5353 2212 5367 2226
rect 5353 2133 5367 2147
rect 5073 2013 5087 2027
rect 5153 1993 5167 2007
rect 5052 1953 5066 1967
rect 5073 1954 5087 1968
rect 5113 1973 5127 1987
rect 5093 1912 5107 1926
rect 5113 1893 5127 1907
rect 5053 1813 5067 1827
rect 5173 1973 5187 1987
rect 5173 1933 5187 1947
rect 5173 1893 5187 1907
rect 5213 1953 5227 1967
rect 5333 1954 5347 1968
rect 5193 1833 5207 1847
rect 5173 1813 5187 1827
rect 5153 1793 5167 1807
rect 5153 1734 5167 1748
rect 5113 1533 5127 1547
rect 5013 1433 5027 1447
rect 5073 1434 5087 1448
rect 5173 1453 5187 1467
rect 5013 1412 5027 1426
rect 5153 1412 5167 1426
rect 5273 1873 5287 1887
rect 5333 1793 5347 1807
rect 5233 1733 5247 1747
rect 5273 1734 5287 1748
rect 5213 1693 5227 1707
rect 5293 1692 5307 1706
rect 5333 1573 5347 1587
rect 5393 2033 5407 2047
rect 5373 1993 5387 2007
rect 5393 1973 5407 1987
rect 5373 1932 5387 1946
rect 5373 1793 5387 1807
rect 5433 2212 5447 2226
rect 5533 2353 5547 2367
rect 5533 2313 5547 2327
rect 5513 2213 5527 2227
rect 5513 2173 5527 2187
rect 5493 2153 5507 2167
rect 5493 2113 5507 2127
rect 5873 2593 5887 2607
rect 5753 2553 5767 2567
rect 5873 2553 5887 2567
rect 5733 2493 5747 2507
rect 5712 2453 5726 2467
rect 5733 2454 5747 2468
rect 5873 2454 5887 2468
rect 5953 2613 5967 2627
rect 6013 2473 6027 2487
rect 5633 2433 5647 2447
rect 5933 2433 5947 2447
rect 5633 2393 5647 2407
rect 5693 2353 5707 2367
rect 5633 2333 5647 2347
rect 5593 2313 5607 2327
rect 5633 2293 5647 2307
rect 5653 2254 5667 2268
rect 5573 2153 5587 2167
rect 5553 2133 5567 2147
rect 5512 2093 5526 2107
rect 5533 2093 5547 2107
rect 5633 2193 5647 2207
rect 5713 2333 5727 2347
rect 5873 2313 5887 2327
rect 5733 2253 5747 2267
rect 5773 2254 5787 2268
rect 5813 2254 5827 2268
rect 5753 2213 5767 2227
rect 5713 2173 5727 2187
rect 5693 2153 5707 2167
rect 5613 2113 5627 2127
rect 5733 2093 5747 2107
rect 5613 2073 5627 2087
rect 5593 2053 5607 2067
rect 5853 2213 5867 2227
rect 5833 2153 5847 2167
rect 5813 2093 5827 2107
rect 5753 2073 5767 2087
rect 5733 2013 5747 2027
rect 5453 1974 5467 1988
rect 5433 1833 5447 1847
rect 5773 1974 5787 1988
rect 5613 1953 5627 1967
rect 5713 1953 5727 1967
rect 5733 1932 5747 1946
rect 5793 1893 5807 1907
rect 5713 1853 5727 1867
rect 5473 1793 5487 1807
rect 5413 1773 5427 1787
rect 5453 1773 5467 1787
rect 5413 1734 5427 1748
rect 5453 1734 5467 1748
rect 5393 1693 5407 1707
rect 5373 1653 5387 1667
rect 5393 1613 5407 1627
rect 5513 1673 5527 1687
rect 5493 1653 5507 1667
rect 5433 1593 5447 1607
rect 5393 1573 5407 1587
rect 5353 1533 5367 1547
rect 5253 1412 5267 1426
rect 5653 1712 5667 1726
rect 5653 1673 5667 1687
rect 5813 1714 5827 1728
rect 5873 2093 5887 2107
rect 5913 2393 5927 2407
rect 5933 2273 5947 2287
rect 5913 2253 5927 2267
rect 5993 2392 6007 2406
rect 5973 2373 5987 2387
rect 5993 2333 6007 2347
rect 6113 2813 6127 2827
rect 6193 2813 6207 2827
rect 6173 2793 6187 2807
rect 6073 2774 6087 2788
rect 6053 2753 6067 2767
rect 6193 2753 6207 2767
rect 6193 2693 6207 2707
rect 6053 2593 6067 2607
rect 6133 2673 6147 2687
rect 6093 2633 6107 2647
rect 6073 2573 6087 2587
rect 6073 2533 6087 2547
rect 6153 2593 6167 2607
rect 6133 2513 6147 2527
rect 6233 3313 6247 3327
rect 6253 3293 6267 3307
rect 6233 3273 6247 3287
rect 6233 3153 6247 3167
rect 6233 3053 6247 3067
rect 6213 2553 6227 2567
rect 6213 2513 6227 2527
rect 6113 2474 6127 2488
rect 6153 2474 6167 2488
rect 6193 2473 6207 2487
rect 6133 2432 6147 2446
rect 6033 2293 6047 2307
rect 5993 2254 6007 2268
rect 6053 2273 6067 2287
rect 6033 2253 6047 2267
rect 5953 2193 5967 2207
rect 5913 2173 5927 2187
rect 5873 2013 5887 2027
rect 5853 1893 5867 1907
rect 5933 2013 5947 2027
rect 5973 2113 5987 2127
rect 5953 1973 5967 1987
rect 5893 1953 5907 1967
rect 6013 2173 6027 2187
rect 6133 2373 6147 2387
rect 6113 2293 6127 2307
rect 6173 2293 6187 2307
rect 6193 2273 6207 2287
rect 6093 2253 6107 2267
rect 6133 2254 6147 2268
rect 6173 2254 6187 2268
rect 6293 3673 6307 3687
rect 6313 3653 6327 3667
rect 6373 4253 6387 4267
rect 6373 4193 6387 4207
rect 6413 4713 6427 4727
rect 6453 5032 6467 5046
rect 6453 4973 6467 4987
rect 6493 5113 6507 5127
rect 6493 5074 6507 5088
rect 6553 5074 6567 5088
rect 6513 4913 6527 4927
rect 6493 4873 6507 4887
rect 6573 4993 6587 5007
rect 6553 4953 6567 4967
rect 6533 4893 6547 4907
rect 6573 4933 6587 4947
rect 6533 4872 6547 4886
rect 6473 4853 6487 4867
rect 6493 4812 6507 4826
rect 6513 4713 6527 4727
rect 6433 4633 6447 4647
rect 6453 4554 6467 4568
rect 6433 4512 6447 4526
rect 6433 4473 6447 4487
rect 6473 4453 6487 4467
rect 6493 4433 6507 4447
rect 6473 4334 6487 4348
rect 6513 4393 6527 4407
rect 6493 4293 6507 4307
rect 6433 4273 6447 4287
rect 6453 4253 6467 4267
rect 6493 4253 6507 4267
rect 6433 4213 6447 4227
rect 6413 4193 6427 4207
rect 6393 4073 6407 4087
rect 6433 4073 6447 4087
rect 6373 4033 6387 4047
rect 6433 4033 6447 4047
rect 6353 3993 6367 4007
rect 6393 3992 6407 4006
rect 6433 3993 6447 4007
rect 6393 3933 6407 3947
rect 6373 3893 6387 3907
rect 6353 3873 6367 3887
rect 6353 3833 6367 3847
rect 6373 3813 6387 3827
rect 6433 3853 6447 3867
rect 6493 4213 6507 4227
rect 6493 4133 6507 4147
rect 6473 4113 6487 4127
rect 6493 4093 6507 4107
rect 6553 4852 6567 4866
rect 6633 5153 6647 5167
rect 6613 5013 6627 5027
rect 6693 5973 6707 5987
rect 6693 5894 6707 5908
rect 6693 5853 6707 5867
rect 6753 6313 6767 6327
rect 6853 6153 6867 6167
rect 6813 6114 6827 6128
rect 6753 6072 6767 6086
rect 6793 6072 6807 6086
rect 6733 6033 6747 6047
rect 6793 6033 6807 6047
rect 6833 6033 6847 6047
rect 6773 5852 6787 5866
rect 6713 5673 6727 5687
rect 6693 5593 6707 5607
rect 6753 5613 6767 5627
rect 6813 5833 6827 5847
rect 6813 5733 6827 5747
rect 6793 5633 6807 5647
rect 6773 5593 6787 5607
rect 6693 5553 6707 5567
rect 6733 5552 6747 5566
rect 6713 5513 6727 5527
rect 6693 5372 6707 5386
rect 6673 5233 6687 5247
rect 6693 5213 6707 5227
rect 6893 5633 6907 5647
rect 6833 5594 6847 5608
rect 6873 5594 6887 5608
rect 6913 5594 6927 5608
rect 6813 5493 6827 5507
rect 6733 5413 6747 5427
rect 6793 5413 6807 5427
rect 6773 5374 6787 5388
rect 6813 5374 6827 5388
rect 6953 5553 6967 5567
rect 6853 5374 6867 5388
rect 6733 5273 6747 5287
rect 6713 5093 6727 5107
rect 6693 5074 6707 5088
rect 6733 5074 6747 5088
rect 6633 4873 6647 4887
rect 6593 4853 6607 4867
rect 6753 5033 6767 5047
rect 6712 5013 6726 5027
rect 6733 5013 6747 5027
rect 6713 4973 6727 4987
rect 6653 4854 6667 4868
rect 6693 4853 6707 4867
rect 6633 4793 6647 4807
rect 6593 4593 6607 4607
rect 6673 4593 6687 4607
rect 6573 4553 6587 4567
rect 6613 4554 6627 4568
rect 6573 4513 6587 4527
rect 6553 4473 6567 4487
rect 6553 4413 6567 4427
rect 6533 4093 6547 4107
rect 6633 4433 6647 4447
rect 6633 4393 6647 4407
rect 6633 4334 6647 4348
rect 6553 4073 6567 4087
rect 6593 4273 6607 4287
rect 6613 4233 6627 4247
rect 6493 4053 6507 4067
rect 6473 3953 6487 3967
rect 6433 3832 6447 3846
rect 6473 3833 6487 3847
rect 6373 3773 6387 3787
rect 6353 3733 6367 3747
rect 6413 3772 6427 3786
rect 6453 3772 6467 3786
rect 6553 4034 6567 4048
rect 6593 4033 6607 4047
rect 6533 3992 6547 4006
rect 6573 3953 6587 3967
rect 6513 3933 6527 3947
rect 6553 3933 6567 3947
rect 6513 3893 6527 3907
rect 6453 3751 6467 3765
rect 6433 3733 6447 3747
rect 6413 3713 6427 3727
rect 6373 3653 6387 3667
rect 6413 3653 6427 3667
rect 6373 3573 6387 3587
rect 6293 3533 6307 3547
rect 6333 3534 6347 3548
rect 6293 3512 6307 3526
rect 6333 3513 6347 3527
rect 6413 3513 6427 3527
rect 6313 3473 6327 3487
rect 6353 3472 6367 3486
rect 6393 3472 6407 3486
rect 6373 3453 6387 3467
rect 6293 3413 6307 3427
rect 6293 3373 6307 3387
rect 6273 3193 6287 3207
rect 6353 3294 6367 3308
rect 6393 3393 6407 3407
rect 6313 3253 6327 3267
rect 6313 3173 6327 3187
rect 6333 3113 6347 3127
rect 6313 3093 6327 3107
rect 6493 3772 6507 3786
rect 6533 3853 6547 3867
rect 6693 4513 6707 4527
rect 6693 4453 6707 4467
rect 6793 5072 6807 5086
rect 6773 4993 6787 5007
rect 6753 4973 6767 4987
rect 6813 5013 6827 5027
rect 6853 5113 6867 5127
rect 6933 5513 6947 5527
rect 6893 5493 6907 5507
rect 6933 5473 6947 5487
rect 6893 5373 6907 5387
rect 6953 5373 6967 5387
rect 6893 5333 6907 5347
rect 6953 5333 6967 5347
rect 6933 5213 6947 5227
rect 6893 5153 6907 5167
rect 6913 5133 6927 5147
rect 6873 5093 6887 5107
rect 6853 5013 6867 5027
rect 6833 4933 6847 4947
rect 6773 4793 6787 4807
rect 6813 4793 6827 4807
rect 6833 4633 6847 4647
rect 6733 4553 6747 4567
rect 6773 4554 6787 4568
rect 6813 4554 6827 4568
rect 6753 4512 6767 4526
rect 6773 4493 6787 4507
rect 6793 4453 6807 4467
rect 6673 4053 6687 4067
rect 6753 4233 6767 4247
rect 6753 4193 6767 4207
rect 6653 3992 6667 4006
rect 6693 3992 6707 4006
rect 6793 4133 6807 4147
rect 6793 4053 6807 4067
rect 6793 3993 6807 4007
rect 6653 3933 6667 3947
rect 6633 3873 6647 3887
rect 6573 3853 6587 3867
rect 6633 3852 6647 3866
rect 6593 3814 6607 3828
rect 6573 3772 6587 3786
rect 6613 3772 6627 3786
rect 6533 3753 6547 3767
rect 6513 3713 6527 3727
rect 6473 3693 6487 3707
rect 6473 3672 6487 3686
rect 6513 3653 6527 3667
rect 6433 3433 6447 3447
rect 6433 3333 6447 3347
rect 6393 3073 6407 3087
rect 6553 3633 6567 3647
rect 6673 3873 6687 3887
rect 6753 3893 6767 3907
rect 6733 3873 6747 3887
rect 6773 3814 6787 3828
rect 6693 3773 6707 3787
rect 6653 3673 6667 3687
rect 6553 3533 6567 3547
rect 6473 3513 6487 3527
rect 6533 3513 6547 3527
rect 6513 3413 6527 3427
rect 6493 3373 6507 3387
rect 6473 3333 6487 3347
rect 6593 3473 6607 3487
rect 6593 3393 6607 3407
rect 6553 3332 6567 3346
rect 6433 3273 6447 3287
rect 6433 3133 6447 3147
rect 6413 3053 6427 3067
rect 6573 3313 6587 3327
rect 6513 3213 6527 3227
rect 6553 3213 6567 3227
rect 6493 3193 6507 3207
rect 6472 3153 6486 3167
rect 6493 3153 6507 3167
rect 6473 3113 6487 3127
rect 6453 3073 6467 3087
rect 6433 3033 6447 3047
rect 6413 2994 6427 3008
rect 6453 2994 6467 3008
rect 6313 2952 6327 2966
rect 6433 2952 6447 2966
rect 6293 2933 6307 2947
rect 6413 2933 6427 2947
rect 6293 2833 6307 2847
rect 6413 2873 6427 2887
rect 6393 2833 6407 2847
rect 6273 2773 6287 2787
rect 6313 2774 6327 2788
rect 6453 2873 6467 2887
rect 6473 2853 6487 2867
rect 6473 2813 6487 2827
rect 6473 2774 6487 2788
rect 6553 3173 6567 3187
rect 6673 3652 6687 3666
rect 6753 3772 6767 3786
rect 6793 3773 6807 3787
rect 6753 3713 6767 3727
rect 6673 3513 6687 3527
rect 6733 3472 6747 3486
rect 6753 3453 6767 3467
rect 6653 3413 6667 3427
rect 6633 3313 6647 3327
rect 6613 3293 6627 3307
rect 6693 3433 6707 3447
rect 6733 3433 6747 3447
rect 6673 3373 6687 3387
rect 6693 3294 6707 3308
rect 6613 3253 6627 3267
rect 6593 3153 6607 3167
rect 6673 3252 6687 3266
rect 6733 3252 6747 3266
rect 6633 3193 6647 3207
rect 6673 3193 6687 3207
rect 6773 3413 6787 3427
rect 6773 3373 6787 3387
rect 6693 3173 6707 3187
rect 6753 3173 6767 3187
rect 6833 4073 6847 4087
rect 6873 4873 6887 4887
rect 6913 4973 6927 4987
rect 6893 4853 6907 4867
rect 6893 4393 6907 4407
rect 6953 5113 6967 5127
rect 6953 5092 6967 5106
rect 6953 4793 6967 4807
rect 6933 4554 6947 4568
rect 6913 4133 6927 4147
rect 6913 4073 6927 4087
rect 6893 4033 6907 4047
rect 6833 3993 6847 4007
rect 6893 3993 6907 4007
rect 6893 3933 6907 3947
rect 6953 4133 6967 4147
rect 6953 3893 6967 3907
rect 6933 3873 6947 3887
rect 6913 3853 6927 3867
rect 6853 3813 6867 3827
rect 6912 3814 6926 3828
rect 6933 3813 6947 3827
rect 6833 3653 6847 3667
rect 6873 3773 6887 3787
rect 6933 3773 6947 3787
rect 6893 3633 6907 3647
rect 6853 3513 6867 3527
rect 6953 3613 6967 3627
rect 6932 3513 6946 3527
rect 6953 3513 6967 3527
rect 6953 3492 6967 3506
rect 6833 3453 6847 3467
rect 6813 3373 6827 3387
rect 6813 3294 6827 3308
rect 6893 3472 6907 3486
rect 6953 3433 6967 3447
rect 6873 3373 6887 3387
rect 6853 3293 6867 3307
rect 6633 3133 6647 3147
rect 6693 3133 6707 3147
rect 6773 3133 6787 3147
rect 6613 3093 6627 3107
rect 6552 3053 6566 3067
rect 6573 3053 6587 3067
rect 6673 3053 6687 3067
rect 6533 2952 6547 2966
rect 6573 2893 6587 2907
rect 6653 2893 6667 2907
rect 6273 2733 6287 2747
rect 6373 2733 6387 2747
rect 6373 2693 6387 2707
rect 6413 2673 6427 2687
rect 6293 2653 6307 2667
rect 6333 2653 6347 2667
rect 6293 2613 6307 2627
rect 6253 2474 6267 2488
rect 6393 2613 6407 2627
rect 6373 2553 6387 2567
rect 6333 2473 6347 2487
rect 6273 2432 6287 2446
rect 6293 2413 6307 2427
rect 6273 2333 6287 2347
rect 6253 2273 6267 2287
rect 6093 2153 6107 2167
rect 6073 2133 6087 2147
rect 6113 2133 6127 2147
rect 6133 2093 6147 2107
rect 6213 2213 6227 2227
rect 6153 2073 6167 2087
rect 6133 2053 6147 2067
rect 6193 2033 6207 2047
rect 6113 2013 6127 2027
rect 5993 1953 6007 1967
rect 5913 1893 5927 1907
rect 5953 1853 5967 1867
rect 5953 1773 5967 1787
rect 5893 1714 5907 1728
rect 5653 1593 5667 1607
rect 5553 1533 5567 1547
rect 5593 1533 5607 1547
rect 5633 1533 5647 1547
rect 5513 1473 5527 1487
rect 5493 1454 5507 1468
rect 5593 1473 5607 1487
rect 5013 1373 5027 1387
rect 5233 1393 5247 1407
rect 5093 1373 5107 1387
rect 5073 1353 5087 1367
rect 5013 1313 5027 1327
rect 5053 1313 5067 1327
rect 4993 1273 5007 1287
rect 4973 1214 4987 1228
rect 4913 1033 4927 1047
rect 4853 973 4867 987
rect 4813 914 4827 928
rect 4873 914 4887 928
rect 4853 872 4867 886
rect 4813 833 4827 847
rect 4853 813 4867 827
rect 4813 793 4827 807
rect 4753 394 4767 408
rect 5053 1273 5067 1287
rect 5133 1253 5147 1267
rect 5153 1172 5167 1186
rect 5113 1093 5127 1107
rect 5193 1053 5207 1067
rect 5013 813 5027 827
rect 5713 1493 5727 1507
rect 5753 1454 5767 1468
rect 5653 1373 5667 1387
rect 5793 1373 5807 1387
rect 5853 1673 5867 1687
rect 6053 1972 6067 1986
rect 6073 1953 6087 1967
rect 6153 1993 6167 2007
rect 6093 1912 6107 1926
rect 6053 1773 6067 1787
rect 6173 1893 6187 1907
rect 6173 1813 6187 1827
rect 6073 1734 6087 1748
rect 6133 1753 6147 1767
rect 5993 1713 6007 1727
rect 6053 1692 6067 1706
rect 6093 1673 6107 1687
rect 5993 1653 6007 1667
rect 5953 1573 5967 1587
rect 5953 1533 5967 1547
rect 5913 1434 5927 1448
rect 5913 1413 5927 1427
rect 6073 1413 6087 1427
rect 5453 1293 5467 1307
rect 5593 1293 5607 1307
rect 5813 1293 5827 1307
rect 5953 1293 5967 1307
rect 6053 1293 6067 1307
rect 5293 1214 5307 1228
rect 5333 1213 5347 1227
rect 5373 1214 5387 1228
rect 5413 1214 5427 1228
rect 5593 1253 5607 1267
rect 5353 1194 5367 1208
rect 5273 1172 5287 1186
rect 5313 973 5327 987
rect 5493 1194 5507 1208
rect 5433 1133 5447 1147
rect 5373 1113 5387 1127
rect 5593 1173 5607 1187
rect 5733 1173 5747 1187
rect 5533 1053 5547 1067
rect 5793 1053 5807 1067
rect 5473 993 5487 1007
rect 5413 953 5427 967
rect 5393 914 5407 928
rect 5313 853 5327 867
rect 5233 813 5247 827
rect 5193 793 5207 807
rect 4893 773 4907 787
rect 5093 773 5107 787
rect 5093 693 5107 707
rect 4993 672 5007 686
rect 5153 613 5167 627
rect 5013 493 5027 507
rect 4873 453 4887 467
rect 4853 394 4867 408
rect 4693 352 4707 366
rect 4733 352 4747 366
rect 4673 193 4687 207
rect 4713 193 4727 207
rect 4353 132 4367 146
rect 4433 132 4447 146
rect 4473 132 4487 146
rect 4513 132 4527 146
rect 4553 132 4567 146
rect 4633 132 4647 146
rect 4693 132 4707 146
rect 4733 132 4747 146
rect 4813 293 4827 307
rect 4793 173 4807 187
rect 4793 132 4807 146
rect 4953 394 4967 408
rect 4973 352 4987 366
rect 4933 293 4947 307
rect 4873 273 4887 287
rect 4933 213 4947 227
rect 4873 174 4887 188
rect 4853 132 4867 146
rect 4873 113 4887 127
rect 4393 93 4407 107
rect 4693 93 4707 107
rect 4773 93 4787 107
rect 4293 73 4307 87
rect 5053 433 5067 447
rect 5033 393 5047 407
rect 5033 352 5047 366
rect 5093 394 5107 408
rect 5233 773 5247 787
rect 5233 713 5247 727
rect 5253 694 5267 708
rect 5473 914 5487 928
rect 5413 873 5427 887
rect 5493 872 5507 886
rect 5393 853 5407 867
rect 5413 833 5427 847
rect 5333 793 5347 807
rect 5593 913 5607 927
rect 5533 793 5547 807
rect 5493 773 5507 787
rect 5413 733 5427 747
rect 5453 694 5467 708
rect 5233 652 5247 666
rect 5333 652 5347 666
rect 5473 652 5487 666
rect 5253 533 5267 547
rect 5293 533 5307 547
rect 5113 352 5127 366
rect 5153 353 5167 367
rect 5053 293 5067 307
rect 5773 873 5787 887
rect 5693 833 5707 847
rect 5773 813 5787 827
rect 6093 1393 6107 1407
rect 6093 1273 6107 1287
rect 6153 1734 6167 1748
rect 6333 2393 6347 2407
rect 6313 2293 6327 2307
rect 6353 2333 6367 2347
rect 6493 2713 6507 2727
rect 6473 2553 6487 2567
rect 6453 2513 6467 2527
rect 6613 2774 6627 2788
rect 6513 2633 6527 2647
rect 6593 2713 6607 2727
rect 6633 2693 6647 2707
rect 6613 2633 6627 2647
rect 6593 2573 6607 2587
rect 6533 2533 6547 2547
rect 6513 2513 6527 2527
rect 6593 2493 6607 2507
rect 6513 2473 6527 2487
rect 6573 2474 6587 2488
rect 6673 2493 6687 2507
rect 6433 2432 6447 2446
rect 6473 2432 6487 2446
rect 6533 2433 6547 2447
rect 6393 2413 6407 2427
rect 6453 2413 6467 2427
rect 6553 2413 6567 2427
rect 6453 2373 6467 2387
rect 6373 2313 6387 2327
rect 6413 2313 6427 2327
rect 6333 2273 6347 2287
rect 6293 2253 6307 2267
rect 6293 2213 6307 2227
rect 6253 2113 6267 2127
rect 6233 2093 6247 2107
rect 6253 2053 6267 2067
rect 6293 2053 6307 2067
rect 6233 1912 6247 1926
rect 6313 2033 6327 2047
rect 6273 1954 6287 1968
rect 6373 1912 6387 1926
rect 6253 1873 6267 1887
rect 6293 1873 6307 1887
rect 6233 1793 6247 1807
rect 6153 1553 6167 1567
rect 6133 1473 6147 1487
rect 6153 1412 6167 1426
rect 6133 1393 6147 1407
rect 6113 1253 6127 1267
rect 6073 1213 6087 1227
rect 5873 993 5887 1007
rect 5833 953 5847 967
rect 5813 913 5827 927
rect 5813 833 5827 847
rect 5633 793 5647 807
rect 5673 733 5687 747
rect 5633 694 5647 708
rect 5573 653 5587 667
rect 6093 1172 6107 1186
rect 5953 1133 5967 1147
rect 5913 973 5927 987
rect 6053 973 6067 987
rect 5893 953 5907 967
rect 5893 872 5907 886
rect 6033 833 6047 847
rect 6113 973 6127 987
rect 6113 872 6127 886
rect 6153 1253 6167 1267
rect 6213 1653 6227 1667
rect 6333 1853 6347 1867
rect 6433 2273 6447 2287
rect 6433 2053 6447 2067
rect 6533 2293 6547 2307
rect 6493 2254 6507 2268
rect 6513 2212 6527 2226
rect 6513 2133 6527 2147
rect 6473 2093 6487 2107
rect 6453 1992 6467 2006
rect 6413 1913 6427 1927
rect 6413 1852 6427 1866
rect 6333 1832 6347 1846
rect 6393 1833 6407 1847
rect 6313 1753 6327 1767
rect 6313 1692 6327 1706
rect 6253 1493 6267 1507
rect 6293 1493 6307 1507
rect 6213 1473 6227 1487
rect 6193 1133 6207 1147
rect 6173 1033 6187 1047
rect 6373 1753 6387 1767
rect 6473 1954 6487 1968
rect 6533 2053 6547 2067
rect 6613 2474 6627 2488
rect 6833 3113 6847 3127
rect 6793 3073 6807 3087
rect 6713 2994 6727 3008
rect 6753 2994 6767 3008
rect 6853 3033 6867 3047
rect 6713 2933 6727 2947
rect 6753 2933 6767 2947
rect 6713 2853 6727 2867
rect 6693 2473 6707 2487
rect 6633 2432 6647 2446
rect 6693 2433 6707 2447
rect 6673 2393 6687 2407
rect 6693 2373 6707 2387
rect 6593 2353 6607 2367
rect 6813 2952 6827 2966
rect 6773 2893 6787 2907
rect 6793 2774 6807 2788
rect 6853 2952 6867 2966
rect 6833 2773 6847 2787
rect 6773 2732 6787 2746
rect 6733 2693 6747 2707
rect 6833 2733 6847 2747
rect 6813 2693 6827 2707
rect 6773 2633 6787 2647
rect 6833 2613 6847 2627
rect 6753 2513 6767 2527
rect 6833 2513 6847 2527
rect 6733 2433 6747 2447
rect 6793 2493 6807 2507
rect 6913 3293 6927 3307
rect 6893 3093 6907 3107
rect 6873 2673 6887 2687
rect 6853 2493 6867 2507
rect 6953 2653 6967 2667
rect 6913 2553 6927 2567
rect 6813 2432 6827 2446
rect 6853 2432 6867 2446
rect 6893 2432 6907 2446
rect 6773 2393 6787 2407
rect 6753 2353 6767 2367
rect 6613 2333 6627 2347
rect 6713 2333 6727 2347
rect 6593 2213 6607 2227
rect 6593 2113 6607 2127
rect 6533 1993 6547 2007
rect 6453 1893 6467 1907
rect 6493 1893 6507 1907
rect 6553 1893 6567 1907
rect 6533 1873 6547 1887
rect 6473 1833 6487 1847
rect 6433 1813 6447 1827
rect 6493 1813 6507 1827
rect 6553 1813 6567 1827
rect 6473 1793 6487 1807
rect 6433 1753 6447 1767
rect 6413 1734 6427 1748
rect 6353 1693 6367 1707
rect 6433 1692 6447 1706
rect 6473 1692 6487 1706
rect 6753 2293 6767 2307
rect 6653 2254 6667 2268
rect 6693 2254 6707 2268
rect 6753 2253 6767 2267
rect 6673 2212 6687 2226
rect 6713 2212 6727 2226
rect 6753 2093 6767 2107
rect 6733 2073 6747 2087
rect 6793 2353 6807 2367
rect 6613 2033 6627 2047
rect 6733 2033 6747 2047
rect 6773 2033 6787 2047
rect 6513 1793 6527 1807
rect 6593 1793 6607 1807
rect 6493 1473 6507 1487
rect 6353 1453 6367 1467
rect 6433 1453 6447 1467
rect 6333 1433 6347 1447
rect 6273 1273 6287 1287
rect 6413 1433 6427 1447
rect 6353 1353 6367 1367
rect 6313 1253 6327 1267
rect 6233 1214 6247 1228
rect 6333 1172 6347 1186
rect 6213 1073 6227 1087
rect 6293 1033 6307 1047
rect 6193 973 6207 987
rect 6333 993 6347 1007
rect 6153 914 6167 928
rect 6273 914 6287 928
rect 6173 872 6187 886
rect 6273 853 6287 867
rect 5913 793 5927 807
rect 6093 793 6107 807
rect 6133 793 6147 807
rect 6173 793 6187 807
rect 5833 733 5847 747
rect 5873 733 5887 747
rect 5773 694 5787 708
rect 5833 694 5847 708
rect 5873 694 5887 708
rect 6173 693 6187 707
rect 5673 632 5687 646
rect 5613 513 5627 527
rect 5393 433 5407 447
rect 5493 433 5507 447
rect 5553 433 5567 447
rect 5253 353 5267 367
rect 5753 593 5767 607
rect 6033 653 6047 667
rect 5873 632 5887 646
rect 6233 713 6247 727
rect 6213 693 6227 707
rect 6193 673 6207 687
rect 6173 613 6187 627
rect 6113 533 6127 547
rect 6033 513 6047 527
rect 5773 493 5787 507
rect 5813 493 5827 507
rect 5613 414 5627 428
rect 5673 414 5687 428
rect 5513 372 5527 386
rect 5673 372 5687 386
rect 5253 313 5267 327
rect 5493 313 5507 327
rect 5653 313 5667 327
rect 5213 233 5227 247
rect 5053 213 5067 227
rect 5393 233 5407 247
rect 5013 174 5027 188
rect 5173 173 5187 187
rect 4933 113 4947 127
rect 5073 132 5087 146
rect 5313 133 5327 147
rect 5873 253 5887 267
rect 6273 613 6287 627
rect 6233 473 6247 487
rect 6213 433 6227 447
rect 6173 413 6187 427
rect 6233 413 6247 427
rect 6253 393 6267 407
rect 6113 353 6127 367
rect 6193 352 6207 366
rect 6153 333 6167 347
rect 5953 233 5967 247
rect 5693 154 5707 168
rect 5833 153 5847 167
rect 5673 113 5687 127
rect 5733 112 5747 126
rect 5573 93 5587 107
rect 5913 112 5927 126
rect 5953 112 5967 126
rect 6113 152 6127 166
rect 6313 893 6327 907
rect 6313 593 6327 607
rect 6293 513 6307 527
rect 6293 413 6307 427
rect 6393 1353 6407 1367
rect 6393 1253 6407 1267
rect 6533 1753 6547 1767
rect 6773 1993 6787 2007
rect 6713 1912 6727 1926
rect 6653 1893 6667 1907
rect 6633 1833 6647 1847
rect 6653 1773 6667 1787
rect 6753 1754 6767 1768
rect 6673 1733 6687 1747
rect 6713 1734 6727 1748
rect 6753 1733 6767 1747
rect 6653 1692 6667 1706
rect 6833 2254 6847 2268
rect 6913 2293 6927 2307
rect 6853 2212 6867 2226
rect 6893 2213 6907 2227
rect 6933 2213 6947 2227
rect 6913 2113 6927 2127
rect 6853 2033 6867 2047
rect 6813 1954 6827 1968
rect 6893 1954 6907 1968
rect 6833 1912 6847 1926
rect 6813 1753 6827 1767
rect 6533 1633 6547 1647
rect 6613 1633 6627 1647
rect 6513 1433 6527 1447
rect 6433 1392 6447 1406
rect 6473 1392 6487 1406
rect 6453 1253 6467 1267
rect 6493 1214 6507 1228
rect 6473 1172 6487 1186
rect 6573 1573 6587 1587
rect 6653 1573 6667 1587
rect 6553 1433 6567 1447
rect 6693 1692 6707 1706
rect 6733 1692 6747 1706
rect 6793 1692 6807 1706
rect 6873 1873 6887 1887
rect 6893 1753 6907 1767
rect 6833 1733 6847 1747
rect 6932 1734 6946 1748
rect 6953 1733 6967 1747
rect 6833 1673 6847 1687
rect 6693 1593 6707 1607
rect 6813 1593 6827 1607
rect 6633 1434 6647 1448
rect 6673 1434 6687 1448
rect 6573 1392 6587 1406
rect 6553 1253 6567 1267
rect 6553 1214 6567 1228
rect 6553 1173 6567 1187
rect 6533 1113 6547 1127
rect 6513 1053 6527 1067
rect 6413 993 6427 1007
rect 6393 973 6407 987
rect 6453 953 6467 967
rect 6353 872 6367 886
rect 6393 872 6407 886
rect 6333 493 6347 507
rect 6333 433 6347 447
rect 6313 394 6327 408
rect 6653 1392 6667 1406
rect 6653 1333 6667 1347
rect 6613 1313 6627 1327
rect 6673 1253 6687 1267
rect 6653 1233 6667 1247
rect 6713 1553 6727 1567
rect 6773 1473 6787 1487
rect 6813 1434 6827 1448
rect 6713 1393 6727 1407
rect 6793 1392 6807 1406
rect 6913 1692 6927 1706
rect 6953 1693 6967 1707
rect 6873 1673 6887 1687
rect 6853 1313 6867 1327
rect 6893 1573 6907 1587
rect 6673 1193 6687 1207
rect 6713 1214 6727 1228
rect 6773 1214 6787 1228
rect 6813 1214 6827 1228
rect 6613 1172 6627 1186
rect 6693 1172 6707 1186
rect 6753 1172 6767 1186
rect 6793 1172 6807 1186
rect 6873 1213 6887 1227
rect 6713 1133 6727 1147
rect 6673 1113 6687 1127
rect 6573 953 6587 967
rect 6653 933 6667 947
rect 6633 914 6647 928
rect 6473 733 6487 747
rect 6453 713 6467 727
rect 6513 694 6527 708
rect 6573 694 6587 708
rect 6713 1093 6727 1107
rect 6833 1093 6847 1107
rect 6673 873 6687 887
rect 6573 633 6587 647
rect 6393 533 6407 547
rect 6573 533 6587 547
rect 6353 413 6367 427
rect 6373 394 6387 408
rect 6433 393 6447 407
rect 6293 333 6307 347
rect 6373 333 6387 347
rect 6353 293 6367 307
rect 6373 253 6387 267
rect 6293 233 6307 247
rect 6353 213 6367 227
rect 6433 293 6447 307
rect 6413 173 6427 187
rect 6393 153 6407 167
rect 6413 133 6427 147
rect 6253 113 6267 127
rect 6473 493 6487 507
rect 6493 433 6507 447
rect 6513 394 6527 408
rect 6673 633 6687 647
rect 6853 1073 6867 1087
rect 6753 973 6767 987
rect 6793 933 6807 947
rect 6773 872 6787 886
rect 6813 833 6827 847
rect 6713 613 6727 627
rect 6813 613 6827 627
rect 6693 533 6707 547
rect 6793 533 6807 547
rect 6633 394 6647 408
rect 6793 473 6807 487
rect 6773 433 6787 447
rect 6733 394 6747 408
rect 6493 353 6507 367
rect 6713 352 6727 366
rect 6553 313 6567 327
rect 6633 313 6647 327
rect 6713 313 6727 327
rect 6553 253 6567 267
rect 6473 213 6487 227
rect 6773 193 6787 207
rect 6513 174 6527 188
rect 6553 174 6567 188
rect 6673 174 6687 188
rect 6493 132 6507 146
rect 6873 833 6887 847
rect 6893 433 6907 447
rect 6933 1673 6947 1687
rect 6933 1333 6947 1347
rect 6813 273 6827 287
rect 6833 193 6847 207
rect 6913 313 6927 327
rect 6953 313 6967 327
rect 6913 273 6927 287
rect 6853 132 6867 146
rect 6933 132 6947 146
rect 6533 113 6547 127
rect 5833 73 5847 87
rect 6013 73 6027 87
rect 6453 73 6467 87
rect 2473 33 2487 47
rect 3613 33 3627 47
rect 4893 33 4907 47
rect 5033 33 5047 47
<< metal3 >>
rect 307 6516 333 6524
rect 2727 6456 2973 6464
rect 3027 6456 3153 6464
rect 3287 6456 4133 6464
rect 4147 6456 4213 6464
rect 4447 6456 4913 6464
rect 4967 6456 5113 6464
rect 6347 6456 6453 6464
rect 2407 6436 2493 6444
rect 3007 6436 3473 6444
rect 3967 6436 3993 6444
rect 5587 6436 5993 6444
rect 6007 6436 6473 6444
rect 6547 6436 6873 6444
rect 167 6416 273 6424
rect 287 6417 413 6425
rect -24 6376 113 6384
rect 436 6344 444 6433
rect 827 6416 913 6424
rect 1387 6416 1733 6424
rect 2036 6420 2453 6424
rect 2033 6416 2453 6420
rect 947 6396 1013 6404
rect 1347 6397 1773 6405
rect 2033 6407 2047 6416
rect 2547 6416 2613 6424
rect 2667 6416 2813 6424
rect 2887 6416 2953 6424
rect 3207 6417 3233 6425
rect 3347 6417 3373 6425
rect 3627 6416 3753 6424
rect 3807 6416 3873 6424
rect 493 6384 507 6393
rect 487 6380 507 6384
rect 487 6376 504 6380
rect 2647 6375 2713 6383
rect 2996 6384 3004 6414
rect 3896 6416 3913 6424
rect 3896 6404 3904 6416
rect 4047 6416 4093 6424
rect 4287 6416 4373 6424
rect 4487 6416 4504 6424
rect 3527 6396 3904 6404
rect 4496 6404 4504 6416
rect 4527 6416 4613 6424
rect 4707 6416 4753 6424
rect 5007 6417 5073 6425
rect 5127 6417 5153 6425
rect 5207 6417 5253 6425
rect 4496 6396 4604 6404
rect 2847 6376 3004 6384
rect 3596 6386 3604 6396
rect 4596 6386 4604 6396
rect 5296 6404 5304 6414
rect 5187 6396 5304 6404
rect 5456 6404 5464 6414
rect 5527 6416 5633 6424
rect 5647 6416 5733 6424
rect 5807 6416 5893 6424
rect 5967 6416 6053 6424
rect 6147 6416 6212 6424
rect 6247 6417 6293 6425
rect 6607 6417 6653 6425
rect 6727 6417 6753 6425
rect 5456 6396 5644 6404
rect 3247 6376 3313 6384
rect 3787 6376 3933 6384
rect 4387 6375 4413 6383
rect 5107 6376 5193 6384
rect 5327 6376 5433 6384
rect 5507 6376 5613 6384
rect 5636 6384 5644 6396
rect 5636 6376 5653 6384
rect 5907 6375 5933 6383
rect 6227 6375 6273 6383
rect 6687 6375 6733 6383
rect 2487 6356 2533 6364
rect 3647 6356 3993 6364
rect 4227 6356 4253 6364
rect 6047 6356 6153 6364
rect 6167 6356 6373 6364
rect 436 6336 473 6344
rect 887 6336 913 6344
rect 927 6336 1333 6344
rect 1347 6336 1373 6344
rect 2787 6336 2973 6344
rect 3167 6336 3733 6344
rect 3887 6336 3973 6344
rect 5447 6336 5973 6344
rect 367 6316 573 6324
rect 2327 6316 2833 6324
rect 3007 6316 3133 6324
rect 3147 6316 3453 6324
rect 4047 6316 4453 6324
rect 4947 6316 5233 6324
rect 5887 6316 6753 6324
rect 4147 6296 4293 6304
rect 4647 6296 5273 6304
rect 5807 6296 6233 6304
rect 587 6276 973 6284
rect 987 6276 1433 6284
rect 1867 6276 2093 6284
rect 2207 6276 2824 6284
rect 2816 6267 2824 6276
rect 4787 6276 5173 6284
rect 5327 6276 5493 6284
rect 5707 6276 6224 6284
rect 1807 6256 2433 6264
rect 2827 6256 3173 6264
rect 3187 6256 3373 6264
rect 3387 6256 4013 6264
rect 6216 6264 6224 6276
rect 6216 6256 6313 6264
rect 687 6236 713 6244
rect 4687 6236 5513 6244
rect 5747 6236 5893 6244
rect 5907 6236 6113 6244
rect 827 6216 933 6224
rect 1447 6216 1893 6224
rect 2227 6216 3193 6224
rect 4696 6216 4813 6224
rect 987 6196 1073 6204
rect 1747 6196 1864 6204
rect 1247 6176 1513 6184
rect 1856 6184 1864 6196
rect 1916 6196 2193 6204
rect 1916 6184 1924 6196
rect 2447 6196 3113 6204
rect 4696 6204 4704 6216
rect 4867 6216 5193 6224
rect 5207 6216 5233 6224
rect 5467 6216 5693 6224
rect 3987 6196 4704 6204
rect 5787 6196 5853 6204
rect 1856 6176 1924 6184
rect 2307 6176 2413 6184
rect 3347 6176 4333 6184
rect 4727 6176 4773 6184
rect 5127 6176 5333 6184
rect 5407 6176 5713 6184
rect 6507 6176 6613 6184
rect 1027 6156 1493 6164
rect 1507 6156 1833 6164
rect 1847 6156 1993 6164
rect 2287 6156 2533 6164
rect 2547 6156 2673 6164
rect 2727 6156 2793 6164
rect 2807 6156 3313 6164
rect 3907 6156 4233 6164
rect 4307 6156 4773 6164
rect 4827 6156 5173 6164
rect 5947 6156 6033 6164
rect 6727 6156 6853 6164
rect 847 6136 893 6144
rect 1147 6136 1433 6144
rect 1647 6136 1713 6144
rect 2047 6136 2313 6144
rect 4847 6136 4933 6144
rect 6367 6136 6613 6144
rect -24 6116 13 6124
rect 187 6117 253 6125
rect 547 6117 653 6125
rect 947 6117 973 6125
rect 1516 6116 1793 6124
rect 796 6104 804 6114
rect 796 6096 864 6104
rect 27 6075 133 6083
rect 267 6075 313 6083
rect 727 6076 813 6084
rect 856 6084 864 6096
rect 1516 6104 1524 6116
rect 2187 6117 2273 6125
rect 2367 6116 2544 6124
rect 1487 6096 1524 6104
rect 2536 6104 2544 6116
rect 2587 6116 2873 6124
rect 2947 6116 3073 6124
rect 3127 6116 3273 6124
rect 3287 6117 3313 6125
rect 3427 6116 3553 6124
rect 3607 6117 3653 6125
rect 3707 6116 3753 6124
rect 4087 6116 4173 6124
rect 2536 6096 2684 6104
rect 856 6076 993 6084
rect 1527 6076 1653 6084
rect 1747 6076 1813 6084
rect 1867 6076 1973 6084
rect 2027 6076 2293 6084
rect 2676 6086 2684 6096
rect 3936 6087 3944 6114
rect 4327 6117 4393 6125
rect 4527 6117 4553 6125
rect 4576 6116 4593 6124
rect 4576 6104 4584 6116
rect 4647 6117 4693 6125
rect 5007 6117 5073 6125
rect 5287 6117 5353 6125
rect 5527 6116 5573 6124
rect 5756 6116 5793 6124
rect 5756 6104 5764 6116
rect 5987 6117 6033 6125
rect 6087 6117 6153 6125
rect 6247 6117 6273 6125
rect 6407 6117 6453 6125
rect 6667 6116 6813 6124
rect 4416 6096 4584 6104
rect 5676 6096 5764 6104
rect 2347 6075 2433 6083
rect 2527 6075 2573 6083
rect 2747 6076 2913 6084
rect 3107 6075 3172 6083
rect 3207 6076 3253 6084
rect 3627 6075 3713 6083
rect 3787 6076 3913 6084
rect 3936 6076 3953 6087
rect 3940 6073 3953 6076
rect 4416 6086 4424 6096
rect 4047 6076 4173 6084
rect 4187 6075 4213 6083
rect 4267 6075 4293 6083
rect 4487 6075 4573 6083
rect 4807 6075 4833 6083
rect 4887 6075 4913 6083
rect 5267 6076 5313 6084
rect 5676 6084 5684 6096
rect 6316 6087 6324 6114
rect 5647 6076 5684 6084
rect 5727 6075 5773 6083
rect 5907 6075 5953 6083
rect 6187 6076 6233 6084
rect 6316 6076 6333 6087
rect 6320 6073 6333 6076
rect 6767 6075 6793 6083
rect 427 6056 493 6064
rect 1067 6056 1504 6064
rect 947 6036 993 6044
rect 1047 6036 1093 6044
rect 1387 6036 1413 6044
rect 1427 6036 1473 6044
rect 1496 6044 1504 6056
rect 4327 6056 4373 6064
rect 4627 6056 4673 6064
rect 5067 6056 5153 6064
rect 5347 6056 5493 6064
rect 6647 6056 6673 6064
rect 1496 6036 2453 6044
rect 2947 6036 2993 6044
rect 4027 6036 4093 6044
rect 4107 6036 4813 6044
rect 5107 6036 5373 6044
rect 5447 6036 5693 6044
rect 5827 6036 6033 6044
rect 6636 6044 6644 6053
rect 6487 6036 6644 6044
rect 6747 6036 6793 6044
rect 6807 6036 6833 6044
rect 1727 6016 2153 6024
rect 2607 6016 2893 6024
rect 3027 6016 3073 6024
rect 3087 6016 3293 6024
rect 3667 6016 3973 6024
rect 4467 6016 4513 6024
rect 4527 6016 4873 6024
rect 5627 6016 5853 6024
rect 6167 6016 6433 6024
rect 907 5996 1052 6004
rect 1087 5996 1613 6004
rect 2647 5996 2813 6004
rect 4067 5996 4133 6004
rect 4707 5996 4852 6004
rect 4876 6004 4884 6012
rect 4876 5996 5573 6004
rect 5967 5996 6133 6004
rect 547 5976 913 5984
rect 1587 5976 1713 5984
rect 3127 5976 3513 5984
rect 3607 5976 3693 5984
rect 4187 5976 4493 5984
rect 4547 5976 4673 5984
rect 5747 5976 5873 5984
rect 6207 5976 6693 5984
rect 867 5956 1073 5964
rect 1127 5956 1193 5964
rect 1487 5956 1993 5964
rect 2007 5956 2253 5964
rect 5027 5956 5293 5964
rect 5607 5956 5653 5964
rect 6067 5956 6433 5964
rect 1687 5936 2384 5944
rect 2376 5924 2384 5936
rect 2587 5936 2753 5944
rect 4007 5936 4253 5944
rect 4307 5936 4364 5944
rect 2376 5916 2413 5924
rect 167 5897 253 5905
rect 787 5896 933 5904
rect 1627 5897 1673 5905
rect 1787 5896 1893 5904
rect 2047 5897 2092 5905
rect 2127 5897 2173 5905
rect 2196 5896 2373 5904
rect 607 5876 764 5884
rect 687 5856 733 5864
rect 756 5864 764 5876
rect 2196 5884 2204 5896
rect 2467 5896 2533 5904
rect 2687 5897 2713 5905
rect 2736 5896 2953 5904
rect 2736 5884 2744 5896
rect 3227 5896 3353 5904
rect 3396 5907 3404 5933
rect 3447 5916 3533 5924
rect 3367 5896 3384 5904
rect 3396 5896 3413 5907
rect 2147 5876 2204 5884
rect 2616 5876 2744 5884
rect 3376 5884 3384 5896
rect 3400 5893 3413 5896
rect 3467 5897 3493 5905
rect 3687 5896 3853 5904
rect 4107 5896 4173 5904
rect 3376 5876 3524 5884
rect 756 5856 813 5864
rect 827 5856 1073 5864
rect 1627 5856 1653 5864
rect 1747 5855 1773 5863
rect 1987 5856 2013 5864
rect 2067 5856 2113 5864
rect 2407 5855 2453 5863
rect 2616 5864 2624 5876
rect 2607 5856 2624 5864
rect 2787 5855 2813 5863
rect 2927 5855 2973 5863
rect 3067 5856 3193 5864
rect 3387 5856 3413 5864
rect 3516 5864 3524 5876
rect 4336 5867 4344 5894
rect 3516 5856 3653 5864
rect 3967 5856 4053 5864
rect 4067 5856 4193 5864
rect 4327 5856 4344 5867
rect 4356 5866 4364 5936
rect 4647 5936 4713 5944
rect 5207 5936 5253 5944
rect 6287 5936 6333 5944
rect 6347 5936 6573 5944
rect 4587 5916 4613 5924
rect 5027 5916 5313 5924
rect 5587 5916 6053 5924
rect 4427 5897 4473 5905
rect 4696 5884 4704 5894
rect 4847 5896 4953 5904
rect 5067 5897 5113 5905
rect 5136 5896 5213 5904
rect 5136 5884 5144 5896
rect 5367 5896 5393 5904
rect 5407 5896 5573 5904
rect 5396 5884 5404 5894
rect 5867 5897 5913 5905
rect 6127 5896 6173 5904
rect 4676 5880 4704 5884
rect 4673 5876 4704 5880
rect 5056 5876 5144 5884
rect 5256 5876 5404 5884
rect 5936 5876 5993 5884
rect 4673 5867 4687 5876
rect 4327 5853 4340 5856
rect 4407 5855 4453 5863
rect 4507 5856 4553 5864
rect 4727 5856 4753 5864
rect 5056 5864 5064 5876
rect 5047 5856 5064 5864
rect 5256 5864 5264 5876
rect 5247 5856 5264 5864
rect 5936 5864 5944 5876
rect 5347 5856 5944 5864
rect 6076 5864 6084 5894
rect 6226 5893 6227 5900
rect 6247 5896 6333 5904
rect 6487 5896 6513 5904
rect 6647 5897 6693 5905
rect 6213 5884 6227 5893
rect 6213 5880 6304 5884
rect 6216 5876 6304 5880
rect 6076 5856 6133 5864
rect 6296 5866 6304 5876
rect 6207 5855 6253 5863
rect 6467 5855 6553 5863
rect 6707 5856 6773 5864
rect 127 5835 193 5843
rect 4236 5836 4653 5844
rect 1007 5816 1093 5824
rect 1447 5816 2133 5824
rect 2187 5816 2353 5824
rect 2527 5816 2633 5824
rect 2847 5816 3133 5824
rect 3147 5816 4033 5824
rect 4236 5824 4244 5836
rect 4707 5836 4973 5844
rect 5527 5836 5973 5844
rect 6027 5836 6093 5844
rect 6107 5836 6353 5844
rect 6556 5844 6564 5852
rect 6556 5836 6813 5844
rect 4047 5816 4244 5824
rect 4256 5816 4312 5824
rect 2387 5796 2653 5804
rect 2667 5796 2733 5804
rect 3307 5796 3833 5804
rect 4256 5804 4264 5816
rect 4347 5816 4593 5824
rect 5167 5816 5253 5824
rect 5387 5816 5593 5824
rect 5727 5816 5873 5824
rect 6007 5816 6193 5824
rect 6587 5816 6653 5824
rect 4107 5796 4264 5804
rect 4287 5796 4753 5804
rect 4867 5796 5033 5804
rect 5087 5796 5333 5804
rect 5427 5796 5553 5804
rect 6347 5796 6373 5804
rect 6427 5796 6653 5804
rect 367 5776 673 5784
rect 687 5776 1033 5784
rect 1107 5776 1313 5784
rect 1327 5776 2293 5784
rect 2647 5776 3013 5784
rect 3247 5776 4153 5784
rect 4547 5776 4673 5784
rect 4947 5776 5013 5784
rect 5147 5776 5193 5784
rect 5207 5776 5292 5784
rect 5327 5776 5753 5784
rect 5767 5776 5853 5784
rect 5927 5776 6293 5784
rect 1967 5756 2373 5764
rect 3667 5756 4213 5764
rect 4267 5756 5144 5764
rect 1507 5736 1873 5744
rect 2507 5736 2573 5744
rect 2587 5736 2873 5744
rect 2927 5736 3573 5744
rect 3847 5736 4473 5744
rect 4627 5736 4693 5744
rect 4907 5736 5033 5744
rect 5047 5736 5113 5744
rect 5136 5744 5144 5756
rect 5347 5756 5633 5764
rect 6147 5756 6473 5764
rect 5136 5736 5773 5744
rect 6207 5736 6813 5744
rect 67 5716 193 5724
rect 207 5716 973 5724
rect 987 5716 1133 5724
rect 1927 5716 2093 5724
rect 2107 5716 2153 5724
rect 2307 5716 2633 5724
rect 3787 5716 4293 5724
rect 4307 5716 6093 5724
rect 1187 5696 1633 5704
rect 2247 5696 2673 5704
rect 3827 5696 4093 5704
rect 4147 5696 4193 5704
rect 4216 5696 5293 5704
rect 967 5676 1784 5684
rect 1776 5667 1784 5676
rect 1827 5676 2113 5684
rect 2967 5676 3593 5684
rect 4216 5684 4224 5696
rect 5607 5696 5793 5704
rect 6167 5696 6313 5704
rect 4127 5676 4224 5684
rect 4427 5676 5104 5684
rect 1787 5656 2233 5664
rect 2687 5656 3053 5664
rect 3967 5656 4313 5664
rect 4327 5656 4753 5664
rect 4967 5656 5053 5664
rect 5096 5664 5104 5676
rect 5507 5676 5953 5684
rect 6107 5676 6633 5684
rect 6647 5676 6713 5684
rect 5096 5656 5513 5664
rect 5567 5656 5613 5664
rect 5887 5656 5973 5664
rect 6387 5656 6573 5664
rect 1027 5636 1153 5644
rect 1427 5636 1913 5644
rect 2067 5636 2273 5644
rect 2287 5636 2484 5644
rect 367 5616 753 5624
rect 807 5616 993 5624
rect 1707 5616 1853 5624
rect 2476 5624 2484 5636
rect 2667 5636 2953 5644
rect 4207 5636 4793 5644
rect 4867 5636 5073 5644
rect 5167 5636 5373 5644
rect 6147 5636 6173 5644
rect 6807 5636 6893 5644
rect 2476 5616 2553 5624
rect 4187 5616 4413 5624
rect 4607 5616 4773 5624
rect 5487 5616 5513 5624
rect 6227 5616 6293 5624
rect 6587 5616 6753 5624
rect -24 5596 113 5604
rect 847 5596 913 5604
rect 1067 5597 1153 5605
rect 1267 5596 1293 5604
rect 1347 5596 1453 5604
rect 1467 5596 1593 5604
rect 1607 5596 1664 5604
rect 1656 5584 1664 5596
rect 1687 5597 1733 5605
rect 1847 5597 1913 5605
rect 1927 5596 2052 5604
rect 2087 5597 2133 5605
rect 2287 5596 2433 5604
rect 2516 5596 2733 5604
rect 2236 5584 2244 5594
rect 607 5576 884 5584
rect 1656 5576 2244 5584
rect 787 5555 833 5563
rect 876 5564 884 5576
rect 2516 5584 2524 5596
rect 2827 5597 2853 5605
rect 3067 5596 3093 5604
rect 3627 5597 3673 5605
rect 3747 5597 3813 5605
rect 3927 5596 4093 5604
rect 4107 5596 4193 5604
rect 2367 5576 2524 5584
rect 876 5556 893 5564
rect 907 5555 933 5563
rect 1007 5556 1033 5564
rect 1127 5555 1173 5563
rect 1287 5555 1333 5563
rect 1587 5555 1633 5563
rect 1767 5555 1813 5563
rect 1867 5556 1893 5564
rect 1947 5556 2093 5564
rect 2147 5556 2193 5564
rect 2307 5555 2493 5563
rect 2607 5555 2633 5563
rect 3087 5555 3133 5563
rect 3216 5564 3224 5594
rect 3576 5584 3584 5594
rect 4267 5596 4413 5604
rect 4467 5597 4493 5605
rect 4587 5596 4724 5604
rect 3576 5576 3624 5584
rect 3616 5567 3624 5576
rect 3187 5556 3224 5564
rect 3287 5556 3593 5564
rect 3616 5556 3633 5567
rect 3620 5553 3633 5556
rect 3687 5556 3753 5564
rect 3987 5556 4033 5564
rect 4047 5555 4073 5563
rect 4207 5555 4233 5563
rect 4287 5555 4313 5563
rect 4447 5556 4593 5564
rect 4716 5564 4724 5596
rect 4887 5596 4953 5604
rect 5127 5597 5193 5605
rect 5207 5596 5333 5604
rect 5387 5597 5433 5605
rect 5727 5596 5813 5604
rect 4793 5584 4807 5593
rect 4956 5584 4964 5594
rect 4793 5580 4924 5584
rect 4796 5576 4924 5580
rect 4956 5576 5073 5584
rect 4916 5566 4924 5576
rect 5287 5584 5300 5587
rect 5556 5584 5564 5594
rect 5827 5596 5873 5604
rect 6107 5597 6173 5605
rect 6356 5596 6373 5604
rect 5287 5573 5304 5584
rect 5556 5576 5644 5584
rect 4716 5556 4733 5564
rect 4787 5555 4813 5563
rect 4927 5555 5133 5563
rect 5156 5556 5173 5564
rect 1327 5536 1433 5544
rect 1547 5536 2193 5544
rect 2427 5536 2513 5544
rect 2887 5536 2953 5544
rect 4627 5536 4693 5544
rect 5156 5544 5164 5556
rect 5296 5564 5304 5573
rect 5296 5556 5393 5564
rect 5547 5556 5613 5564
rect 5007 5536 5164 5544
rect 5227 5536 5252 5544
rect 5287 5536 5513 5544
rect 5636 5544 5644 5576
rect 5787 5564 5800 5567
rect 5787 5553 5804 5564
rect 5636 5536 5693 5544
rect 5796 5544 5804 5553
rect 5907 5556 5973 5564
rect 5796 5536 5873 5544
rect 6056 5544 6064 5594
rect 6256 5567 6264 5594
rect 6356 5567 6364 5596
rect 6187 5556 6233 5564
rect 6256 5556 6273 5567
rect 6260 5553 6273 5556
rect 6416 5547 6424 5594
rect 6507 5596 6553 5604
rect 6596 5567 6604 5594
rect 6847 5597 6873 5605
rect 6696 5567 6704 5593
rect 6447 5556 6493 5564
rect 6596 5556 6613 5567
rect 6600 5553 6613 5556
rect 6776 5564 6784 5593
rect 6747 5556 6784 5564
rect 6916 5564 6924 5594
rect 6916 5556 6953 5564
rect 5947 5536 6064 5544
rect 6307 5536 6392 5544
rect 747 5516 853 5524
rect 907 5516 1233 5524
rect 1567 5516 1713 5524
rect 2067 5516 2173 5524
rect 2847 5516 3033 5524
rect 3047 5516 3113 5524
rect 3327 5516 3553 5524
rect 3727 5516 4033 5524
rect 4487 5516 5133 5524
rect 5187 5516 5293 5524
rect 5307 5516 5353 5524
rect 5647 5516 5733 5524
rect 5927 5516 6153 5524
rect 6487 5516 6573 5524
rect 6727 5516 6933 5524
rect 167 5496 513 5504
rect 887 5496 1333 5504
rect 2127 5496 2413 5504
rect 2647 5496 2673 5504
rect 2807 5496 2973 5504
rect 2987 5496 3124 5504
rect 267 5476 393 5484
rect 647 5476 1053 5484
rect 1167 5476 1293 5484
rect 1307 5476 1553 5484
rect 2207 5476 2353 5484
rect 2467 5476 3073 5484
rect 3116 5484 3124 5496
rect 3147 5496 3233 5504
rect 3647 5496 3984 5504
rect 3116 5476 3193 5484
rect 3207 5476 3233 5484
rect 3367 5476 3433 5484
rect 3447 5476 3613 5484
rect 3847 5476 3933 5484
rect 3976 5484 3984 5496
rect 4007 5496 4393 5504
rect 4687 5496 4813 5504
rect 4907 5496 4953 5504
rect 4967 5496 5113 5504
rect 5347 5496 5473 5504
rect 5687 5496 5713 5504
rect 5807 5496 6273 5504
rect 6287 5496 6413 5504
rect 6827 5496 6893 5504
rect 3976 5476 4093 5484
rect 4167 5476 4253 5484
rect 4587 5476 5213 5484
rect 5227 5476 5453 5484
rect 5667 5476 5773 5484
rect 5827 5476 6033 5484
rect 6667 5476 6933 5484
rect 247 5456 333 5464
rect 1587 5456 1873 5464
rect 1887 5456 2133 5464
rect 2387 5456 2413 5464
rect 4487 5456 4853 5464
rect 5367 5456 5433 5464
rect 5487 5456 5533 5464
rect 5547 5456 5633 5464
rect 5687 5456 5753 5464
rect 5856 5456 5933 5464
rect 5856 5447 5864 5456
rect 6207 5456 6353 5464
rect 787 5436 853 5444
rect 947 5436 1533 5444
rect 2687 5436 2713 5444
rect 3187 5436 3713 5444
rect 3807 5436 3893 5444
rect 3967 5436 4153 5444
rect 4207 5436 4293 5444
rect 4307 5436 4693 5444
rect 4947 5436 5053 5444
rect 5167 5436 5333 5444
rect 5467 5436 5604 5444
rect 487 5416 593 5424
rect 1047 5416 1393 5424
rect 2327 5416 2453 5424
rect 2747 5416 2893 5424
rect 3407 5416 3684 5424
rect 547 5396 753 5404
rect 2507 5396 2553 5404
rect 2607 5396 2653 5404
rect 3027 5396 3053 5404
rect 3676 5404 3684 5416
rect 4027 5416 4493 5424
rect 5087 5416 5273 5424
rect 5527 5416 5573 5424
rect 5596 5424 5604 5436
rect 5647 5436 5853 5444
rect 5967 5436 6033 5444
rect 6167 5436 6293 5444
rect 6387 5436 6453 5444
rect 5596 5416 5913 5424
rect 6407 5416 6453 5424
rect 6747 5416 6793 5424
rect 3676 5396 3753 5404
rect 4047 5396 4353 5404
rect 4567 5396 4624 5404
rect 707 5376 793 5384
rect 896 5376 933 5384
rect 40 5364 53 5367
rect 36 5353 53 5364
rect 387 5357 493 5365
rect 507 5356 873 5364
rect 16 5327 24 5353
rect 36 5326 44 5353
rect 547 5335 573 5343
rect 627 5335 693 5343
rect 747 5336 813 5344
rect 896 5327 904 5376
rect 987 5384 1000 5387
rect 987 5373 1004 5384
rect 1047 5380 1144 5384
rect 1047 5376 1147 5380
rect 996 5326 1004 5373
rect 1133 5367 1147 5376
rect 1447 5376 1533 5384
rect 1687 5377 1733 5385
rect 1967 5377 2013 5385
rect 2600 5384 2613 5387
rect 2376 5364 2384 5374
rect 2596 5373 2613 5384
rect 2787 5377 2853 5385
rect 3007 5377 3273 5385
rect 3347 5376 3373 5384
rect 3447 5376 3513 5384
rect 2596 5364 2604 5373
rect 2076 5356 2424 5364
rect 1767 5335 1853 5343
rect 2076 5344 2084 5356
rect 1867 5336 2084 5344
rect 2167 5336 2393 5344
rect 2416 5327 2424 5356
rect 2576 5356 2604 5364
rect 2576 5346 2584 5356
rect 3576 5347 3584 5374
rect 3627 5376 3773 5384
rect 3787 5376 3833 5384
rect 3887 5376 3904 5384
rect 3896 5347 3904 5376
rect 3987 5384 4000 5387
rect 3987 5373 4004 5384
rect 4107 5376 4184 5384
rect 2467 5335 2533 5343
rect 2667 5335 2713 5343
rect 2827 5336 2873 5344
rect 3127 5336 3253 5344
rect 3527 5335 3553 5343
rect 3576 5336 3593 5347
rect 3580 5333 3593 5336
rect 3647 5336 3693 5344
rect 3767 5336 3813 5344
rect 3996 5346 4004 5373
rect 4176 5364 4184 5376
rect 4547 5377 4593 5385
rect 4176 5356 4453 5364
rect 4616 5364 4624 5396
rect 4807 5396 5033 5404
rect 5787 5396 5853 5404
rect 6187 5396 6313 5404
rect 6567 5396 6633 5404
rect 4747 5377 4773 5385
rect 4987 5377 5073 5385
rect 5187 5377 5253 5385
rect 5367 5377 5413 5385
rect 5427 5376 5493 5384
rect 5727 5377 5753 5385
rect 5947 5376 6053 5384
rect 6127 5376 6164 5384
rect 4616 5356 4704 5364
rect 4047 5335 4113 5343
rect 4307 5335 4373 5343
rect 4607 5336 4673 5344
rect 4696 5344 4704 5356
rect 5653 5364 5667 5373
rect 5147 5360 5667 5364
rect 6156 5364 6164 5376
rect 6267 5376 6324 5384
rect 5147 5356 5664 5360
rect 6156 5356 6244 5364
rect 4696 5336 4853 5344
rect 4927 5336 4973 5344
rect 1607 5316 1713 5324
rect 2416 5316 2433 5327
rect 2420 5313 2433 5316
rect 2767 5316 3313 5324
rect 3407 5316 3473 5324
rect 4976 5324 4984 5333
rect 5067 5336 5233 5344
rect 5447 5336 5733 5344
rect 6236 5346 6244 5356
rect 6316 5347 6324 5376
rect 6427 5376 6533 5384
rect 6707 5376 6773 5384
rect 6827 5377 6853 5385
rect 6896 5347 6904 5373
rect 6956 5347 6964 5373
rect 5927 5336 5953 5344
rect 6407 5335 6433 5343
rect 6567 5335 6593 5343
rect 4976 5316 5273 5324
rect 5287 5316 5353 5324
rect 5687 5316 5793 5324
rect 6067 5316 6093 5324
rect 6167 5316 6333 5324
rect 6487 5316 6633 5324
rect 207 5296 473 5304
rect 1027 5296 1133 5304
rect 1747 5296 2073 5304
rect 2707 5296 3333 5304
rect 3347 5296 3533 5304
rect 4227 5296 4333 5304
rect 4347 5296 4493 5304
rect 4687 5296 4733 5304
rect 4807 5296 4853 5304
rect 5187 5296 5253 5304
rect 5547 5296 5653 5304
rect 5727 5296 5853 5304
rect 6027 5296 6293 5304
rect 27 5276 53 5284
rect 407 5276 433 5284
rect 967 5276 1053 5284
rect 2687 5276 2713 5284
rect 2727 5276 2753 5284
rect 3087 5276 3413 5284
rect 4927 5276 4953 5284
rect 4967 5276 5113 5284
rect 5307 5276 5333 5284
rect 5727 5276 5992 5284
rect 6027 5276 6224 5284
rect 1927 5256 2353 5264
rect 2447 5256 2993 5264
rect 3447 5256 3953 5264
rect 4856 5256 4904 5264
rect 1067 5236 1293 5244
rect 1436 5236 1493 5244
rect 787 5216 913 5224
rect 1436 5224 1444 5236
rect 1507 5236 2033 5244
rect 2427 5236 2673 5244
rect 2687 5236 2833 5244
rect 2947 5236 3013 5244
rect 3267 5236 3593 5244
rect 4856 5244 4864 5256
rect 3907 5236 4864 5244
rect 4896 5244 4904 5256
rect 5007 5256 5053 5264
rect 5247 5256 5373 5264
rect 5687 5256 6193 5264
rect 6216 5264 6224 5276
rect 6547 5276 6733 5284
rect 6216 5256 6373 5264
rect 4896 5236 5133 5244
rect 5667 5236 6133 5244
rect 6627 5236 6673 5244
rect 927 5216 1444 5224
rect 2867 5216 3053 5224
rect 4027 5216 4233 5224
rect 4247 5216 4653 5224
rect 4887 5216 5153 5224
rect 5207 5216 5313 5224
rect 5387 5216 5473 5224
rect 5627 5216 5733 5224
rect 6307 5216 6413 5224
rect 6527 5216 6593 5224
rect 6707 5216 6933 5224
rect 267 5196 333 5204
rect 827 5196 1073 5204
rect 1167 5196 1233 5204
rect 1467 5196 1973 5204
rect 3247 5196 3433 5204
rect 3747 5196 3793 5204
rect 5507 5196 5713 5204
rect 5767 5196 5873 5204
rect 5887 5196 5973 5204
rect 6147 5196 6473 5204
rect 2247 5176 2493 5184
rect 2987 5176 3333 5184
rect 3867 5176 3973 5184
rect 4187 5176 4213 5184
rect 4487 5176 4693 5184
rect 4767 5176 5313 5184
rect 5387 5176 5653 5184
rect 6007 5176 6253 5184
rect 6367 5176 6453 5184
rect 467 5156 1093 5164
rect 1647 5156 2533 5164
rect 2547 5156 3353 5164
rect 3827 5156 4053 5164
rect 4607 5156 4792 5164
rect 4827 5156 4993 5164
rect 5316 5164 5324 5173
rect 5316 5156 5813 5164
rect 5907 5156 6244 5164
rect 707 5136 873 5144
rect 2567 5136 2633 5144
rect 2747 5136 3153 5144
rect 3347 5136 3633 5144
rect 3947 5136 4073 5144
rect 4087 5136 4513 5144
rect 4527 5136 4573 5144
rect 5036 5136 5093 5144
rect 367 5116 613 5124
rect 627 5116 893 5124
rect 1567 5116 1813 5124
rect 1827 5116 1853 5124
rect 1867 5116 2213 5124
rect 2607 5116 3273 5124
rect 3787 5116 3873 5124
rect 4267 5116 4713 5124
rect 5036 5124 5044 5136
rect 5107 5136 5613 5144
rect 5847 5136 6093 5144
rect 6147 5136 6213 5144
rect 6236 5144 6244 5156
rect 6307 5156 6584 5164
rect 6236 5136 6432 5144
rect 6576 5144 6584 5156
rect 6647 5156 6893 5164
rect 6467 5136 6544 5144
rect 6576 5136 6913 5144
rect 4727 5116 5044 5124
rect 5067 5116 5433 5124
rect 5447 5116 5693 5124
rect 5707 5116 5773 5124
rect 5927 5116 5993 5124
rect 6267 5116 6493 5124
rect 6536 5124 6544 5136
rect 6536 5116 6853 5124
rect 6967 5124 6980 5127
rect 6967 5113 6984 5124
rect 747 5096 933 5104
rect 1307 5096 1433 5104
rect 2267 5096 2373 5104
rect 3587 5096 3653 5104
rect 4567 5096 4633 5104
rect 4907 5096 4933 5104
rect 5147 5096 5373 5104
rect 5827 5096 5893 5104
rect 5967 5096 6053 5104
rect 6107 5096 6133 5104
rect 6207 5096 6284 5104
rect -24 5076 113 5084
rect 187 5077 293 5085
rect 416 5076 553 5084
rect 416 5064 424 5076
rect 767 5077 813 5085
rect 1087 5076 1153 5084
rect 1347 5077 1373 5085
rect 1427 5076 1453 5084
rect 1467 5077 1553 5085
rect 1727 5077 1813 5085
rect 2327 5077 2353 5085
rect 2667 5076 2793 5084
rect 2847 5077 2893 5085
rect 3027 5076 3133 5084
rect 3227 5076 3473 5084
rect 3707 5077 3793 5085
rect 3847 5077 3893 5085
rect 3987 5076 4093 5084
rect 4167 5076 4313 5084
rect 376 5056 424 5064
rect 3933 5064 3947 5073
rect 3933 5060 4024 5064
rect 3936 5056 4024 5060
rect 376 5044 384 5056
rect 4016 5047 4024 5056
rect 4356 5064 4364 5074
rect 4267 5056 4364 5064
rect 4967 5076 5013 5084
rect 5407 5076 5513 5084
rect 5527 5077 5573 5085
rect 5627 5077 5692 5085
rect 5727 5076 5933 5084
rect 5956 5076 6173 5084
rect 4613 5064 4627 5073
rect 4613 5060 4684 5064
rect 4616 5056 4684 5060
rect 167 5036 384 5044
rect 667 5035 693 5043
rect 847 5035 893 5043
rect 1027 5035 1053 5043
rect 1107 5036 1133 5044
rect 1387 5036 1473 5044
rect 1567 5036 1633 5044
rect 1647 5036 1753 5044
rect 2387 5035 2433 5043
rect 2487 5035 2573 5043
rect 2827 5036 2872 5044
rect 2907 5036 2953 5044
rect 3167 5036 3313 5044
rect 3587 5035 3653 5043
rect 3747 5035 3773 5043
rect 4016 5036 4033 5047
rect 4020 5033 4033 5036
rect 4107 5035 4133 5043
rect 4187 5035 4233 5043
rect 4347 5036 4493 5044
rect 4587 5035 4633 5043
rect 4676 5044 4684 5056
rect 4676 5036 4813 5044
rect 4916 5044 4924 5073
rect 5047 5056 5184 5064
rect 4836 5036 4933 5044
rect 727 5016 993 5024
rect 2447 5016 2613 5024
rect 3907 5016 3953 5024
rect 4027 5016 4473 5024
rect 4836 5024 4844 5036
rect 5107 5036 5153 5044
rect 5176 5044 5184 5056
rect 5956 5064 5964 5076
rect 5847 5056 5964 5064
rect 6276 5064 6284 5096
rect 6887 5096 6953 5104
rect 6387 5076 6433 5084
rect 6507 5077 6553 5085
rect 6696 5064 6704 5074
rect 6276 5056 6364 5064
rect 5176 5036 5213 5044
rect 5287 5035 5313 5043
rect 5487 5036 5553 5044
rect 5647 5036 5753 5044
rect 5767 5036 5853 5044
rect 6356 5046 6364 5056
rect 6596 5056 6704 5064
rect 6596 5044 6604 5056
rect 6467 5036 6604 5044
rect 6716 5044 6724 5093
rect 6747 5077 6793 5085
rect 6716 5036 6753 5044
rect 4787 5016 4844 5024
rect 5596 5024 5604 5032
rect 5407 5016 5604 5024
rect 5807 5016 5844 5024
rect 247 4996 333 5004
rect 407 4996 653 5004
rect 787 4996 973 5004
rect 1247 4996 1313 5004
rect 2607 4996 2773 5004
rect 3507 4996 3853 5004
rect 3967 4996 3993 5004
rect 4007 4996 4253 5004
rect 4467 4996 5033 5004
rect 5227 4996 5813 5004
rect 5836 5004 5844 5016
rect 6627 5016 6712 5024
rect 6747 5016 6813 5024
rect 6976 5024 6984 5113
rect 6867 5016 6984 5024
rect 5836 4996 5913 5004
rect 5927 4996 6073 5004
rect 6187 4996 6213 5004
rect 6287 4996 6393 5004
rect 6407 4996 6573 5004
rect 6787 5004 6800 5007
rect 6787 4993 6804 5004
rect 1567 4976 1673 4984
rect 1687 4976 1913 4984
rect 2367 4976 2573 4984
rect 2587 4976 2993 4984
rect 3007 4976 3213 4984
rect 3387 4976 4013 4984
rect 4427 4976 4753 4984
rect 5347 4976 5493 4984
rect 5787 4976 5973 4984
rect 6207 4976 6453 4984
rect 6727 4976 6753 4984
rect 6796 4984 6804 4993
rect 6796 4976 6913 4984
rect 1027 4956 1273 4964
rect 1407 4956 1493 4964
rect 2307 4956 2453 4964
rect 2687 4956 2893 4964
rect 4036 4956 4693 4964
rect 1276 4944 1284 4953
rect 1276 4936 1473 4944
rect 1527 4936 1844 4944
rect 767 4916 1213 4924
rect 1836 4924 1844 4936
rect 2367 4936 2593 4944
rect 2896 4944 2904 4953
rect 4036 4947 4044 4956
rect 4827 4956 4913 4964
rect 5247 4956 5533 4964
rect 5627 4956 5673 4964
rect 5747 4956 5833 4964
rect 6007 4956 6073 4964
rect 6187 4956 6553 4964
rect 2896 4936 3453 4944
rect 3567 4936 3673 4944
rect 3827 4936 3873 4944
rect 4027 4936 4044 4947
rect 4027 4933 4040 4936
rect 4067 4936 4413 4944
rect 4487 4936 4933 4944
rect 5707 4936 6573 4944
rect 6587 4936 6833 4944
rect 1836 4916 1953 4924
rect 3707 4916 3813 4924
rect 3827 4916 4293 4924
rect 4447 4916 4853 4924
rect 4867 4916 4973 4924
rect 5127 4916 5273 4924
rect 5547 4916 5633 4924
rect 5767 4916 6173 4924
rect 6327 4916 6513 4924
rect 1467 4896 1753 4904
rect 2287 4896 2333 4904
rect 2747 4896 2913 4904
rect 3047 4896 3253 4904
rect 3787 4896 3913 4904
rect 4707 4896 5053 4904
rect 5667 4896 5693 4904
rect 5847 4896 5893 4904
rect 6027 4896 6053 4904
rect 6347 4896 6533 4904
rect 1887 4876 1913 4884
rect 2427 4876 2533 4884
rect 3327 4876 3404 4884
rect 287 4856 433 4864
rect 847 4857 893 4865
rect 916 4826 924 4873
rect 947 4857 973 4865
rect -24 4816 113 4824
rect 1096 4807 1104 4854
rect 1487 4857 1713 4865
rect 1847 4856 2033 4864
rect 2047 4856 2133 4864
rect 2267 4857 2313 4865
rect 2447 4856 2513 4864
rect 2607 4856 2813 4864
rect 2927 4857 2973 4865
rect 3027 4856 3073 4864
rect 1136 4824 1144 4853
rect 1327 4835 1453 4843
rect 2393 4844 2407 4853
rect 3116 4844 3124 4854
rect 3207 4856 3293 4864
rect 3307 4856 3353 4864
rect 2393 4840 2464 4844
rect 2396 4836 2464 4840
rect 3116 4836 3233 4844
rect 1136 4820 1184 4824
rect 1136 4816 1187 4820
rect 1173 4807 1187 4816
rect 1747 4815 1793 4823
rect 2207 4816 2333 4824
rect 2387 4815 2433 4823
rect 2456 4824 2464 4836
rect 2456 4816 2793 4824
rect 3087 4815 3133 4823
rect 3287 4815 3373 4823
rect 3396 4824 3404 4876
rect 3447 4876 3553 4884
rect 3627 4876 4113 4884
rect 4307 4876 4573 4884
rect 4687 4876 4813 4884
rect 4967 4876 5093 4884
rect 6507 4876 6533 4884
rect 6647 4876 6873 4884
rect 3487 4857 3513 4865
rect 3647 4856 4013 4864
rect 4136 4844 4144 4854
rect 4187 4856 4273 4864
rect 4296 4856 4313 4864
rect 4296 4844 4304 4856
rect 4507 4856 4633 4864
rect 4947 4856 5053 4864
rect 5167 4857 5233 4865
rect 5307 4856 5413 4864
rect 5427 4857 5493 4865
rect 5547 4856 5593 4864
rect 4136 4836 4304 4844
rect 3396 4816 3453 4824
rect 3727 4816 3793 4824
rect 3907 4815 3933 4823
rect 3987 4815 4033 4823
rect 4247 4816 4333 4824
rect 4487 4816 4733 4824
rect 4807 4815 4912 4823
rect 4947 4815 4973 4823
rect 5187 4815 5373 4823
rect 5656 4807 5664 4854
rect 6020 4864 6033 4867
rect 6016 4853 6033 4864
rect 6127 4856 6253 4864
rect 5740 4844 5753 4847
rect 5736 4833 5753 4844
rect 5736 4824 5744 4833
rect 5956 4827 5964 4853
rect 5687 4816 5744 4824
rect 6016 4824 6024 4853
rect 6007 4816 6024 4824
rect 6287 4815 6313 4823
rect 6476 4824 6484 4853
rect 6567 4856 6593 4864
rect 6367 4816 6484 4824
rect 6656 4824 6664 4854
rect 6707 4856 6893 4864
rect 6507 4816 6664 4824
rect 507 4796 613 4804
rect 667 4796 713 4804
rect 727 4796 753 4804
rect 1707 4796 1813 4804
rect 1827 4796 1893 4804
rect 2547 4796 2673 4804
rect 3367 4796 3613 4804
rect 4807 4796 5173 4804
rect 5287 4796 5353 4804
rect 5447 4796 5653 4804
rect 5787 4796 5813 4804
rect 6147 4796 6193 4804
rect 6647 4796 6773 4804
rect 6827 4796 6953 4804
rect 487 4776 633 4784
rect 647 4776 1153 4784
rect 2027 4776 2373 4784
rect 3107 4776 3193 4784
rect 3327 4776 3373 4784
rect 3387 4776 3673 4784
rect 4307 4776 4373 4784
rect 4427 4776 4513 4784
rect 4647 4776 5213 4784
rect 5367 4776 5444 4784
rect 87 4756 593 4764
rect 927 4756 973 4764
rect 1667 4756 2493 4764
rect 2507 4756 2813 4764
rect 4047 4756 4213 4764
rect 4227 4756 4933 4764
rect 4987 4756 5233 4764
rect 5247 4756 5413 4764
rect 5436 4764 5444 4776
rect 5867 4776 6113 4784
rect 5436 4756 5833 4764
rect 5887 4756 6073 4764
rect 6147 4756 6213 4764
rect 2267 4736 2593 4744
rect 2687 4736 2893 4744
rect 2907 4736 3273 4744
rect 3367 4736 3513 4744
rect 3527 4736 3724 4744
rect 707 4716 1073 4724
rect 1087 4716 1513 4724
rect 2807 4716 3033 4724
rect 3716 4724 3724 4736
rect 3747 4736 4093 4744
rect 4167 4736 4533 4744
rect 4667 4736 4853 4744
rect 4927 4736 5133 4744
rect 5187 4736 5213 4744
rect 5287 4736 5353 4744
rect 5787 4736 6053 4744
rect 3716 4716 3892 4724
rect 3927 4716 4353 4724
rect 4487 4716 4793 4724
rect 4947 4716 5513 4724
rect 5667 4716 6053 4724
rect 6247 4716 6413 4724
rect 6427 4716 6513 4724
rect 1127 4696 1413 4704
rect 1907 4696 2093 4704
rect 2347 4696 2453 4704
rect 2467 4696 2613 4704
rect 2627 4696 3453 4704
rect 3567 4696 3653 4704
rect 3667 4696 4373 4704
rect 4387 4696 4433 4704
rect 5136 4696 5333 4704
rect 47 4676 193 4684
rect 207 4676 313 4684
rect 2787 4676 2993 4684
rect 3067 4676 3413 4684
rect 3687 4676 4053 4684
rect 4400 4684 4413 4687
rect 4067 4676 4364 4684
rect 567 4656 1104 4664
rect 1096 4644 1104 4656
rect 2067 4656 2113 4664
rect 2127 4656 2173 4664
rect 2187 4656 3233 4664
rect 3927 4656 4333 4664
rect 4356 4664 4364 4676
rect 4396 4673 4413 4684
rect 4467 4676 4913 4684
rect 5136 4684 5144 4696
rect 5647 4696 6073 4704
rect 6127 4696 6333 4704
rect 4967 4676 5144 4684
rect 5307 4676 5433 4684
rect 5667 4676 6013 4684
rect 6067 4676 6373 4684
rect 4396 4664 4404 4673
rect 4356 4656 4404 4664
rect 4427 4656 5073 4664
rect 5147 4656 5253 4664
rect 5387 4656 5853 4664
rect 5987 4656 6233 4664
rect 1096 4636 1893 4644
rect 2847 4636 3373 4644
rect 3627 4636 3873 4644
rect 4267 4636 4513 4644
rect 5067 4636 5213 4644
rect 5387 4636 5433 4644
rect 5507 4636 5653 4644
rect 5727 4636 5813 4644
rect 5907 4636 6313 4644
rect 6447 4636 6833 4644
rect 2167 4616 2313 4624
rect 2527 4616 2753 4624
rect 2867 4616 3353 4624
rect 3527 4616 3793 4624
rect 4147 4616 4593 4624
rect 4787 4616 4873 4624
rect 4896 4616 5473 4624
rect 347 4596 404 4604
rect 233 4584 247 4593
rect 233 4580 384 4584
rect 236 4576 384 4580
rect -24 4556 113 4564
rect 353 4544 367 4553
rect 216 4540 367 4544
rect 216 4536 364 4540
rect 216 4526 224 4536
rect 167 4515 213 4523
rect 376 4504 384 4576
rect 396 4564 404 4596
rect 507 4596 913 4604
rect 1207 4596 1293 4604
rect 2827 4596 3053 4604
rect 3396 4596 3953 4604
rect 867 4576 953 4584
rect 1107 4576 1253 4584
rect 2287 4576 2353 4584
rect 2667 4576 2693 4584
rect 2707 4576 2853 4584
rect 2880 4584 2893 4587
rect 2876 4573 2893 4584
rect 3396 4584 3404 4596
rect 4007 4596 4213 4604
rect 4227 4596 4293 4604
rect 4447 4596 4633 4604
rect 4896 4604 4904 4616
rect 5607 4616 6344 4624
rect 6336 4607 6344 4616
rect 4707 4596 4904 4604
rect 4987 4596 5353 4604
rect 5527 4596 6052 4604
rect 6087 4596 6173 4604
rect 6336 4596 6353 4607
rect 6340 4593 6353 4596
rect 6607 4596 6673 4604
rect 3367 4576 3404 4584
rect 3427 4576 3553 4584
rect 3707 4576 3873 4584
rect 4107 4576 4173 4584
rect 4407 4576 4453 4584
rect 4467 4576 4653 4584
rect 4947 4576 5233 4584
rect 5256 4576 5333 4584
rect 396 4556 753 4564
rect 1027 4557 1073 4565
rect 1487 4556 1553 4564
rect 1807 4557 1833 4565
rect 1947 4556 2093 4564
rect 2107 4556 2153 4564
rect 2207 4556 2253 4564
rect 2387 4556 2453 4564
rect 2876 4564 2884 4573
rect 5256 4568 5264 4576
rect 5647 4576 5784 4584
rect 2856 4556 2884 4564
rect 547 4516 613 4524
rect 667 4515 733 4523
rect 787 4515 853 4523
rect 947 4516 1033 4524
rect 1107 4516 1173 4524
rect 1227 4516 1313 4524
rect 1707 4515 1812 4523
rect 1847 4515 1913 4523
rect 2127 4516 2233 4524
rect 2247 4515 2273 4523
rect 2347 4515 2433 4523
rect 2487 4516 2553 4524
rect 2567 4515 2593 4523
rect 2676 4524 2684 4553
rect 2676 4516 2793 4524
rect 2856 4524 2864 4556
rect 2907 4556 2973 4564
rect 2987 4556 3113 4564
rect 3167 4557 3213 4565
rect 3227 4556 3293 4564
rect 3667 4556 3764 4564
rect 3756 4544 3764 4556
rect 3847 4556 3864 4564
rect 3756 4536 3804 4544
rect 2847 4516 2864 4524
rect 3007 4515 3373 4523
rect 3487 4516 3533 4524
rect 3747 4515 3773 4523
rect 3796 4524 3804 4536
rect 3796 4516 3813 4524
rect 3856 4524 3864 4556
rect 4247 4557 4293 4565
rect 4536 4556 4693 4564
rect 4193 4544 4207 4553
rect 3907 4540 4207 4544
rect 3907 4536 4204 4540
rect 4156 4526 4164 4536
rect 3856 4516 4113 4524
rect 4327 4515 4393 4523
rect 4536 4524 4544 4556
rect 5027 4556 5073 4564
rect 5187 4556 5224 4564
rect 4940 4544 4953 4547
rect 4587 4536 4684 4544
rect 4527 4516 4544 4524
rect 4676 4526 4684 4536
rect 4936 4533 4953 4544
rect 5216 4544 5224 4556
rect 5527 4556 5653 4564
rect 5707 4557 5753 4565
rect 5776 4564 5784 4576
rect 5807 4576 5873 4584
rect 5776 4556 5993 4564
rect 6187 4557 6253 4565
rect 6367 4557 6453 4565
rect 5216 4536 5244 4544
rect 4607 4516 4633 4524
rect 4687 4516 4873 4524
rect 4936 4524 4944 4533
rect 4887 4516 4944 4524
rect 5127 4516 5193 4524
rect 5236 4524 5244 4536
rect 5416 4527 5424 4553
rect 5236 4516 5293 4524
rect 247 4496 384 4504
rect 907 4496 1073 4504
rect 2927 4496 2953 4504
rect 3067 4496 3313 4504
rect 3327 4496 3353 4504
rect 3967 4496 4013 4504
rect 607 4476 833 4484
rect 896 4484 904 4493
rect 4647 4496 4893 4504
rect 5287 4496 5433 4504
rect 847 4476 904 4484
rect 1147 4476 1193 4484
rect 1587 4476 1733 4484
rect 1747 4476 1773 4484
rect 1827 4476 1953 4484
rect 1967 4476 2893 4484
rect 3087 4476 3133 4484
rect 3407 4476 3453 4484
rect 3567 4476 3613 4484
rect 4387 4476 4453 4484
rect 4587 4476 4933 4484
rect 5307 4476 5373 4484
rect 5496 4486 5504 4553
rect 6036 4544 6044 4554
rect 6587 4556 6613 4564
rect 6747 4556 6773 4564
rect 6827 4557 6933 4565
rect 6036 4536 6113 4544
rect 6576 4527 6584 4553
rect 5547 4515 5593 4523
rect 5767 4516 5813 4524
rect 5907 4516 6053 4524
rect 6187 4516 6293 4524
rect 6387 4515 6433 4523
rect 6707 4516 6753 4524
rect 6776 4507 6784 4554
rect 5527 4496 5673 4504
rect 5947 4496 6012 4504
rect 6047 4496 6093 4504
rect 6147 4476 6193 4484
rect 6327 4476 6353 4484
rect 6447 4476 6553 4484
rect 3887 4456 4193 4464
rect 4487 4456 4533 4464
rect 4747 4456 4932 4464
rect 4967 4456 5033 4464
rect 5487 4456 5792 4464
rect 5827 4456 6213 4464
rect 6287 4456 6473 4464
rect 6707 4456 6793 4464
rect 267 4436 373 4444
rect 1007 4436 1153 4444
rect 2447 4436 2533 4444
rect 2547 4436 2973 4444
rect 3807 4436 4033 4444
rect 4167 4436 4293 4444
rect 4567 4436 4812 4444
rect 4847 4436 4893 4444
rect 5447 4436 5753 4444
rect 6127 4436 6233 4444
rect 6247 4436 6493 4444
rect 6507 4436 6633 4444
rect 2247 4416 3073 4424
rect 3307 4416 3433 4424
rect 3447 4416 3633 4424
rect 3707 4416 4013 4424
rect 4227 4416 4533 4424
rect 4816 4416 4953 4424
rect 247 4396 313 4404
rect 2087 4396 2133 4404
rect 2547 4396 3113 4404
rect 3127 4396 3193 4404
rect 3207 4396 3313 4404
rect 3327 4396 3933 4404
rect 4127 4396 4513 4404
rect 4816 4404 4824 4416
rect 5007 4416 5073 4424
rect 5327 4416 5893 4424
rect 5987 4416 6553 4424
rect 4567 4396 4824 4404
rect 4847 4396 4893 4404
rect 4947 4396 5173 4404
rect 5187 4396 5273 4404
rect 5527 4396 5573 4404
rect 5707 4396 5853 4404
rect 6127 4396 6233 4404
rect 6247 4396 6273 4404
rect 6327 4396 6513 4404
rect 6647 4396 6893 4404
rect 1207 4376 1273 4384
rect 1507 4376 1593 4384
rect 1967 4376 2193 4384
rect 2747 4376 2793 4384
rect 2947 4376 3033 4384
rect 3047 4376 3084 4384
rect 1647 4356 2324 4364
rect 167 4337 193 4345
rect 207 4336 273 4344
rect 287 4336 493 4344
rect 116 4324 124 4334
rect 587 4336 633 4344
rect 1167 4337 1233 4345
rect 1367 4337 1413 4345
rect 1487 4336 1524 4344
rect 116 4316 264 4324
rect -24 4296 13 4304
rect 256 4306 264 4316
rect 536 4316 993 4324
rect 536 4307 544 4316
rect 1067 4317 1433 4325
rect 87 4296 133 4304
rect 16 4284 24 4293
rect 267 4295 293 4303
rect 487 4296 533 4304
rect 1516 4306 1524 4336
rect 1687 4336 1704 4344
rect 827 4296 1213 4304
rect 1536 4304 1544 4334
rect 1696 4324 1704 4336
rect 1727 4336 1793 4344
rect 1816 4336 1853 4344
rect 1816 4324 1824 4336
rect 1867 4336 2033 4344
rect 2096 4336 2233 4344
rect 1696 4316 1824 4324
rect 1536 4296 1573 4304
rect 2096 4306 2104 4336
rect 2316 4344 2324 4356
rect 2687 4356 2713 4364
rect 3076 4364 3084 4376
rect 4107 4376 4204 4384
rect 3076 4356 3133 4364
rect 3147 4356 3373 4364
rect 3587 4356 3653 4364
rect 4196 4364 4204 4376
rect 4827 4376 4913 4384
rect 5027 4376 5093 4384
rect 6087 4376 6293 4384
rect 3976 4356 4184 4364
rect 4196 4356 4533 4364
rect 2287 4336 2304 4344
rect 2316 4336 2393 4344
rect 2296 4307 2304 4336
rect 2407 4336 2512 4344
rect 2547 4344 2560 4347
rect 2547 4333 2564 4344
rect 2587 4336 2653 4344
rect 2707 4344 2720 4347
rect 2707 4333 2724 4344
rect 2747 4336 2873 4344
rect 2927 4336 3053 4344
rect 3427 4336 3533 4344
rect 1747 4295 1773 4303
rect 1927 4295 1953 4303
rect 2187 4295 2213 4303
rect 2556 4306 2564 4333
rect 2716 4306 2724 4333
rect 3436 4307 3444 4336
rect 3596 4307 3604 4333
rect 3676 4307 3684 4333
rect 2607 4296 2713 4304
rect 3087 4295 3113 4303
rect 3167 4296 3193 4304
rect 3247 4296 3313 4304
rect 3507 4296 3553 4304
rect 3696 4304 3704 4334
rect 3787 4336 3853 4344
rect 3976 4347 3984 4356
rect 4067 4336 4144 4344
rect 3973 4324 3987 4333
rect 3916 4320 3987 4324
rect 3916 4316 3984 4320
rect 3696 4296 3833 4304
rect 3916 4304 3924 4316
rect 4136 4307 4144 4336
rect 3887 4296 3924 4304
rect 3947 4295 3993 4303
rect 4176 4306 4184 4356
rect 4867 4356 4913 4364
rect 4987 4356 5033 4364
rect 5600 4364 5613 4367
rect 5207 4356 5324 4364
rect 4247 4336 4273 4344
rect 4367 4337 4433 4345
rect 4567 4337 4593 4345
rect 4656 4336 4693 4344
rect 4656 4307 4664 4336
rect 4827 4344 4840 4347
rect 4827 4333 4844 4344
rect 4307 4295 4333 4303
rect 4447 4296 4533 4304
rect 4836 4306 4844 4333
rect 5047 4336 5293 4344
rect 4953 4324 4967 4333
rect 4953 4320 5024 4324
rect 4956 4316 5027 4320
rect 5013 4307 5027 4316
rect 5316 4306 5324 4356
rect 5596 4353 5613 4364
rect 5147 4295 5233 4303
rect 5436 4304 5444 4334
rect 5547 4336 5573 4344
rect 5436 4300 5484 4304
rect 5436 4296 5487 4300
rect 5473 4287 5487 4296
rect 16 4276 553 4284
rect 567 4276 593 4284
rect 1387 4276 1493 4284
rect 1707 4276 1873 4284
rect 2067 4276 2253 4284
rect 3047 4276 3133 4284
rect 4307 4276 4373 4284
rect 5307 4276 5393 4284
rect 247 4256 333 4264
rect 447 4256 573 4264
rect 587 4256 653 4264
rect 2707 4256 2753 4264
rect 2767 4256 2953 4264
rect 2967 4256 3293 4264
rect 3407 4256 3472 4264
rect 3507 4256 4313 4264
rect 4607 4256 4733 4264
rect 5087 4256 5193 4264
rect 5327 4256 5453 4264
rect 5596 4264 5604 4353
rect 5727 4356 5773 4364
rect 5927 4356 5953 4364
rect 5907 4336 5973 4344
rect 6067 4336 6093 4344
rect 6227 4344 6240 4347
rect 6227 4333 6244 4344
rect 6347 4336 6473 4344
rect 5616 4316 5873 4324
rect 5616 4306 5624 4316
rect 6236 4324 6244 4333
rect 6236 4316 6384 4324
rect 6107 4296 6173 4304
rect 6327 4296 6353 4304
rect 5927 4276 5993 4284
rect 6227 4276 6313 4284
rect 6376 4284 6384 4316
rect 6476 4307 6484 4334
rect 6476 4296 6493 4307
rect 6480 4293 6493 4296
rect 6376 4276 6433 4284
rect 6636 4284 6644 4334
rect 6607 4276 6644 4284
rect 5596 4256 5633 4264
rect 5947 4256 5973 4264
rect 1427 4236 1573 4244
rect 1587 4236 2073 4244
rect 2087 4236 2293 4244
rect 3007 4236 3053 4244
rect 3227 4236 3353 4244
rect 3667 4236 3713 4244
rect 3727 4236 4113 4244
rect 4227 4236 4713 4244
rect 4767 4236 5113 4244
rect 5247 4236 5753 4244
rect 6013 4244 6027 4253
rect 6287 4256 6373 4264
rect 6467 4256 6493 4264
rect 5947 4240 6027 4244
rect 5947 4236 6024 4240
rect 6047 4236 6153 4244
rect 6627 4236 6753 4244
rect 1087 4216 1213 4224
rect 1567 4216 2173 4224
rect 3947 4216 4073 4224
rect 4787 4216 5133 4224
rect 5936 4224 5944 4232
rect 5327 4216 5944 4224
rect 6447 4216 6493 4224
rect 547 4196 853 4204
rect 1447 4196 1693 4204
rect 3127 4196 3433 4204
rect 3487 4196 3773 4204
rect 3827 4196 4653 4204
rect 4676 4196 5153 4204
rect 887 4176 1064 4184
rect 727 4156 813 4164
rect 1056 4164 1064 4176
rect 2227 4176 2493 4184
rect 3427 4176 3453 4184
rect 3967 4176 4073 4184
rect 4676 4184 4684 4196
rect 5207 4196 5673 4204
rect 6087 4196 6113 4204
rect 6247 4196 6373 4204
rect 6427 4196 6753 4204
rect 4547 4176 4684 4184
rect 4696 4176 4793 4184
rect 1056 4156 1153 4164
rect 2187 4156 2633 4164
rect 3236 4156 4093 4164
rect 847 4136 1013 4144
rect 2527 4136 2933 4144
rect 3236 4144 3244 4156
rect 4207 4156 4304 4164
rect 3207 4136 3244 4144
rect 3647 4136 4273 4144
rect 4296 4144 4304 4156
rect 4407 4156 4513 4164
rect 4696 4164 4704 4176
rect 4867 4176 5353 4184
rect 5647 4176 5833 4184
rect 5967 4176 6193 4184
rect 6207 4176 6333 4184
rect 4527 4156 4704 4164
rect 4747 4156 5653 4164
rect 5667 4156 5693 4164
rect 5707 4156 5893 4164
rect 5907 4156 6133 4164
rect 4296 4136 4813 4144
rect 5007 4136 5053 4144
rect 5107 4136 5273 4144
rect 5367 4136 5633 4144
rect 5916 4136 6073 4144
rect 807 4116 913 4124
rect 927 4116 953 4124
rect 1607 4116 1673 4124
rect 1687 4116 1753 4124
rect 3087 4116 3533 4124
rect 3927 4116 4093 4124
rect 4327 4116 4753 4124
rect 5127 4116 5173 4124
rect 5367 4116 5713 4124
rect 5916 4124 5924 4136
rect 6087 4136 6304 4144
rect 5767 4116 5924 4124
rect 6027 4116 6213 4124
rect 6296 4124 6304 4136
rect 6507 4136 6793 4144
rect 6927 4136 6953 4144
rect 6296 4116 6473 4124
rect 187 4096 213 4104
rect 227 4096 1353 4104
rect 2327 4096 2533 4104
rect 2547 4096 2633 4104
rect 2687 4096 2713 4104
rect 2727 4096 2773 4104
rect 3707 4096 3793 4104
rect 4147 4096 4213 4104
rect 4447 4096 4664 4104
rect 4656 4087 4664 4096
rect 4707 4096 4913 4104
rect 4927 4096 5373 4104
rect 6507 4096 6533 4104
rect 827 4076 944 4084
rect 447 4056 733 4064
rect 936 4064 944 4076
rect 967 4076 1113 4084
rect 1127 4076 1193 4084
rect 1556 4076 1613 4084
rect 936 4056 1073 4064
rect 1307 4056 1433 4064
rect -24 4036 113 4044
rect 266 4033 267 4040
rect 287 4036 424 4044
rect 253 4024 267 4033
rect 253 4020 393 4024
rect 255 4016 393 4020
rect 247 3996 293 4004
rect 416 3984 424 4036
rect 1067 4037 1093 4045
rect 1487 4037 1513 4045
rect 1556 4047 1564 4076
rect 1907 4076 1993 4084
rect 2567 4076 2653 4084
rect 2987 4076 3293 4084
rect 3787 4076 3973 4084
rect 4667 4076 4904 4084
rect 2527 4056 2673 4064
rect 2747 4056 2793 4064
rect 2927 4056 3133 4064
rect 3347 4056 3372 4064
rect 3407 4056 3593 4064
rect 3613 4064 3627 4073
rect 3613 4060 3873 4064
rect 3616 4056 3873 4060
rect 3887 4056 4133 4064
rect 4287 4056 4353 4064
rect 4467 4056 4573 4064
rect 4587 4056 4833 4064
rect 4896 4064 4904 4076
rect 5027 4076 5133 4084
rect 5267 4076 5513 4084
rect 5587 4076 5613 4084
rect 5747 4076 5793 4084
rect 6327 4076 6393 4084
rect 6447 4076 6553 4084
rect 6847 4076 6913 4084
rect 4896 4056 5213 4064
rect 5287 4056 5553 4064
rect 5687 4056 5884 4064
rect 547 4017 673 4025
rect 727 4015 853 4023
rect 947 3996 1033 4004
rect 1636 4006 1644 4053
rect 1807 4036 1873 4044
rect 1887 4037 1933 4045
rect 1987 4036 2033 4044
rect 2427 4037 2453 4045
rect 3007 4037 3033 4045
rect 3456 4036 3753 4044
rect 1367 3996 1413 4004
rect 1567 3995 1593 4003
rect 1727 3995 1773 4003
rect 2087 3995 2153 4003
rect 2347 3995 2393 4003
rect 2507 3995 2533 4003
rect 2827 3995 2893 4003
rect 2947 3995 2973 4003
rect 3456 4006 3464 4036
rect 4027 4036 4433 4044
rect 4487 4036 4544 4044
rect 4067 4016 4373 4024
rect 4536 4007 4544 4036
rect 4887 4036 4953 4044
rect 5007 4036 5113 4044
rect 5347 4037 5433 4045
rect 5507 4036 5533 4044
rect 5556 4044 5564 4053
rect 5556 4036 5573 4044
rect 5876 4044 5884 4056
rect 6056 4056 6093 4064
rect 5876 4036 5953 4044
rect 5256 4016 5473 4024
rect 3087 3996 3133 4004
rect 3247 3995 3313 4003
rect 3507 3995 3533 4003
rect 4107 3996 4153 4004
rect 4287 3995 4353 4003
rect 5256 4006 5264 4016
rect 5527 4024 5540 4027
rect 5527 4013 5544 4024
rect 4607 3995 4633 4003
rect 4827 3995 4853 4003
rect 5027 3995 5073 4003
rect 5347 3996 5453 4004
rect 5536 4004 5544 4013
rect 5536 3996 5693 4004
rect 5716 4004 5724 4034
rect 5756 4024 5764 4034
rect 5756 4016 5784 4024
rect 5776 4004 5784 4016
rect 5716 4000 5764 4004
rect 5716 3996 5767 4000
rect 5776 3996 5873 4004
rect 416 3976 433 3984
rect 447 3976 773 3984
rect 1287 3976 1333 3984
rect 1967 3976 2113 3984
rect 2396 3984 2404 3992
rect 5753 3987 5767 3996
rect 5927 3996 6013 4004
rect 6056 4006 6064 4056
rect 6507 4056 6544 4064
rect 6127 4036 6173 4044
rect 6116 4004 6124 4034
rect 6216 4036 6233 4044
rect 6216 4024 6224 4036
rect 6316 4036 6373 4044
rect 6187 4016 6224 4024
rect 6316 4007 6324 4036
rect 6436 4007 6444 4033
rect 6116 3996 6213 4004
rect 6307 3996 6324 4007
rect 6307 3993 6320 3996
rect 6367 3996 6393 4004
rect 6536 4006 6544 4056
rect 6687 4056 6793 4064
rect 6567 4036 6593 4044
rect 6896 4007 6904 4033
rect 6667 3995 6693 4003
rect 6807 3996 6833 4004
rect 2396 3976 3993 3984
rect 4507 3976 4564 3984
rect 207 3956 353 3964
rect 1227 3956 1473 3964
rect 3147 3956 3293 3964
rect 3307 3956 3793 3964
rect 4467 3956 4513 3964
rect 4556 3964 4564 3976
rect 4727 3976 4793 3984
rect 4807 3976 4893 3984
rect 5587 3976 5613 3984
rect 5947 3976 5973 3984
rect 6147 3976 6173 3984
rect 4556 3956 4893 3964
rect 5647 3956 5733 3964
rect 5787 3956 5953 3964
rect 6127 3956 6253 3964
rect 6487 3956 6573 3964
rect 476 3940 753 3944
rect 473 3936 753 3940
rect 473 3927 487 3936
rect 767 3936 793 3944
rect 1087 3936 1153 3944
rect 1567 3936 2293 3944
rect 2807 3936 2913 3944
rect 3007 3936 3693 3944
rect 3967 3936 4493 3944
rect 4547 3936 4792 3944
rect 4827 3936 4904 3944
rect 27 3916 413 3924
rect 547 3916 673 3924
rect 867 3916 1373 3924
rect 3387 3916 3884 3924
rect 1127 3896 1193 3904
rect 1827 3896 2413 3904
rect 2867 3896 3833 3904
rect 3876 3904 3884 3916
rect 4027 3916 4253 3924
rect 4387 3916 4753 3924
rect 4896 3924 4904 3936
rect 5167 3936 5313 3944
rect 6287 3936 6393 3944
rect 6527 3936 6553 3944
rect 6667 3936 6893 3944
rect 4896 3916 4993 3924
rect 5147 3916 5253 3924
rect 5547 3916 5673 3924
rect 6007 3916 6133 3924
rect 6187 3916 6253 3924
rect 3876 3896 4493 3904
rect 4507 3896 5173 3904
rect 5187 3896 5333 3904
rect 5347 3896 5513 3904
rect 5567 3896 5713 3904
rect 5827 3896 5973 3904
rect 6387 3896 6513 3904
rect 6767 3896 6953 3904
rect 407 3876 613 3884
rect 987 3876 1053 3884
rect 1067 3876 1084 3884
rect 1076 3864 1084 3876
rect 1216 3876 1493 3884
rect 1216 3864 1224 3876
rect 1647 3876 2213 3884
rect 2667 3876 3033 3884
rect 3047 3876 3433 3884
rect 3867 3876 3913 3884
rect 3927 3876 4053 3884
rect 4067 3876 4233 3884
rect 4247 3876 4404 3884
rect 1076 3856 1224 3864
rect 2467 3856 2673 3864
rect 2827 3856 2944 3864
rect 347 3836 393 3844
rect 927 3836 993 3844
rect 1827 3836 1853 3844
rect 2936 3844 2944 3856
rect 3567 3856 3633 3864
rect 4396 3864 4404 3876
rect 4607 3876 4824 3884
rect 4396 3856 4453 3864
rect 4816 3864 4824 3876
rect 4867 3876 5073 3884
rect 5627 3876 5793 3884
rect 5976 3876 6113 3884
rect 4816 3856 5033 3864
rect 5427 3856 5473 3864
rect 5976 3864 5984 3876
rect 6187 3876 6233 3884
rect 6287 3876 6353 3884
rect 6647 3876 6673 3884
rect 6747 3876 6933 3884
rect 5787 3856 5984 3864
rect 6007 3856 6053 3864
rect 6447 3856 6533 3864
rect 6587 3856 6633 3864
rect 6876 3856 6913 3864
rect 2936 3836 3033 3844
rect 3267 3836 3353 3844
rect 3427 3836 3493 3844
rect 4087 3836 4533 3844
rect 4647 3836 4753 3844
rect 4807 3836 5153 3844
rect 5440 3844 5453 3847
rect 5436 3833 5453 3844
rect 5827 3836 5913 3844
rect 6107 3836 6213 3844
rect 147 3816 253 3824
rect 267 3817 313 3825
rect 667 3817 713 3825
rect 1087 3816 1204 3824
rect 796 3787 804 3814
rect 1087 3796 1172 3804
rect 1196 3806 1204 3816
rect 1407 3816 1573 3824
rect 1887 3817 1953 3825
rect 2287 3816 2352 3824
rect 2387 3817 2493 3825
rect 2627 3816 2713 3824
rect 2736 3816 2873 3824
rect 1347 3796 1504 3804
rect 167 3775 193 3783
rect 207 3776 293 3784
rect 347 3776 604 3784
rect 267 3756 333 3764
rect 596 3764 604 3776
rect 787 3776 804 3787
rect 787 3773 800 3776
rect 867 3776 973 3784
rect 1496 3784 1504 3796
rect 2736 3804 2744 3816
rect 2927 3817 2953 3825
rect 3087 3816 3233 3824
rect 3407 3816 3473 3824
rect 3607 3816 3673 3824
rect 3687 3816 3733 3824
rect 4107 3816 4284 3824
rect 2187 3796 2744 3804
rect 3187 3796 3333 3804
rect 3776 3804 3784 3814
rect 3527 3796 3784 3804
rect 1496 3776 1553 3784
rect 1687 3775 1753 3783
rect 1807 3776 1933 3784
rect 1947 3776 2053 3784
rect 2227 3775 2293 3783
rect 2367 3775 2473 3783
rect 2907 3776 2924 3784
rect 596 3756 633 3764
rect 747 3755 1033 3763
rect 2916 3764 2924 3776
rect 3107 3775 3133 3783
rect 3427 3776 3493 3784
rect 4276 3786 4284 3816
rect 4307 3817 4373 3825
rect 4627 3824 4640 3827
rect 4627 3813 4644 3824
rect 4667 3816 4733 3824
rect 4847 3817 4913 3825
rect 5187 3816 5233 3824
rect 5436 3824 5444 3833
rect 5276 3816 5444 3824
rect 3647 3776 3713 3784
rect 3807 3776 4113 3784
rect 4636 3786 4644 3813
rect 5276 3804 5284 3816
rect 5807 3816 5833 3824
rect 5896 3816 5953 3824
rect 5216 3800 5284 3804
rect 5213 3796 5284 3800
rect 5696 3796 5773 3804
rect 5213 3787 5227 3796
rect 4387 3776 4473 3784
rect 4527 3775 4553 3783
rect 4687 3776 4813 3784
rect 4887 3776 4933 3784
rect 4947 3775 4993 3783
rect 5107 3775 5153 3783
rect 5427 3775 5453 3783
rect 2916 3760 3084 3764
rect 2916 3756 3087 3760
rect 3073 3747 3087 3756
rect 3207 3756 3393 3764
rect 3416 3756 3573 3764
rect 727 3736 853 3744
rect 1487 3736 2033 3744
rect 2227 3736 2433 3744
rect 3416 3744 3424 3756
rect 4367 3756 4453 3764
rect 4767 3756 4833 3764
rect 5187 3756 5393 3764
rect 5696 3764 5704 3796
rect 5896 3786 5904 3816
rect 5967 3816 6053 3824
rect 6173 3826 6187 3836
rect 6367 3836 6433 3844
rect 6487 3836 6624 3844
rect 6387 3816 6424 3824
rect 6293 3804 6307 3813
rect 6293 3800 6384 3804
rect 6296 3796 6387 3800
rect 6373 3787 6387 3796
rect 6147 3776 6253 3784
rect 6416 3786 6424 3816
rect 6456 3816 6593 3824
rect 6456 3786 6464 3816
rect 6616 3824 6624 3836
rect 6616 3816 6773 3824
rect 6876 3827 6884 3856
rect 6776 3804 6784 3814
rect 6867 3816 6884 3827
rect 6867 3813 6880 3816
rect 6776 3800 6804 3804
rect 6776 3796 6807 3800
rect 6793 3787 6807 3796
rect 6507 3775 6573 3783
rect 6627 3776 6693 3784
rect 6707 3776 6753 3784
rect 6916 3784 6924 3814
rect 6936 3787 6944 3813
rect 6887 3776 6924 3784
rect 5407 3756 5704 3764
rect 5747 3756 5813 3764
rect 6107 3756 6213 3764
rect 6467 3756 6533 3764
rect 3347 3736 3424 3744
rect 3447 3736 3853 3744
rect 4347 3736 4513 3744
rect 4607 3736 4633 3744
rect 4927 3736 5033 3744
rect 5047 3736 5213 3744
rect 5787 3736 5993 3744
rect 6236 3736 6304 3744
rect 6236 3727 6244 3736
rect 67 3716 353 3724
rect 927 3716 1453 3724
rect 1527 3716 1933 3724
rect 2267 3716 2293 3724
rect 2427 3716 2913 3724
rect 2967 3716 3053 3724
rect 3247 3716 4113 3724
rect 4327 3716 4733 3724
rect 4967 3716 5192 3724
rect 5227 3716 5552 3724
rect 5587 3716 5673 3724
rect 5767 3716 5953 3724
rect 6007 3716 6113 3724
rect 6227 3716 6244 3727
rect 6296 3724 6304 3736
rect 6367 3736 6433 3744
rect 6296 3716 6413 3724
rect 6227 3713 6240 3716
rect 6527 3716 6753 3724
rect 787 3696 1473 3704
rect 2367 3696 2693 3704
rect 3087 3696 3213 3704
rect 3687 3696 4073 3704
rect 4087 3696 4433 3704
rect 4587 3696 4673 3704
rect 5087 3696 5773 3704
rect 5827 3696 6093 3704
rect 6287 3696 6473 3704
rect 427 3676 544 3684
rect 536 3664 544 3676
rect 1367 3676 1633 3684
rect 1867 3676 2373 3684
rect 3667 3676 3873 3684
rect 4467 3676 4713 3684
rect 5167 3676 5233 3684
rect 5667 3676 6044 3684
rect 536 3656 853 3664
rect 1987 3656 2173 3664
rect 2196 3656 2633 3664
rect 127 3636 433 3644
rect 447 3636 473 3644
rect 527 3636 1293 3644
rect 2196 3644 2204 3656
rect 2787 3656 2913 3664
rect 3227 3656 3473 3664
rect 3487 3656 3613 3664
rect 3627 3656 3933 3664
rect 3947 3656 4333 3664
rect 4467 3656 4693 3664
rect 4747 3656 4853 3664
rect 5336 3656 5733 3664
rect 5336 3647 5344 3656
rect 5867 3656 5993 3664
rect 6036 3664 6044 3676
rect 6147 3676 6172 3684
rect 6207 3676 6293 3684
rect 6487 3676 6653 3684
rect 6036 3656 6093 3664
rect 6107 3656 6313 3664
rect 6387 3656 6413 3664
rect 6427 3656 6513 3664
rect 6687 3656 6833 3664
rect 1747 3636 2204 3644
rect 2527 3636 3293 3644
rect 3316 3636 3753 3644
rect 467 3616 653 3624
rect 1727 3616 2713 3624
rect 2867 3616 2933 3624
rect 3316 3624 3324 3636
rect 4187 3636 4253 3644
rect 4447 3636 5333 3644
rect 5567 3636 5693 3644
rect 6567 3636 6893 3644
rect 2947 3616 3324 3624
rect 3487 3616 3633 3624
rect 3847 3616 3913 3624
rect 4087 3616 4413 3624
rect 4527 3616 4653 3624
rect 4707 3616 4733 3624
rect 4776 3616 5173 3624
rect 507 3596 593 3604
rect 707 3596 753 3604
rect 847 3596 893 3604
rect 1307 3596 1393 3604
rect 2676 3596 3053 3604
rect 2676 3587 2684 3596
rect 3067 3596 3513 3604
rect 4127 3596 4413 3604
rect 4776 3604 4784 3616
rect 5516 3616 5913 3624
rect 4727 3596 4784 3604
rect 5516 3604 5524 3616
rect 6227 3616 6953 3624
rect 5147 3596 5524 3604
rect 5587 3596 5633 3604
rect 5647 3596 5813 3604
rect 5967 3596 6104 3604
rect 176 3580 673 3584
rect 173 3576 673 3580
rect 173 3567 187 3576
rect 1107 3576 1153 3584
rect 1167 3576 1393 3584
rect 1767 3576 2133 3584
rect 2627 3576 2673 3584
rect 4207 3576 4473 3584
rect 4787 3576 4893 3584
rect 4907 3576 5033 3584
rect 5427 3576 5533 3584
rect 5547 3576 5853 3584
rect 6096 3584 6104 3596
rect 6127 3596 6153 3604
rect 6096 3576 6213 3584
rect 6267 3576 6373 3584
rect 367 3556 493 3564
rect 767 3556 873 3564
rect 887 3556 913 3564
rect 2827 3556 2893 3564
rect 3267 3556 3353 3564
rect 4387 3556 4533 3564
rect 4807 3556 4872 3564
rect 4907 3556 5133 3564
rect 5567 3556 5673 3564
rect 5687 3556 5813 3564
rect 5827 3556 5933 3564
rect 6027 3556 6073 3564
rect 47 3536 93 3544
rect 1607 3536 1713 3544
rect 1867 3536 1893 3544
rect 2007 3536 2104 3544
rect 647 3516 773 3524
rect 967 3517 993 3525
rect 1107 3516 1173 3524
rect 1187 3516 1253 3524
rect 1347 3517 1433 3525
rect 1547 3516 1673 3524
rect 2096 3524 2104 3536
rect 2267 3536 2433 3544
rect 2447 3536 2633 3544
rect 2747 3536 2793 3544
rect 2807 3536 3033 3544
rect 3087 3536 3113 3544
rect 3127 3536 3173 3544
rect 3327 3536 3364 3544
rect 2096 3516 2113 3524
rect 2507 3516 2553 3524
rect 2847 3516 2993 3524
rect 193 3504 207 3513
rect 193 3500 353 3504
rect 196 3496 353 3500
rect 2176 3496 2213 3504
rect 87 3476 453 3484
rect 547 3476 573 3484
rect 687 3476 893 3484
rect 1387 3476 1493 3484
rect 1827 3476 1873 3484
rect 2176 3484 2184 3496
rect 2107 3476 2184 3484
rect 2727 3476 2813 3484
rect 2867 3475 2893 3483
rect 2947 3475 2973 3483
rect 3047 3476 3113 3484
rect 3136 3467 3144 3514
rect 3167 3475 3192 3483
rect 3227 3476 3273 3484
rect 3356 3486 3364 3536
rect 3596 3536 3653 3544
rect 3456 3500 3573 3504
rect 3453 3496 3573 3500
rect 3453 3487 3467 3496
rect 3596 3504 3604 3536
rect 3987 3537 4013 3545
rect 4507 3536 4553 3544
rect 4756 3536 4793 3544
rect 4087 3516 4213 3524
rect 4393 3524 4407 3533
rect 4287 3516 4624 3524
rect 3587 3496 3664 3504
rect 3656 3484 3664 3496
rect 3687 3497 3813 3505
rect 4616 3507 4624 3516
rect 4707 3516 4733 3524
rect 4756 3524 4764 3536
rect 5067 3536 5153 3544
rect 5507 3536 5613 3544
rect 5627 3536 5793 3544
rect 5987 3536 6133 3544
rect 6280 3544 6293 3547
rect 6276 3533 6293 3544
rect 6540 3544 6553 3547
rect 6347 3540 6484 3544
rect 6347 3536 6487 3540
rect 4747 3516 4764 3524
rect 4867 3517 4913 3525
rect 4927 3516 5193 3524
rect 5247 3516 5293 3524
rect 5387 3516 5413 3524
rect 5516 3516 5552 3524
rect 3947 3496 4053 3504
rect 4616 3496 4633 3507
rect 4620 3493 4633 3496
rect 4813 3504 4827 3513
rect 4813 3500 5073 3504
rect 4816 3496 5073 3500
rect 5267 3496 5433 3504
rect 3656 3476 3924 3484
rect 767 3456 1013 3464
rect 1076 3456 1333 3464
rect 1076 3447 1084 3456
rect 2207 3456 2273 3464
rect 2667 3456 2753 3464
rect 407 3436 433 3444
rect 447 3436 833 3444
rect 847 3436 1073 3444
rect 1336 3444 1344 3453
rect 3227 3456 3313 3464
rect 3427 3456 3493 3464
rect 3916 3464 3924 3476
rect 4087 3476 4113 3484
rect 5516 3486 5524 3516
rect 5587 3516 5633 3524
rect 5833 3524 5847 3533
rect 5816 3520 5847 3524
rect 5816 3516 5844 3520
rect 5816 3504 5824 3516
rect 6027 3517 6073 3525
rect 5696 3496 5824 3504
rect 6276 3504 6284 3533
rect 6473 3527 6487 3536
rect 6536 3533 6553 3544
rect 6536 3527 6544 3533
rect 6307 3516 6333 3524
rect 6400 3524 6413 3527
rect 6396 3513 6413 3524
rect 6616 3516 6673 3524
rect 6276 3496 6304 3504
rect 4667 3475 4713 3483
rect 4907 3475 5013 3483
rect 5307 3475 5353 3483
rect 5696 3484 5704 3496
rect 5567 3476 5704 3484
rect 5727 3476 5833 3484
rect 5887 3475 5993 3483
rect 6087 3476 6153 3484
rect 6207 3475 6233 3483
rect 3916 3456 4053 3464
rect 4067 3456 4393 3464
rect 4487 3456 4653 3464
rect 5047 3456 5233 3464
rect 5327 3456 5473 3464
rect 6296 3464 6304 3496
rect 6396 3486 6404 3513
rect 6616 3487 6624 3516
rect 6946 3513 6947 3520
rect 6967 3516 7004 3524
rect 6327 3476 6353 3484
rect 6607 3476 6624 3487
rect 6607 3473 6620 3476
rect 6856 3484 6864 3513
rect 6933 3507 6947 3513
rect 6933 3506 6960 3507
rect 6933 3500 6953 3506
rect 6936 3496 6953 3500
rect 6940 3493 6953 3496
rect 6747 3476 6893 3484
rect 6296 3456 6373 3464
rect 6767 3456 6833 3464
rect 1336 3436 1733 3444
rect 2187 3436 2473 3444
rect 3607 3436 4273 3444
rect 4367 3436 4453 3444
rect 4607 3436 4753 3444
rect 5407 3436 5553 3444
rect 5947 3436 6153 3444
rect 6447 3436 6693 3444
rect 6747 3436 6953 3444
rect 487 3416 753 3424
rect 947 3416 1413 3424
rect 1967 3416 2733 3424
rect 3007 3416 3273 3424
rect 3547 3416 4072 3424
rect 4107 3416 4153 3424
rect 4307 3416 4553 3424
rect 4576 3416 4733 3424
rect 1007 3396 1233 3404
rect 1487 3396 1553 3404
rect 1567 3396 1813 3404
rect 2147 3396 2213 3404
rect 2227 3396 2313 3404
rect 3367 3396 3433 3404
rect 4576 3404 4584 3416
rect 5247 3416 5333 3424
rect 5627 3416 5673 3424
rect 5847 3416 5893 3424
rect 6107 3416 6213 3424
rect 6307 3416 6513 3424
rect 6667 3416 6773 3424
rect 4267 3396 4584 3404
rect 4596 3396 4813 3404
rect 427 3376 653 3384
rect 2867 3376 3053 3384
rect 3927 3376 3993 3384
rect 4367 3376 4473 3384
rect 4596 3384 4604 3396
rect 4827 3396 4973 3404
rect 5287 3396 5393 3404
rect 5627 3396 5773 3404
rect 6407 3396 6593 3404
rect 4527 3376 4604 3384
rect 4647 3376 4793 3384
rect 4836 3376 4964 3384
rect 1327 3356 1353 3364
rect 1547 3356 1773 3364
rect 4836 3364 4844 3376
rect 4787 3356 4844 3364
rect 4956 3364 4964 3376
rect 5507 3376 5753 3384
rect 6047 3376 6093 3384
rect 6307 3376 6493 3384
rect 6687 3376 6773 3384
rect 6827 3376 6873 3384
rect 4956 3356 5413 3364
rect 5607 3356 5673 3364
rect 387 3336 473 3344
rect 1207 3336 1264 3344
rect 1187 3316 1224 3324
rect 127 3297 173 3305
rect 287 3296 553 3304
rect 607 3296 733 3304
rect 787 3297 833 3305
rect 1216 3307 1224 3316
rect 947 3296 993 3304
rect 1216 3296 1233 3307
rect 1220 3293 1233 3296
rect 1256 3287 1264 3336
rect 2247 3336 2273 3344
rect 2287 3336 2393 3344
rect 2547 3336 2653 3344
rect 3047 3336 3253 3344
rect 3327 3336 3433 3344
rect 3527 3336 3633 3344
rect 3687 3336 4213 3344
rect 5547 3336 5573 3344
rect 6127 3336 6433 3344
rect 6487 3336 6553 3344
rect 1516 3316 1613 3324
rect 1327 3296 1373 3304
rect 1387 3296 1473 3304
rect 1256 3276 1273 3287
rect 1260 3273 1273 3276
rect 1516 3267 1524 3316
rect 1707 3316 1853 3324
rect 1987 3316 2033 3324
rect 4047 3316 4113 3324
rect 4956 3316 5093 3324
rect 1587 3297 1633 3305
rect 1947 3296 2053 3304
rect 1776 3284 1784 3294
rect 2327 3296 2373 3304
rect 2467 3297 2573 3305
rect 2747 3297 2773 3305
rect 2827 3297 2913 3305
rect 2967 3296 3053 3304
rect 3367 3296 3473 3304
rect 4956 3307 4964 3316
rect 5427 3316 5473 3324
rect 6147 3316 6233 3324
rect 6587 3316 6633 3324
rect 1756 3280 1784 3284
rect 1753 3276 1784 3280
rect 3156 3284 3164 3294
rect 3647 3296 3713 3304
rect 4307 3304 4320 3307
rect 4307 3293 4324 3304
rect 4436 3300 4873 3304
rect 3156 3276 3233 3284
rect 1753 3267 1767 3276
rect 3887 3276 3993 3284
rect 587 3255 653 3263
rect 847 3256 913 3264
rect 967 3256 1073 3264
rect 1627 3255 1693 3263
rect 1807 3256 2164 3264
rect 147 3236 333 3244
rect 347 3236 393 3244
rect 627 3236 693 3244
rect 707 3236 773 3244
rect 827 3236 953 3244
rect 2156 3244 2164 3256
rect 2387 3255 2433 3263
rect 2807 3256 2933 3264
rect 3067 3255 3133 3263
rect 3267 3255 3293 3263
rect 3727 3256 3853 3264
rect 2156 3236 2173 3244
rect 2187 3236 2293 3244
rect 2487 3236 2733 3244
rect 3207 3236 3333 3244
rect 3576 3244 3584 3252
rect 4316 3247 4324 3293
rect 4433 3296 4873 3300
rect 4433 3287 4447 3296
rect 4947 3296 4964 3307
rect 4947 3293 4960 3296
rect 5447 3296 5513 3304
rect 5767 3297 6093 3305
rect 6267 3296 6353 3304
rect 6600 3304 6613 3307
rect 6596 3293 6613 3304
rect 6707 3296 6813 3304
rect 6867 3296 6913 3304
rect 4887 3255 4973 3263
rect 5053 3264 5067 3273
rect 5107 3275 5193 3283
rect 5387 3277 5453 3285
rect 5616 3267 5624 3293
rect 5936 3276 6093 3284
rect 5053 3260 5084 3264
rect 5056 3256 5084 3260
rect 5076 3247 5084 3256
rect 5936 3264 5944 3276
rect 6107 3276 6133 3284
rect 6247 3280 6324 3284
rect 6247 3276 6327 3280
rect 5707 3256 5944 3264
rect 6176 3247 6184 3273
rect 6313 3267 6327 3276
rect 6596 3284 6604 3293
rect 6447 3276 6604 3284
rect 6596 3267 6604 3276
rect 6596 3256 6613 3267
rect 6600 3253 6613 3256
rect 6687 3255 6733 3263
rect 3576 3236 3633 3244
rect 4607 3236 4853 3244
rect 4867 3236 5053 3244
rect 5076 3236 5093 3247
rect 5080 3233 5093 3236
rect 5347 3236 5624 3244
rect 1747 3216 1953 3224
rect 2087 3216 2113 3224
rect 2127 3216 2153 3224
rect 3407 3216 3613 3224
rect 4347 3216 4433 3224
rect 4876 3216 5193 3224
rect 187 3196 793 3204
rect 1067 3196 1173 3204
rect 1667 3196 1793 3204
rect 1887 3196 1953 3204
rect 2707 3196 3353 3204
rect 3447 3196 4133 3204
rect 507 3176 1393 3184
rect 1867 3176 1993 3184
rect 2007 3176 2253 3184
rect 2896 3176 3073 3184
rect 1287 3156 1333 3164
rect 2896 3164 2904 3176
rect 4876 3184 4884 3216
rect 5347 3216 5392 3224
rect 5427 3216 5553 3224
rect 5567 3216 5593 3224
rect 5616 3224 5624 3236
rect 5727 3236 5884 3244
rect 5616 3216 5853 3224
rect 5876 3224 5884 3236
rect 5876 3216 6133 3224
rect 6527 3216 6553 3224
rect 5467 3196 5692 3204
rect 5727 3196 6093 3204
rect 6287 3196 6493 3204
rect 6647 3196 6673 3204
rect 4487 3176 4884 3184
rect 5367 3176 5393 3184
rect 5447 3176 5773 3184
rect 5847 3176 5953 3184
rect 6327 3176 6553 3184
rect 6707 3176 6753 3184
rect 1427 3156 2904 3164
rect 4187 3156 4353 3164
rect 5067 3156 5413 3164
rect 6147 3156 6233 3164
rect 6247 3156 6472 3164
rect 6507 3156 6593 3164
rect 1727 3136 2393 3144
rect 2407 3136 2553 3144
rect 2567 3136 2833 3144
rect 2947 3136 3413 3144
rect 3527 3136 3653 3144
rect 4047 3136 4453 3144
rect 4587 3136 4793 3144
rect 5207 3136 5593 3144
rect 5647 3136 5673 3144
rect 6107 3136 6193 3144
rect 6447 3136 6633 3144
rect 6707 3136 6773 3144
rect 207 3116 253 3124
rect 447 3116 993 3124
rect 1347 3116 1493 3124
rect 2647 3116 2773 3124
rect 2987 3116 3173 3124
rect 4567 3116 4833 3124
rect 5047 3116 5233 3124
rect 5427 3116 5453 3124
rect 5707 3116 5733 3124
rect 5787 3116 6133 3124
rect 6196 3124 6204 3133
rect 6196 3116 6333 3124
rect 6487 3116 6833 3124
rect 4027 3096 4053 3104
rect 4067 3096 4293 3104
rect 5036 3104 5044 3113
rect 4307 3096 5044 3104
rect 5107 3096 5173 3104
rect 5307 3096 5393 3104
rect 5467 3096 5513 3104
rect 5527 3096 5633 3104
rect 5947 3096 6313 3104
rect 6627 3096 6893 3104
rect 1547 3076 2413 3084
rect 2507 3076 2653 3084
rect 4087 3076 4473 3084
rect 5247 3076 5733 3084
rect 6087 3076 6112 3084
rect 6147 3076 6393 3084
rect 6467 3076 6793 3084
rect 407 3056 773 3064
rect 1167 3056 1413 3064
rect 3427 3056 3553 3064
rect 3627 3056 4013 3064
rect 4596 3056 4753 3064
rect 487 3036 2673 3044
rect 3376 3036 3593 3044
rect 47 3016 93 3024
rect 1267 3016 1313 3024
rect 1807 3016 1893 3024
rect 2347 3016 2393 3024
rect 2947 3016 2973 3024
rect 607 2996 673 3004
rect 987 2997 1053 3005
rect 1187 2997 1233 3005
rect 1467 2997 1493 3005
rect 1667 2997 1713 3005
rect 736 2984 744 2994
rect 736 2976 924 2984
rect 87 2956 333 2964
rect 447 2956 513 2964
rect 587 2956 713 2964
rect 807 2955 893 2963
rect 916 2964 924 2976
rect 916 2956 1073 2964
rect 1096 2964 1104 2994
rect 1096 2956 1133 2964
rect 1147 2956 1253 2964
rect 1616 2964 1624 2994
rect 1767 2996 1893 3004
rect 2287 2996 2433 3004
rect 2447 2996 2593 3004
rect 2607 2996 2733 3004
rect 2156 2967 2164 2993
rect 2867 2996 2913 3004
rect 3007 2996 3033 3004
rect 3187 2997 3233 3005
rect 3287 2996 3353 3004
rect 3376 3004 3384 3036
rect 3707 3036 4073 3044
rect 4596 3044 4604 3056
rect 4827 3056 5184 3064
rect 4227 3036 4604 3044
rect 5176 3044 5184 3056
rect 5327 3056 5513 3064
rect 5607 3056 5713 3064
rect 6247 3056 6413 3064
rect 6566 3053 6567 3060
rect 6587 3056 6673 3064
rect 4807 3036 4944 3044
rect 5176 3036 5473 3044
rect 3887 3016 4093 3024
rect 4627 3016 4653 3024
rect 4667 3016 4773 3024
rect 4867 3024 4880 3027
rect 4867 3013 4884 3024
rect 4936 3024 4944 3036
rect 5747 3036 5773 3044
rect 6147 3036 6433 3044
rect 6553 3044 6567 3053
rect 6553 3040 6853 3044
rect 6556 3036 6853 3040
rect 4936 3016 5373 3024
rect 5627 3016 5693 3024
rect 3367 2996 3384 3004
rect 3447 2997 3472 3005
rect 3507 2997 3593 3005
rect 3787 2997 3833 3005
rect 3947 2996 3993 3004
rect 2187 2976 2333 2984
rect 1616 2956 1673 2964
rect 1787 2955 1993 2963
rect 2067 2955 2093 2963
rect 2227 2956 2293 2964
rect 2427 2956 2472 2964
rect 2507 2955 2573 2963
rect 2767 2956 2893 2964
rect 3107 2956 3193 2964
rect 3307 2956 3513 2964
rect 3627 2956 3653 2964
rect 3736 2947 3744 2994
rect 4287 2996 4313 3004
rect 4367 2997 4433 3005
rect 4596 2996 4813 3004
rect 4596 2984 4604 2996
rect 4876 3004 4884 3013
rect 4876 2996 4904 3004
rect 4896 2986 4904 2996
rect 4916 2987 4924 3013
rect 5296 2996 5493 3004
rect 3956 2976 4604 2984
rect 3956 2966 3964 2976
rect 3887 2955 3913 2963
rect 4007 2955 4133 2963
rect 4147 2956 4253 2964
rect 4327 2955 4413 2963
rect 4667 2955 4773 2963
rect 907 2936 1113 2944
rect 1487 2936 1713 2944
rect 1976 2936 2793 2944
rect 387 2916 473 2924
rect 487 2916 713 2924
rect 1976 2924 1984 2936
rect 3227 2936 3253 2944
rect 3396 2936 3453 2944
rect 1027 2916 1984 2924
rect 2007 2916 2253 2924
rect 3027 2916 3093 2924
rect 3396 2924 3404 2936
rect 4867 2936 4933 2944
rect 5076 2944 5084 2974
rect 5207 2976 5273 2984
rect 5296 2964 5304 2996
rect 6427 2997 6453 3005
rect 6727 2997 6753 3005
rect 5807 2976 5912 2984
rect 5247 2956 5304 2964
rect 5407 2955 5433 2963
rect 5447 2956 5573 2964
rect 5076 2936 5213 2944
rect 3167 2916 3404 2924
rect 3427 2916 3493 2924
rect 3587 2916 3753 2924
rect 4056 2916 4353 2924
rect 767 2896 993 2904
rect 1467 2896 2133 2904
rect 2687 2896 3293 2904
rect 4056 2904 4064 2916
rect 4447 2916 4833 2924
rect 5427 2916 5693 2924
rect 3656 2896 4064 2904
rect 1247 2876 1773 2884
rect 2107 2876 2193 2884
rect 2667 2876 2933 2884
rect 3067 2876 3113 2884
rect 3656 2884 3664 2896
rect 4087 2896 4333 2904
rect 5056 2896 5253 2904
rect 3467 2876 3664 2884
rect 3676 2876 3813 2884
rect 1407 2856 1653 2864
rect 1727 2856 1813 2864
rect 2707 2856 2833 2864
rect 3367 2856 3433 2864
rect 3676 2864 3684 2876
rect 4107 2876 4213 2884
rect 4467 2876 4833 2884
rect 4887 2876 4953 2884
rect 3647 2856 3684 2864
rect 3867 2856 3933 2864
rect 4027 2856 4273 2864
rect 5056 2864 5064 2896
rect 5307 2896 5493 2904
rect 5107 2876 5313 2884
rect 5367 2876 5453 2884
rect 5547 2876 5593 2884
rect 5807 2876 5893 2884
rect 5936 2884 5944 2974
rect 6087 2975 6113 2983
rect 6327 2956 6344 2964
rect 6187 2936 6293 2944
rect 6336 2944 6344 2956
rect 6447 2955 6533 2963
rect 6827 2955 6853 2963
rect 6336 2936 6413 2944
rect 6727 2936 6753 2944
rect 6087 2916 6153 2924
rect 6207 2896 6573 2904
rect 6667 2896 6773 2904
rect 5936 2876 5973 2884
rect 6427 2876 6453 2884
rect 5027 2856 5064 2864
rect 5507 2856 6133 2864
rect 6487 2856 6713 2864
rect 67 2836 233 2844
rect 427 2836 813 2844
rect 827 2836 873 2844
rect 887 2836 1093 2844
rect 1447 2836 1613 2844
rect 1627 2836 1693 2844
rect 1947 2836 2233 2844
rect 2607 2836 2673 2844
rect 2787 2836 2813 2844
rect 2927 2836 3073 2844
rect 3187 2836 3473 2844
rect 3487 2836 3573 2844
rect 3587 2836 3793 2844
rect 3807 2836 4433 2844
rect 4627 2836 4673 2844
rect 5127 2836 5173 2844
rect 5487 2836 5533 2844
rect 6047 2836 6073 2844
rect 6307 2836 6393 2844
rect 107 2816 193 2824
rect 947 2816 973 2824
rect 1187 2816 1573 2824
rect 1707 2816 1733 2824
rect 1747 2816 2173 2824
rect 2867 2816 3133 2824
rect 3207 2816 3353 2824
rect 3827 2816 4173 2824
rect 4787 2816 4833 2824
rect 4847 2816 5093 2824
rect 5667 2816 5813 2824
rect 5967 2816 6113 2824
rect 6207 2816 6473 2824
rect 427 2796 673 2804
rect 3707 2796 3773 2804
rect 4367 2796 4493 2804
rect 4547 2796 4573 2804
rect 5147 2796 5233 2804
rect 5767 2796 6173 2804
rect 167 2777 213 2785
rect 116 2727 124 2774
rect 276 2747 284 2774
rect 316 2764 324 2774
rect 787 2776 853 2784
rect 867 2777 913 2785
rect 1007 2777 1053 2785
rect 267 2736 284 2747
rect 296 2756 324 2764
rect 336 2756 393 2764
rect 267 2733 280 2736
rect 296 2727 304 2756
rect 336 2746 344 2756
rect 547 2755 693 2763
rect 1456 2747 1464 2773
rect 1507 2776 1533 2784
rect 947 2736 973 2744
rect 1087 2736 1253 2744
rect 1267 2736 1413 2744
rect 1556 2746 1564 2793
rect 1787 2777 1833 2785
rect 1967 2777 2133 2785
rect 2227 2776 2493 2784
rect 2827 2777 2873 2785
rect 3007 2777 3053 2785
rect 3327 2777 3473 2785
rect 3547 2777 3613 2785
rect 3747 2776 3833 2784
rect 3816 2747 3824 2776
rect 3927 2776 4053 2784
rect 4176 2764 4184 2774
rect 4307 2776 4633 2784
rect 4707 2777 4753 2785
rect 4767 2777 4893 2785
rect 4176 2756 4253 2764
rect 1607 2736 1673 2744
rect 1687 2736 1753 2744
rect 1847 2736 1913 2744
rect 2007 2735 2033 2743
rect 2296 2736 2353 2744
rect 287 2716 304 2727
rect 287 2713 300 2716
rect 407 2716 433 2724
rect 2296 2724 2304 2736
rect 2587 2735 2653 2743
rect 2807 2735 2893 2743
rect 2967 2736 3113 2744
rect 3127 2736 3173 2744
rect 4207 2736 4333 2744
rect 4527 2735 4613 2743
rect 4687 2736 4713 2744
rect 4767 2735 4793 2743
rect 5056 2744 5064 2774
rect 5127 2776 5333 2784
rect 5467 2776 5493 2784
rect 5516 2776 5573 2784
rect 5516 2764 5524 2776
rect 5396 2756 5524 2764
rect 5696 2764 5704 2774
rect 5696 2756 6053 2764
rect 5007 2736 5064 2744
rect 5107 2735 5153 2743
rect 5167 2735 5193 2743
rect 5396 2744 5404 2756
rect 6076 2764 6084 2774
rect 6487 2776 6613 2784
rect 6076 2756 6193 2764
rect 6276 2747 6284 2773
rect 5387 2736 5404 2744
rect 5567 2735 5613 2743
rect 5947 2736 5973 2744
rect 6316 2744 6324 2774
rect 6316 2736 6364 2744
rect 2227 2716 2304 2724
rect 3807 2716 3853 2724
rect 5067 2716 5113 2724
rect 5687 2716 5873 2724
rect 6356 2724 6364 2736
rect 6387 2736 6773 2744
rect 6356 2716 6493 2724
rect 6507 2716 6593 2724
rect 6796 2724 6804 2774
rect 6836 2747 6844 2773
rect 6607 2716 6804 2724
rect 87 2696 133 2704
rect 207 2696 373 2704
rect 1287 2696 1693 2704
rect 1847 2696 1993 2704
rect 2247 2696 2693 2704
rect 3627 2696 4673 2704
rect 5867 2696 6013 2704
rect 6207 2696 6373 2704
rect 6647 2696 6733 2704
rect 6747 2696 6813 2704
rect 1787 2676 1813 2684
rect 3787 2676 3973 2684
rect 3987 2676 4293 2684
rect 4307 2676 5053 2684
rect 5107 2676 5233 2684
rect 5247 2676 5533 2684
rect 5827 2676 6133 2684
rect 6427 2676 6873 2684
rect 127 2656 173 2664
rect 247 2656 353 2664
rect 1247 2656 1553 2664
rect 1927 2656 2013 2664
rect 2027 2656 2333 2664
rect 2347 2656 2473 2664
rect 2887 2656 3093 2664
rect 3107 2656 3913 2664
rect 4267 2656 4373 2664
rect 4567 2656 4753 2664
rect 4807 2656 4913 2664
rect 5847 2656 5932 2664
rect 5967 2656 6293 2664
rect 6347 2656 6953 2664
rect 227 2636 853 2644
rect 1687 2636 1953 2644
rect 2047 2636 2213 2644
rect 2507 2636 2593 2644
rect 4947 2636 5293 2644
rect 5367 2636 5433 2644
rect 5856 2636 5904 2644
rect 307 2616 1133 2624
rect 3827 2616 4993 2624
rect 5096 2616 5273 2624
rect 467 2596 1213 2604
rect 1387 2596 1553 2604
rect 1667 2596 2513 2604
rect 3407 2596 3713 2604
rect 3847 2596 4013 2604
rect 4307 2596 4553 2604
rect 4607 2596 4733 2604
rect 5096 2604 5104 2616
rect 5856 2624 5864 2636
rect 5527 2616 5864 2624
rect 5896 2624 5904 2636
rect 6107 2636 6513 2644
rect 6627 2636 6773 2644
rect 5896 2616 5953 2624
rect 6307 2616 6393 2624
rect 6536 2616 6833 2624
rect 4867 2596 5104 2604
rect 5427 2596 5453 2604
rect 5887 2596 6053 2604
rect 6536 2604 6544 2616
rect 6167 2596 6544 2604
rect 707 2576 993 2584
rect 1676 2576 2493 2584
rect 967 2556 1253 2564
rect 1676 2564 1684 2576
rect 2947 2576 3653 2584
rect 3787 2576 3813 2584
rect 3907 2576 3953 2584
rect 4427 2576 5213 2584
rect 5387 2576 5733 2584
rect 6087 2576 6593 2584
rect 1567 2556 1684 2564
rect 2407 2556 2813 2564
rect 3847 2556 4153 2564
rect 4647 2556 4693 2564
rect 5767 2556 5873 2564
rect 6227 2556 6373 2564
rect 6487 2556 6913 2564
rect 316 2536 793 2544
rect 316 2527 324 2536
rect 1427 2536 1673 2544
rect 1927 2536 2033 2544
rect 2087 2536 2153 2544
rect 4987 2536 5133 2544
rect 5507 2536 5593 2544
rect 6087 2536 6533 2544
rect 127 2516 253 2524
rect 267 2516 313 2524
rect 687 2516 833 2524
rect 847 2516 1373 2524
rect 1716 2516 1773 2524
rect 1716 2504 1724 2516
rect 1827 2516 2373 2524
rect 2547 2516 2933 2524
rect 3107 2516 3553 2524
rect 3927 2516 4413 2524
rect 4527 2516 4553 2524
rect 4567 2516 4813 2524
rect 5387 2516 5473 2524
rect 5647 2516 5713 2524
rect 6147 2516 6213 2524
rect 6467 2516 6513 2524
rect 6767 2516 6833 2524
rect 1587 2496 1724 2504
rect 2127 2496 2393 2504
rect 2487 2496 2993 2504
rect 3496 2496 3653 2504
rect 547 2476 753 2484
rect 1067 2477 1093 2485
rect 1247 2476 1493 2484
rect 1687 2477 1733 2485
rect 1536 2447 1544 2473
rect 1616 2447 1624 2474
rect 2207 2477 2273 2485
rect 2687 2476 2873 2484
rect 2927 2477 2973 2485
rect 3047 2476 3173 2484
rect 3227 2476 3333 2484
rect 3347 2476 3473 2484
rect 1667 2456 1813 2464
rect 307 2435 353 2443
rect 507 2436 593 2444
rect 607 2436 693 2444
rect 827 2436 973 2444
rect 1167 2435 1233 2443
rect 1616 2436 1633 2447
rect 1620 2433 1633 2436
rect 1976 2444 1984 2473
rect 1887 2436 1984 2444
rect 2107 2436 2193 2444
rect 2307 2436 2353 2444
rect 3496 2446 3504 2496
rect 3667 2496 3833 2504
rect 4027 2496 4113 2504
rect 4447 2496 4584 2504
rect 3540 2484 3553 2487
rect 2727 2436 2853 2444
rect 2867 2435 2953 2443
rect 3367 2435 3393 2443
rect 3516 2427 3524 2474
rect 3536 2473 3553 2484
rect 3767 2476 3873 2484
rect 3887 2476 4173 2484
rect 4187 2476 4313 2484
rect 4576 2487 4584 2496
rect 5027 2496 5053 2504
rect 5236 2496 5353 2504
rect 4566 2473 4567 2480
rect 4587 2477 4753 2485
rect 4847 2476 4893 2484
rect 4947 2476 5084 2484
rect 3536 2446 3544 2473
rect 4553 2467 4567 2473
rect 4553 2466 4580 2467
rect 4553 2460 4573 2466
rect 4556 2456 4573 2460
rect 4560 2453 4573 2456
rect 5076 2447 5084 2476
rect 5236 2484 5244 2496
rect 5506 2493 5507 2500
rect 5527 2496 5573 2504
rect 5587 2497 5633 2505
rect 5093 2464 5107 2473
rect 5176 2476 5244 2484
rect 5493 2484 5507 2493
rect 5747 2496 5944 2504
rect 5493 2480 5564 2484
rect 5496 2476 5567 2480
rect 5093 2460 5133 2464
rect 5096 2456 5133 2460
rect 5176 2466 5184 2476
rect 5553 2467 5567 2476
rect 3807 2435 3993 2443
rect 4047 2435 4073 2443
rect 4127 2435 4153 2443
rect 4207 2435 4393 2443
rect 4467 2436 4493 2444
rect 4507 2436 4653 2444
rect 4667 2436 4873 2444
rect 5007 2435 5033 2443
rect 5076 2436 5093 2447
rect 5080 2433 5093 2436
rect 5356 2444 5364 2454
rect 5387 2460 5484 2464
rect 5387 2456 5487 2460
rect 5227 2436 5364 2444
rect 5473 2447 5487 2456
rect 5726 2453 5727 2460
rect 5747 2457 5873 2465
rect 5620 2444 5633 2447
rect 5616 2433 5633 2444
rect 5713 2444 5727 2453
rect 5936 2447 5944 2496
rect 6607 2496 6673 2504
rect 6807 2496 6853 2504
rect 6027 2476 6113 2484
rect 6127 2477 6153 2485
rect 6207 2476 6253 2484
rect 6276 2476 6333 2484
rect 6276 2464 6284 2476
rect 6527 2476 6564 2484
rect 6176 2456 6284 2464
rect 6556 2464 6564 2476
rect 6587 2477 6613 2485
rect 6556 2456 6624 2464
rect 5713 2440 5924 2444
rect 5716 2436 5924 2440
rect 787 2416 873 2424
rect 967 2416 1013 2424
rect 1567 2416 1673 2424
rect 1687 2416 1773 2424
rect 1847 2416 1933 2424
rect 3847 2416 3953 2424
rect 4287 2416 4413 2424
rect 4547 2416 4573 2424
rect 5616 2424 5624 2433
rect 5527 2416 5624 2424
rect 5916 2424 5924 2436
rect 6176 2444 6184 2456
rect 6147 2436 6184 2444
rect 6287 2436 6433 2444
rect 6487 2436 6533 2444
rect 6616 2444 6624 2456
rect 6696 2447 6704 2473
rect 6616 2436 6633 2444
rect 6747 2436 6813 2444
rect 6867 2435 6893 2443
rect 5916 2416 6124 2424
rect 147 2396 173 2404
rect 187 2396 433 2404
rect 447 2396 533 2404
rect 947 2396 1113 2404
rect 1167 2396 1193 2404
rect 2107 2396 2153 2404
rect 3687 2396 3753 2404
rect 4007 2396 4053 2404
rect 4367 2396 4393 2404
rect 4407 2396 4693 2404
rect 4847 2396 5073 2404
rect 5187 2396 5213 2404
rect 5647 2396 5913 2404
rect 6000 2406 6020 2407
rect 6007 2404 6020 2406
rect 6116 2404 6124 2416
rect 6307 2416 6393 2424
rect 6467 2416 6553 2424
rect 6007 2393 6024 2404
rect 6116 2396 6333 2404
rect 6687 2396 6773 2404
rect 1507 2376 1553 2384
rect 2987 2376 3173 2384
rect 4867 2376 4913 2384
rect 5696 2380 5973 2384
rect 5693 2376 5973 2380
rect 5693 2367 5707 2376
rect 6016 2384 6024 2393
rect 6016 2376 6133 2384
rect 6467 2376 6693 2384
rect 787 2356 1653 2364
rect 2507 2356 3433 2364
rect 3487 2356 3773 2364
rect 4227 2356 4333 2364
rect 4667 2356 4933 2364
rect 4987 2356 5013 2364
rect 5036 2356 5173 2364
rect 67 2336 193 2344
rect 487 2336 853 2344
rect 1927 2336 1993 2344
rect 2407 2336 2512 2344
rect 2547 2336 2613 2344
rect 2767 2336 2973 2344
rect 3916 2336 4513 2344
rect 256 2304 264 2333
rect 3916 2327 3924 2336
rect 5036 2344 5044 2356
rect 5227 2356 5484 2364
rect 4907 2336 5044 2344
rect 5476 2344 5484 2356
rect 5507 2356 5533 2364
rect 6607 2356 6753 2364
rect 6767 2356 6793 2364
rect 5476 2336 5633 2344
rect 5727 2336 5993 2344
rect 6287 2336 6353 2344
rect 6627 2336 6713 2344
rect 927 2316 1473 2324
rect 1767 2316 2013 2324
rect 2027 2316 2073 2324
rect 3127 2316 3633 2324
rect 3767 2316 3853 2324
rect 3907 2316 3924 2327
rect 3907 2313 3920 2316
rect 4127 2316 4233 2324
rect 4547 2316 4713 2324
rect 4787 2316 4833 2324
rect 4887 2316 5113 2324
rect 5467 2316 5493 2324
rect 5547 2316 5593 2324
rect 5736 2316 5873 2324
rect 236 2296 264 2304
rect 236 2264 244 2296
rect 1227 2296 1333 2304
rect 1547 2296 1733 2304
rect 1887 2296 1953 2304
rect 2387 2296 2573 2304
rect 2947 2296 3073 2304
rect 3707 2296 3733 2304
rect 3947 2296 4013 2304
rect 4267 2296 4493 2304
rect 5147 2296 5333 2304
rect 5736 2304 5744 2316
rect 5887 2316 5964 2324
rect 5647 2296 5744 2304
rect 5956 2304 5964 2316
rect 6387 2316 6413 2324
rect 5956 2296 6033 2304
rect 6127 2296 6173 2304
rect 6327 2296 6533 2304
rect 6547 2296 6684 2304
rect 387 2276 733 2284
rect 1847 2276 2033 2284
rect 2047 2276 2064 2284
rect 216 2256 244 2264
rect 56 2204 64 2233
rect 216 2227 224 2256
rect 947 2257 993 2265
rect 1107 2256 1153 2264
rect 1267 2257 1293 2265
rect 1513 2264 1527 2273
rect 1513 2260 1553 2264
rect 1516 2256 1553 2260
rect 1807 2257 1853 2265
rect 1616 2227 1624 2254
rect 1867 2257 1893 2265
rect 2056 2267 2064 2276
rect 3247 2276 3433 2284
rect 3527 2276 3593 2284
rect 3607 2276 3893 2284
rect 4527 2276 4793 2284
rect 4867 2276 4913 2284
rect 4936 2276 4993 2284
rect 2067 2256 2153 2264
rect 2247 2256 2313 2264
rect 2336 2244 2344 2273
rect 2407 2257 2433 2265
rect 2907 2257 3033 2265
rect 3207 2257 3233 2265
rect 3287 2256 3373 2264
rect 3807 2256 3873 2264
rect 3987 2257 4033 2265
rect 4047 2256 4153 2264
rect 4467 2257 4493 2265
rect 4936 2264 4944 2276
rect 5427 2276 5473 2284
rect 5947 2276 6053 2284
rect 6207 2276 6253 2284
rect 6347 2276 6433 2284
rect 4547 2256 4584 2264
rect 207 2216 224 2227
rect 207 2213 220 2216
rect 607 2215 673 2223
rect 887 2216 933 2224
rect 1027 2216 1073 2224
rect 1127 2216 1173 2224
rect 1187 2216 1433 2224
rect 1607 2216 1624 2227
rect 1636 2236 2344 2244
rect 1636 2226 1644 2236
rect 2336 2226 2344 2236
rect 4027 2236 4393 2244
rect 1607 2213 1620 2216
rect 1687 2215 1893 2223
rect 1987 2215 2052 2223
rect 2087 2215 2133 2223
rect 2187 2215 2233 2223
rect 2513 2224 2527 2233
rect 2467 2220 2527 2224
rect 2467 2216 2524 2220
rect 2747 2216 2933 2224
rect 2987 2215 3053 2223
rect 3187 2215 3293 2223
rect 3387 2215 3453 2223
rect 3887 2215 3913 2223
rect 4067 2215 4133 2223
rect 4247 2215 4273 2223
rect 4396 2224 4404 2233
rect 4576 2227 4584 2256
rect 4916 2256 4944 2264
rect 4396 2216 4473 2224
rect 4487 2216 4513 2224
rect 4916 2226 4924 2256
rect 5047 2256 5093 2264
rect 5207 2257 5253 2265
rect 5307 2256 5373 2264
rect 5667 2256 5733 2264
rect 5827 2256 5913 2264
rect 5776 2227 5784 2254
rect 5067 2216 5213 2224
rect 5227 2215 5273 2223
rect 5327 2215 5353 2223
rect 5447 2216 5513 2224
rect 5767 2216 5784 2227
rect 5767 2213 5780 2216
rect 5996 2224 6004 2254
rect 6047 2256 6084 2264
rect 6076 2244 6084 2256
rect 6107 2256 6133 2264
rect 6176 2244 6184 2254
rect 6507 2256 6653 2264
rect 6293 2244 6307 2253
rect 6076 2236 6164 2244
rect 6176 2240 6307 2244
rect 6176 2236 6304 2240
rect 5867 2216 6004 2224
rect 6156 2224 6164 2236
rect 6156 2216 6213 2224
rect 6236 2224 6244 2236
rect 6236 2216 6293 2224
rect 6527 2216 6593 2224
rect 6676 2226 6684 2296
rect 6767 2296 6913 2304
rect 6707 2256 6753 2264
rect 6847 2256 7004 2264
rect 6836 2224 6844 2254
rect 6727 2216 6844 2224
rect 6867 2216 6893 2224
rect 6907 2216 6933 2224
rect 6996 2216 7004 2256
rect 47 2196 64 2204
rect 1527 2196 2284 2204
rect 2276 2187 2284 2196
rect 3707 2196 3773 2204
rect 3867 2196 4093 2204
rect 4327 2196 4533 2204
rect 4807 2196 4953 2204
rect 4967 2196 5033 2204
rect 5647 2196 5953 2204
rect 647 2176 1473 2184
rect 1667 2176 1733 2184
rect 2027 2176 2173 2184
rect 2287 2176 2393 2184
rect 2907 2176 3013 2184
rect 3267 2176 3413 2184
rect 3427 2176 3613 2184
rect 4227 2176 4733 2184
rect 5527 2176 5713 2184
rect 5927 2176 6013 2184
rect 727 2156 913 2164
rect 1767 2156 1933 2164
rect 2967 2156 3093 2164
rect 4147 2156 4193 2164
rect 4547 2156 5493 2164
rect 5587 2156 5693 2164
rect 5847 2156 6093 2164
rect 1327 2136 1493 2144
rect 2167 2136 2253 2144
rect 2547 2136 3973 2144
rect 3987 2136 4293 2144
rect 4307 2136 4453 2144
rect 5367 2136 5553 2144
rect 6087 2136 6113 2144
rect 6127 2136 6513 2144
rect 487 2116 573 2124
rect 1607 2116 2244 2124
rect 427 2096 753 2104
rect 1227 2096 1313 2104
rect 1487 2096 2093 2104
rect 2107 2096 2193 2104
rect 2236 2104 2244 2116
rect 3107 2116 3733 2124
rect 3747 2116 3953 2124
rect 4107 2116 4853 2124
rect 5107 2116 5493 2124
rect 5627 2116 5973 2124
rect 5987 2116 6253 2124
rect 6607 2116 6913 2124
rect 2236 2096 2293 2104
rect 2607 2096 2673 2104
rect 3167 2096 3433 2104
rect 4207 2096 4533 2104
rect 5087 2096 5512 2104
rect 5547 2096 5733 2104
rect 5827 2096 5873 2104
rect 6147 2096 6233 2104
rect 6487 2096 6753 2104
rect 3547 2076 3913 2084
rect 4647 2076 4873 2084
rect 5187 2076 5613 2084
rect 5767 2076 6153 2084
rect 6167 2076 6733 2084
rect 807 2056 1513 2064
rect 1647 2056 1853 2064
rect 3387 2056 4013 2064
rect 4067 2056 4313 2064
rect 5607 2056 6133 2064
rect 6267 2056 6293 2064
rect 6447 2056 6533 2064
rect 447 2036 493 2044
rect 2547 2036 2853 2044
rect 3907 2036 4193 2044
rect 4567 2036 5033 2044
rect 5047 2036 5093 2044
rect 5596 2044 5604 2053
rect 5407 2036 5604 2044
rect 6207 2036 6313 2044
rect 6327 2036 6613 2044
rect 6747 2036 6773 2044
rect 6787 2036 6853 2044
rect 1047 2016 1693 2024
rect 4427 2016 5073 2024
rect 5747 2016 5873 2024
rect 5947 2016 6113 2024
rect 527 1996 673 2004
rect 1487 1996 1553 2004
rect 1727 1996 1953 2004
rect 2427 1996 2733 2004
rect 2847 1996 2953 2004
rect 3647 1996 3913 2004
rect 4527 1996 4613 2004
rect 5167 1996 5373 2004
rect 6167 1996 6453 2004
rect 6547 1996 6773 2004
rect 1587 1976 1613 1984
rect 1827 1976 2053 1984
rect 3027 1977 3073 1985
rect 3087 1976 3344 1984
rect 267 1957 293 1965
rect 607 1957 633 1965
rect 767 1957 833 1965
rect 1247 1956 1373 1964
rect 1387 1956 1413 1964
rect 116 1927 124 1954
rect 107 1916 124 1927
rect 107 1913 120 1916
rect 156 1907 164 1954
rect 187 1916 253 1924
rect 336 1904 344 1954
rect 476 1944 484 1954
rect 376 1936 484 1944
rect 876 1944 884 1954
rect 876 1936 924 1944
rect 376 1924 384 1936
rect 367 1916 384 1924
rect 407 1916 493 1924
rect 707 1915 793 1923
rect 916 1924 924 1936
rect 916 1916 1173 1924
rect 307 1896 344 1904
rect 907 1896 1053 1904
rect 1196 1887 1204 1954
rect 1567 1957 1773 1965
rect 2027 1957 2113 1965
rect 2247 1956 2313 1964
rect 2327 1956 2353 1964
rect 2467 1956 2513 1964
rect 3336 1964 3344 1976
rect 3436 1976 3473 1984
rect 3436 1964 3444 1976
rect 3787 1976 4053 1984
rect 4267 1976 4313 1984
rect 4396 1976 4693 1984
rect 3336 1956 3444 1964
rect 3876 1956 4073 1964
rect 2647 1936 2833 1944
rect 2907 1936 3053 1944
rect 3187 1937 3453 1945
rect 3876 1946 3884 1956
rect 4167 1957 4193 1965
rect 4247 1957 4333 1965
rect 4396 1964 4404 1976
rect 4347 1956 4404 1964
rect 4596 1967 4604 1976
rect 4747 1976 4773 1984
rect 5127 1976 5173 1984
rect 5467 1977 5773 1985
rect 5967 1976 6053 1984
rect 4447 1956 4493 1964
rect 5087 1956 5213 1964
rect 4660 1944 4673 1947
rect 4656 1933 4673 1944
rect 1507 1916 1673 1924
rect 1727 1916 1813 1924
rect 2127 1916 2213 1924
rect 3987 1915 4013 1923
rect 4067 1916 4153 1924
rect 4267 1915 4313 1923
rect 4656 1924 4664 1933
rect 4427 1916 4664 1924
rect 4867 1915 4913 1923
rect 5055 1924 5063 1953
rect 5336 1944 5344 1954
rect 5187 1936 5344 1944
rect 5396 1944 5404 1973
rect 5627 1956 5713 1964
rect 6007 1956 6044 1964
rect 5387 1936 5404 1944
rect 5893 1944 5907 1953
rect 5747 1940 5907 1944
rect 6036 1944 6044 1956
rect 6087 1956 6273 1964
rect 6287 1957 6473 1965
rect 6827 1957 6893 1965
rect 5747 1936 5904 1940
rect 6036 1936 6104 1944
rect 6096 1926 6104 1936
rect 5055 1916 5093 1924
rect 6247 1915 6373 1923
rect 6387 1916 6413 1924
rect 6727 1915 6833 1923
rect 1587 1896 1893 1904
rect 2087 1896 2153 1904
rect 2327 1896 2493 1904
rect 2547 1896 2573 1904
rect 3447 1896 3793 1904
rect 5127 1896 5173 1904
rect 5807 1896 5853 1904
rect 5927 1896 6173 1904
rect 6467 1896 6493 1904
rect 6567 1896 6653 1904
rect 707 1876 773 1884
rect 1187 1876 1204 1887
rect 1187 1873 1200 1876
rect 1347 1876 1493 1884
rect 1667 1876 1713 1884
rect 2987 1876 3373 1884
rect 3467 1876 3804 1884
rect 267 1856 593 1864
rect 667 1856 913 1864
rect 1227 1856 1413 1864
rect 2187 1856 2373 1864
rect 2387 1856 2413 1864
rect 2467 1856 2553 1864
rect 3467 1856 3773 1864
rect 3796 1864 3804 1876
rect 3927 1876 4213 1884
rect 4236 1876 4573 1884
rect 4236 1864 4244 1876
rect 4707 1876 4793 1884
rect 4887 1876 4953 1884
rect 4976 1876 5273 1884
rect 3796 1856 4244 1864
rect 4976 1864 4984 1876
rect 6267 1876 6293 1884
rect 6547 1876 6873 1884
rect 4627 1856 4984 1864
rect 5727 1856 5953 1864
rect 6347 1856 6413 1864
rect 1027 1836 1533 1844
rect 1967 1836 2053 1844
rect 2227 1836 2293 1844
rect 2827 1836 3353 1844
rect 3367 1836 3433 1844
rect 3447 1836 3813 1844
rect 3827 1836 3853 1844
rect 3867 1836 4573 1844
rect 4587 1836 5193 1844
rect 5207 1836 5433 1844
rect 6347 1836 6393 1844
rect 6487 1836 6633 1844
rect 867 1816 2033 1824
rect 2707 1816 2973 1824
rect 3327 1816 3393 1824
rect 3967 1816 4033 1824
rect 4307 1816 4373 1824
rect 4627 1816 4653 1824
rect 4847 1816 4973 1824
rect 5067 1816 5173 1824
rect 6187 1816 6433 1824
rect 6507 1816 6553 1824
rect 327 1796 393 1804
rect 1407 1796 1453 1804
rect 1467 1796 1513 1804
rect 3667 1796 4133 1804
rect 107 1776 493 1784
rect 1947 1776 2033 1784
rect 2747 1776 4153 1784
rect 4387 1776 4473 1784
rect 4527 1776 4553 1784
rect 787 1756 993 1764
rect 1287 1756 1593 1764
rect 2987 1756 3553 1764
rect 127 1736 353 1744
rect 367 1737 413 1745
rect 667 1737 733 1745
rect 807 1737 853 1745
rect 1047 1737 1093 1745
rect 1227 1737 1253 1745
rect 1307 1736 1353 1744
rect 1427 1736 1553 1744
rect 1687 1736 1793 1744
rect 1907 1737 1973 1745
rect 2027 1736 2113 1744
rect 2247 1736 2693 1744
rect 2707 1736 2733 1744
rect 3876 1736 3933 1744
rect 2176 1707 2184 1714
rect 2427 1715 2553 1723
rect 2647 1717 2673 1725
rect 227 1695 273 1703
rect 447 1695 473 1703
rect 727 1696 753 1704
rect 967 1696 1013 1704
rect 1207 1695 1293 1703
rect 1547 1695 1693 1703
rect 1827 1696 1913 1704
rect 2067 1695 2093 1703
rect 2167 1696 2184 1707
rect 2167 1693 2180 1696
rect 1187 1676 1333 1684
rect 1887 1676 1953 1684
rect 2567 1676 2733 1684
rect 3076 1684 3084 1713
rect 3267 1715 3453 1723
rect 3876 1724 3884 1736
rect 4007 1736 4093 1744
rect 4207 1736 4253 1744
rect 4307 1736 4413 1744
rect 4467 1736 4504 1744
rect 3656 1716 3884 1724
rect 3527 1696 3633 1704
rect 3656 1704 3664 1716
rect 4496 1707 4504 1736
rect 4756 1726 4764 1813
rect 5167 1796 5333 1804
rect 5387 1796 5473 1804
rect 6247 1796 6473 1804
rect 6527 1796 6593 1804
rect 5427 1776 5453 1784
rect 5967 1776 6053 1784
rect 6476 1784 6484 1793
rect 6476 1776 6653 1784
rect 5656 1756 6133 1764
rect 5167 1736 5233 1744
rect 5247 1736 5273 1744
rect 5467 1736 5524 1744
rect 4887 1716 4953 1724
rect 5416 1724 5424 1734
rect 5396 1720 5424 1724
rect 5393 1716 5424 1720
rect 5393 1707 5407 1716
rect 3647 1696 3664 1704
rect 3687 1695 3713 1703
rect 4287 1696 4373 1704
rect 4387 1695 4433 1703
rect 5227 1696 5293 1704
rect 5516 1687 5524 1736
rect 5656 1726 5664 1756
rect 6327 1756 6373 1764
rect 6447 1756 6533 1764
rect 6740 1764 6753 1767
rect 6736 1754 6753 1764
rect 6736 1753 6760 1754
rect 6827 1756 6893 1764
rect 6087 1737 6153 1745
rect 6356 1736 6413 1744
rect 5827 1717 5893 1725
rect 5907 1716 5993 1724
rect 6356 1707 6364 1736
rect 6687 1736 6713 1744
rect 6067 1695 6313 1703
rect 6736 1706 6744 1753
rect 6767 1736 6833 1744
rect 6936 1707 6944 1734
rect 6967 1744 6980 1747
rect 6967 1733 6984 1744
rect 6447 1695 6473 1703
rect 6667 1695 6693 1703
rect 6807 1695 6913 1703
rect 6936 1696 6953 1707
rect 6940 1693 6953 1696
rect 3047 1676 3093 1684
rect 3107 1675 3253 1683
rect 5667 1676 5853 1684
rect 5867 1676 6093 1684
rect 6847 1676 6873 1684
rect 6976 1684 6984 1733
rect 6947 1676 6984 1684
rect 1667 1656 1753 1664
rect 2167 1656 2233 1664
rect 3967 1656 4073 1664
rect 4087 1656 4853 1664
rect 4927 1656 5373 1664
rect 5387 1656 5493 1664
rect 6007 1656 6213 1664
rect 307 1636 353 1644
rect 867 1636 893 1644
rect 1267 1636 1493 1644
rect 1507 1636 2013 1644
rect 2027 1636 2073 1644
rect 3427 1636 3673 1644
rect 6547 1636 6613 1644
rect 687 1616 873 1624
rect 2147 1616 2673 1624
rect 3467 1616 3993 1624
rect 4347 1616 5393 1624
rect 287 1596 733 1604
rect 747 1596 824 1604
rect 816 1584 824 1596
rect 1727 1596 3233 1604
rect 5447 1596 5653 1604
rect 6707 1596 6813 1604
rect 816 1576 893 1584
rect 1327 1576 1553 1584
rect 2287 1576 2353 1584
rect 2887 1576 2933 1584
rect 4127 1576 4833 1584
rect 5347 1576 5393 1584
rect 5967 1576 6573 1584
rect 6667 1576 6893 1584
rect 207 1556 433 1564
rect 807 1556 1004 1564
rect 996 1547 1004 1556
rect 1087 1556 1253 1564
rect 1267 1556 1713 1564
rect 3827 1556 3873 1564
rect 3887 1556 3993 1564
rect 4907 1556 4953 1564
rect 6167 1556 6713 1564
rect 527 1536 773 1544
rect 1007 1536 1413 1544
rect 2767 1536 2973 1544
rect 3087 1536 3193 1544
rect 3236 1536 3433 1544
rect 167 1516 433 1524
rect 447 1516 633 1524
rect 827 1516 873 1524
rect 1127 1516 1313 1524
rect 1987 1516 2033 1524
rect 2047 1516 2153 1524
rect 2207 1516 2433 1524
rect 3236 1524 3244 1536
rect 3487 1536 4373 1544
rect 4387 1536 4533 1544
rect 5127 1536 5353 1544
rect 5567 1536 5593 1544
rect 5647 1536 5953 1544
rect 2527 1516 3244 1524
rect 3267 1516 3453 1524
rect 3807 1516 3893 1524
rect 4047 1516 4313 1524
rect 4627 1516 4753 1524
rect 487 1496 513 1504
rect 1627 1496 1773 1504
rect 1907 1496 3913 1504
rect 3927 1496 4233 1504
rect 4247 1496 4853 1504
rect 5727 1496 6253 1504
rect 6267 1496 6293 1504
rect 247 1476 333 1484
rect 627 1476 833 1484
rect 847 1476 1053 1484
rect 1467 1476 1513 1484
rect 1967 1476 2033 1484
rect 2047 1476 2113 1484
rect 2127 1476 2393 1484
rect 2487 1476 2513 1484
rect 2587 1476 2864 1484
rect 2856 1468 2864 1476
rect 2947 1476 3153 1484
rect 3247 1476 3373 1484
rect 4147 1476 4473 1484
rect 4887 1476 4973 1484
rect 5527 1476 5593 1484
rect 6147 1476 6213 1484
rect 6507 1476 6773 1484
rect 987 1456 1113 1464
rect 1347 1456 1433 1464
rect 1647 1456 1904 1464
rect 1896 1448 1904 1456
rect 2867 1457 2913 1465
rect 3207 1456 3253 1464
rect 3267 1456 3413 1464
rect 3467 1457 3493 1465
rect 4567 1456 4613 1464
rect 5136 1456 5173 1464
rect 127 1437 213 1445
rect 587 1436 693 1444
rect 707 1437 753 1445
rect 907 1436 933 1444
rect 947 1437 1013 1445
rect 1207 1437 1293 1445
rect 1827 1437 1853 1445
rect 1907 1437 1933 1445
rect 1073 1424 1087 1433
rect 1036 1420 1087 1424
rect 1036 1416 1084 1420
rect 87 1396 133 1404
rect 407 1396 593 1404
rect 787 1396 833 1404
rect 1036 1404 1044 1416
rect 927 1396 1044 1404
rect 1067 1395 1093 1403
rect 1187 1396 1273 1404
rect 1627 1396 1693 1404
rect 1707 1396 1793 1404
rect 2007 1395 2033 1403
rect 2136 1404 2144 1453
rect 2287 1437 2373 1445
rect 3127 1437 3173 1445
rect 3307 1437 3333 1445
rect 2156 1424 2164 1434
rect 3947 1436 4053 1444
rect 4247 1437 4293 1445
rect 4427 1437 4453 1445
rect 4587 1436 4653 1444
rect 4707 1437 4793 1445
rect 4807 1436 4824 1444
rect 2156 1420 2264 1424
rect 2156 1416 2267 1420
rect 2253 1407 2267 1416
rect 2887 1416 2953 1424
rect 3367 1416 3533 1424
rect 4816 1424 4824 1436
rect 4847 1436 4913 1444
rect 4987 1436 5013 1444
rect 5027 1437 5073 1445
rect 3667 1416 4064 1424
rect 4816 1416 5013 1424
rect 2136 1396 2164 1404
rect 2156 1384 2164 1396
rect 2307 1396 2353 1404
rect 2427 1396 2453 1404
rect 2987 1396 3093 1404
rect 3167 1396 3273 1404
rect 4007 1395 4033 1403
rect 4056 1404 4064 1416
rect 4056 1396 4213 1404
rect 4407 1396 4693 1404
rect 4787 1395 4833 1403
rect 4947 1395 4973 1403
rect 5136 1404 5144 1456
rect 5507 1457 5753 1465
rect 6367 1456 6433 1464
rect 5927 1436 6144 1444
rect 5167 1415 5253 1423
rect 5927 1416 6073 1424
rect 6136 1424 6144 1436
rect 6347 1436 6413 1444
rect 6427 1436 6513 1444
rect 6567 1436 6633 1444
rect 6687 1437 6813 1445
rect 6136 1416 6153 1424
rect 5136 1396 5233 1404
rect 6107 1396 6133 1404
rect 6447 1395 6473 1403
rect 6587 1395 6653 1403
rect 6727 1396 6793 1404
rect 2156 1376 2193 1384
rect 2247 1376 2273 1384
rect 3407 1376 3833 1384
rect 4607 1376 4873 1384
rect 5027 1376 5093 1384
rect 5667 1376 5793 1384
rect 787 1356 813 1364
rect 887 1356 953 1364
rect 1387 1356 1613 1364
rect 1867 1356 2133 1364
rect 2887 1356 4024 1364
rect 1507 1336 1953 1344
rect 2267 1336 2553 1344
rect 3187 1336 3893 1344
rect 4016 1344 4024 1356
rect 4987 1356 5073 1364
rect 6367 1356 6393 1364
rect 4016 1336 4453 1344
rect 4467 1336 4553 1344
rect 6667 1336 6933 1344
rect 707 1316 933 1324
rect 1147 1316 1413 1324
rect 2107 1316 2173 1324
rect 2407 1316 2633 1324
rect 2867 1316 2893 1324
rect 2967 1316 3033 1324
rect 3047 1316 3233 1324
rect 3527 1316 4133 1324
rect 5027 1316 5053 1324
rect 6627 1316 6853 1324
rect 467 1296 493 1304
rect 507 1296 553 1304
rect 2467 1296 2493 1304
rect 3347 1296 4232 1304
rect 4267 1296 4333 1304
rect 4347 1296 4433 1304
rect 4447 1296 4693 1304
rect 4767 1296 4933 1304
rect 5467 1296 5593 1304
rect 5827 1296 5953 1304
rect 6616 1304 6624 1313
rect 6067 1296 6624 1304
rect 147 1276 213 1284
rect 227 1276 393 1284
rect 407 1276 593 1284
rect 647 1276 1153 1284
rect 1707 1276 2113 1284
rect 2207 1276 2373 1284
rect 2527 1276 3513 1284
rect 3567 1276 3733 1284
rect 3747 1276 4993 1284
rect 5007 1276 5053 1284
rect 6107 1276 6273 1284
rect 267 1256 293 1264
rect 1727 1256 1993 1264
rect 2147 1256 2233 1264
rect 3007 1256 3053 1264
rect 3867 1256 4073 1264
rect 4307 1256 4553 1264
rect 4747 1256 4793 1264
rect 5147 1256 5593 1264
rect 6127 1256 6153 1264
rect 6327 1256 6393 1264
rect 6467 1256 6553 1264
rect 6567 1256 6673 1264
rect 547 1236 1093 1244
rect 1107 1236 1173 1244
rect 1827 1236 1873 1244
rect 2127 1236 2213 1244
rect 2227 1236 2513 1244
rect 6236 1236 6653 1244
rect 187 1216 233 1224
rect 367 1216 453 1224
rect 647 1217 673 1225
rect 1227 1216 1273 1224
rect 1436 1204 1444 1233
rect 1467 1217 1693 1225
rect 1196 1196 1304 1204
rect 1436 1196 1464 1204
rect 327 1175 353 1183
rect 407 1175 433 1183
rect 487 1175 553 1183
rect 567 1175 673 1183
rect 1196 1184 1204 1196
rect 1147 1176 1204 1184
rect 1296 1184 1304 1196
rect 1296 1176 1433 1184
rect 1456 1184 1464 1196
rect 1456 1176 1493 1184
rect 1756 1186 1764 1233
rect 6236 1228 6244 1236
rect 1787 1216 1953 1224
rect 2067 1216 2153 1224
rect 2267 1216 2333 1224
rect 2387 1217 2413 1225
rect 2687 1216 2733 1224
rect 2787 1217 2833 1225
rect 2947 1217 2993 1225
rect 3387 1216 3413 1224
rect 3427 1216 3793 1224
rect 4007 1217 4113 1225
rect 4207 1217 4273 1225
rect 4527 1217 4593 1225
rect 4687 1216 4753 1224
rect 4987 1216 5293 1224
rect 5307 1216 5333 1224
rect 5387 1217 5413 1225
rect 6507 1217 6553 1225
rect 6727 1217 6773 1225
rect 6827 1216 6873 1224
rect 5367 1197 5493 1205
rect 1647 1175 1713 1183
rect 2087 1175 2133 1183
rect 2187 1175 2233 1183
rect 2247 1176 2353 1184
rect 2816 1176 3013 1184
rect 127 1156 193 1164
rect 747 1156 853 1164
rect 1227 1156 1473 1164
rect 1567 1156 1593 1164
rect 2707 1156 2773 1164
rect 2816 1164 2824 1176
rect 3447 1176 3633 1184
rect 4107 1176 4193 1184
rect 4347 1175 4413 1183
rect 4627 1175 4673 1183
rect 5167 1176 5273 1184
rect 5607 1176 5733 1184
rect 6076 1184 6084 1213
rect 6687 1196 6804 1204
rect 6076 1176 6093 1184
rect 6347 1176 6473 1184
rect 6796 1186 6804 1196
rect 6567 1176 6613 1184
rect 6707 1175 6753 1183
rect 2787 1156 2824 1164
rect 4267 1156 4573 1164
rect 287 1136 613 1144
rect 947 1136 993 1144
rect 1596 1144 1604 1153
rect 1267 1136 1444 1144
rect 1596 1136 1833 1144
rect 627 1116 713 1124
rect 1436 1124 1444 1136
rect 2027 1136 2253 1144
rect 2587 1136 2893 1144
rect 3927 1136 4013 1144
rect 4256 1144 4264 1153
rect 4027 1136 4264 1144
rect 4307 1136 4513 1144
rect 5447 1136 5953 1144
rect 6207 1136 6713 1144
rect 1436 1116 1933 1124
rect 2016 1124 2024 1133
rect 1947 1116 2024 1124
rect 2547 1116 2973 1124
rect 2987 1116 3073 1124
rect 4687 1116 5373 1124
rect 6547 1116 6673 1124
rect 1087 1096 1133 1104
rect 1147 1096 1293 1104
rect 1427 1096 1493 1104
rect 1707 1096 1793 1104
rect 2027 1096 2313 1104
rect 2327 1096 2453 1104
rect 2467 1096 2513 1104
rect 2567 1096 2853 1104
rect 2907 1096 3433 1104
rect 3807 1096 4373 1104
rect 4667 1096 5113 1104
rect 6727 1096 6833 1104
rect 1207 1076 1313 1084
rect 3607 1076 4393 1084
rect 6227 1076 6853 1084
rect 2327 1056 2393 1064
rect 4147 1056 4733 1064
rect 5207 1056 5533 1064
rect 5807 1056 6513 1064
rect 527 1036 793 1044
rect 2007 1036 2933 1044
rect 3467 1036 3853 1044
rect 3867 1036 4093 1044
rect 4227 1036 4293 1044
rect 4507 1036 4913 1044
rect 6187 1036 6293 1044
rect 1647 1016 1893 1024
rect 1907 1016 2333 1024
rect 2427 1016 3504 1024
rect 2336 1004 2344 1013
rect 2336 996 2953 1004
rect 2967 996 3433 1004
rect 3496 1004 3504 1016
rect 3496 996 3693 1004
rect 3967 996 4213 1004
rect 4707 996 4773 1004
rect 5487 996 5873 1004
rect 6347 996 6413 1004
rect 687 976 793 984
rect 1827 976 2553 984
rect 3027 976 3293 984
rect 4007 976 4193 984
rect 4247 976 4673 984
rect 4867 976 5313 984
rect 5927 976 6053 984
rect 6127 976 6193 984
rect 6407 976 6753 984
rect 207 956 513 964
rect 1587 956 1653 964
rect 1667 956 1753 964
rect 2147 956 2453 964
rect 2467 956 2573 964
rect 2667 956 3373 964
rect 4047 956 4193 964
rect 4207 956 4533 964
rect 4767 956 5413 964
rect 5847 956 5893 964
rect 6467 956 6573 964
rect 6587 956 6644 964
rect 547 936 573 944
rect 6636 928 6644 956
rect 6667 936 6793 944
rect 147 917 213 925
rect 287 917 353 925
rect 447 917 473 925
rect 667 916 873 924
rect 1727 917 1833 925
rect 2187 917 2233 925
rect 207 876 273 884
rect 347 876 433 884
rect 687 876 752 884
rect 787 876 833 884
rect 907 876 1233 884
rect 1287 875 1353 883
rect 1536 884 1544 913
rect 1896 904 1904 914
rect 2487 916 2533 924
rect 2727 916 2813 924
rect 2867 916 3093 924
rect 3136 916 3153 924
rect 1836 896 1904 904
rect 1536 876 1553 884
rect 1836 884 1844 896
rect 1787 876 1844 884
rect 1867 876 1913 884
rect 2267 876 2313 884
rect 2587 875 2653 883
rect 2747 875 2792 883
rect 2827 875 2873 883
rect 2887 876 2973 884
rect 3136 884 3144 916
rect 3207 916 3413 924
rect 3567 917 3673 925
rect 3967 916 3993 924
rect 4167 917 4253 925
rect 4427 917 4473 925
rect 4527 916 4733 924
rect 4827 917 4873 925
rect 5407 917 5473 925
rect 5607 916 5813 924
rect 6167 917 6273 925
rect 6276 904 6284 914
rect 6276 896 6313 904
rect 3047 876 3144 884
rect 3487 875 3533 883
rect 3827 875 3853 883
rect 4247 875 4353 883
rect 4567 875 4633 883
rect 4787 875 4853 883
rect 5427 876 5493 884
rect 5787 876 5893 884
rect 6127 875 6173 883
rect 6187 876 6264 884
rect 6256 867 6264 876
rect 6367 875 6393 883
rect 6687 876 6773 884
rect 867 856 933 864
rect 2067 856 2213 864
rect 3007 856 3033 864
rect 3087 856 3133 864
rect 3387 856 3453 864
rect 4127 856 4193 864
rect 4447 856 4513 864
rect 5327 856 5393 864
rect 6256 856 6273 867
rect 6260 853 6273 856
rect 627 836 673 844
rect 807 836 1033 844
rect 1127 836 1453 844
rect 1647 836 1733 844
rect 1807 836 1893 844
rect 1907 836 2013 844
rect 2347 836 2393 844
rect 3287 836 3953 844
rect 4627 836 4673 844
rect 4800 844 4813 847
rect 4796 833 4813 844
rect 5427 836 5693 844
rect 5827 836 6033 844
rect 6827 836 6873 844
rect 1456 824 1464 833
rect 1456 816 1713 824
rect 1767 816 2093 824
rect 2107 816 2173 824
rect 2527 816 2693 824
rect 3447 816 3573 824
rect 3787 816 4413 824
rect 4427 816 4553 824
rect 4796 824 4804 833
rect 4727 816 4804 824
rect 4867 816 5013 824
rect 5247 816 5773 824
rect 167 796 453 804
rect 547 796 973 804
rect 987 796 1853 804
rect 1867 796 2053 804
rect 2727 796 3393 804
rect 4827 796 5193 804
rect 5347 796 5533 804
rect 5547 796 5633 804
rect 5927 796 6093 804
rect 6147 796 6173 804
rect 1067 776 1133 784
rect 1327 776 1433 784
rect 1447 776 1793 784
rect 1847 776 1953 784
rect 1967 776 1993 784
rect 2087 776 2133 784
rect 2227 776 2733 784
rect 2747 776 3193 784
rect 3867 776 4233 784
rect 4296 776 4433 784
rect 107 756 233 764
rect 4296 764 4304 776
rect 4527 776 4633 784
rect 4907 776 5093 784
rect 5247 776 5493 784
rect 3827 756 4304 764
rect 4327 756 4393 764
rect 647 736 733 744
rect 847 736 973 744
rect 1727 736 1773 744
rect 2347 736 2573 744
rect 2887 736 2933 744
rect 3067 736 3433 744
rect 3447 736 3593 744
rect 3847 736 4073 744
rect 4187 736 4213 744
rect 4227 736 4313 744
rect 4547 736 4613 744
rect 4627 736 5413 744
rect 5687 736 5833 744
rect 5887 736 6473 744
rect 127 716 153 724
rect 2007 716 2033 724
rect 3087 716 3113 724
rect 3647 716 3693 724
rect 4756 716 5233 724
rect 167 697 213 705
rect 307 696 553 704
rect 907 697 933 705
rect 987 696 1253 704
rect 1327 697 1413 705
rect 1507 696 1573 704
rect 1596 696 1833 704
rect 1596 666 1604 696
rect 2507 697 2533 705
rect 2627 697 2713 705
rect 2847 697 2913 705
rect 3727 697 3773 705
rect 3796 696 3833 704
rect 2247 675 2333 683
rect 3796 684 3804 696
rect 3887 696 3993 704
rect 4047 696 4113 704
rect 4367 697 4393 705
rect 4756 707 4764 716
rect 6247 716 6453 724
rect 4507 696 4573 704
rect 4587 696 4593 704
rect 4647 696 4753 704
rect 4996 696 5093 704
rect 4996 686 5004 696
rect 5267 697 5453 705
rect 5647 696 5773 704
rect 5847 697 5873 705
rect 6187 696 6213 704
rect 6527 697 6573 705
rect 3636 676 3804 684
rect 147 656 313 664
rect 487 656 613 664
rect 807 655 973 663
rect 1127 656 1233 664
rect 1247 656 1433 664
rect 1447 655 1493 663
rect 1647 655 1673 663
rect 1767 655 1853 663
rect 1907 656 1933 664
rect 2107 656 2553 664
rect 2567 655 2653 663
rect 2907 656 2993 664
rect 3087 655 3113 663
rect 3636 664 3644 676
rect 3627 656 3644 664
rect 3707 655 3753 663
rect 3907 655 3933 663
rect 4147 655 4173 663
rect 4227 655 4253 663
rect 4447 655 4513 663
rect 4627 655 4653 663
rect 5247 655 5333 663
rect 5487 656 5573 664
rect 6193 664 6207 673
rect 6047 660 6207 664
rect 6047 656 6204 660
rect 1287 636 1313 644
rect 2407 635 2473 643
rect 2627 636 2833 644
rect 5687 635 5873 643
rect 6587 636 6673 644
rect 207 616 973 624
rect 3267 616 4033 624
rect 5676 624 5684 632
rect 5167 616 5684 624
rect 6187 616 6273 624
rect 6727 616 6813 624
rect 3467 596 3893 604
rect 5767 596 6313 604
rect 2847 576 3653 584
rect 3667 576 4113 584
rect 4127 576 4693 584
rect 2467 556 2513 564
rect 2607 556 3253 564
rect 3567 556 3713 564
rect 3987 556 4493 564
rect 127 536 233 544
rect 1347 536 1493 544
rect 1687 536 2033 544
rect 2047 536 2273 544
rect 2287 536 2373 544
rect 3647 536 3873 544
rect 5267 536 5293 544
rect 6127 536 6393 544
rect 6587 536 6693 544
rect 6707 536 6793 544
rect 1547 516 2493 524
rect 2507 516 2573 524
rect 2767 516 3493 524
rect 5627 516 6033 524
rect 6047 516 6293 524
rect 287 496 453 504
rect 467 496 993 504
rect 1347 496 1833 504
rect 2756 504 2764 513
rect 2547 496 2764 504
rect 2947 496 3073 504
rect 3087 496 3273 504
rect 3496 504 3504 513
rect 3496 496 5013 504
rect 5787 496 5813 504
rect 6347 496 6473 504
rect 167 476 213 484
rect 227 476 2473 484
rect 2667 476 3213 484
rect 3387 476 3793 484
rect 6247 476 6793 484
rect 787 456 913 464
rect 927 456 953 464
rect 1007 456 1213 464
rect 1227 456 1353 464
rect 1367 456 1533 464
rect 2036 456 4053 464
rect 2036 447 2044 456
rect 4387 456 4873 464
rect 947 436 1713 444
rect 1727 436 2032 444
rect 2067 436 2133 444
rect 2147 436 2593 444
rect 2847 436 3293 444
rect 3447 436 3853 444
rect 3867 436 4653 444
rect 5067 436 5393 444
rect 5507 436 5553 444
rect 6227 436 6333 444
rect 6347 436 6493 444
rect 6787 436 6893 444
rect 567 416 633 424
rect 1147 416 1173 424
rect 1187 416 1333 424
rect 2476 416 2793 424
rect 507 396 593 404
rect 607 396 833 404
rect 987 397 1393 405
rect 1416 396 1433 404
rect 1416 384 1424 396
rect 1607 396 1673 404
rect 1907 396 2093 404
rect 2327 396 2433 404
rect 2476 404 2484 416
rect 2807 416 2853 424
rect 3627 416 3824 424
rect 2447 396 2484 404
rect 2547 397 2613 405
rect 2687 397 2773 405
rect 2787 396 2893 404
rect 3667 397 3793 405
rect 3816 404 3824 416
rect 5627 417 5673 425
rect 6187 416 6233 424
rect 6307 416 6353 424
rect 3816 396 3973 404
rect 4047 397 4153 405
rect 4247 397 4273 405
rect 4327 397 4353 405
rect 4407 397 4433 405
rect 4627 396 4673 404
rect 4767 396 4853 404
rect 4867 397 4953 405
rect 5047 396 5093 404
rect 6267 396 6313 404
rect 6327 397 6373 405
rect 6447 396 6513 404
rect 6647 397 6733 405
rect 1367 376 1424 384
rect 147 356 253 364
rect 527 356 553 364
rect 707 356 752 364
rect 787 355 813 363
rect 947 356 993 364
rect 1227 355 1253 363
rect 1307 355 1333 363
rect 1467 355 1512 363
rect 1547 356 1573 364
rect 1687 355 1753 363
rect 1847 355 1873 363
rect 2047 355 2073 363
rect 2167 355 2333 363
rect 2607 356 2693 364
rect 2767 356 2953 364
rect 2967 356 3033 364
rect 3347 356 3513 364
rect 3527 355 3633 363
rect 4067 355 4093 363
rect 4147 356 4233 364
rect 4307 356 4393 364
rect 4496 364 4504 393
rect 5527 375 5673 383
rect 4467 356 4504 364
rect 4707 355 4733 363
rect 4987 355 5033 363
rect 5127 356 5153 364
rect 5167 356 5253 364
rect 6127 356 6193 364
rect 6507 356 6713 364
rect 307 336 473 344
rect 487 336 573 344
rect 867 336 1033 344
rect 1047 336 1113 344
rect 2467 336 2533 344
rect 6167 336 6293 344
rect 6307 336 6373 344
rect 667 316 753 324
rect 1116 324 1124 333
rect 1116 316 1653 324
rect 1667 316 1713 324
rect 1727 316 2653 324
rect 2667 316 2813 324
rect 2927 316 3053 324
rect 3147 316 3373 324
rect 3787 316 3913 324
rect 4367 316 4593 324
rect 4607 316 5253 324
rect 5507 316 5653 324
rect 6567 316 6633 324
rect 6647 316 6713 324
rect 6927 316 6953 324
rect 647 296 733 304
rect 1427 296 1493 304
rect 1967 296 2833 304
rect 3567 296 3713 304
rect 3867 296 4033 304
rect 4667 296 4813 304
rect 4947 296 5053 304
rect 6367 296 6433 304
rect 2347 276 2693 284
rect 4887 276 5664 284
rect 1927 256 1993 264
rect 2307 256 2673 264
rect 2907 256 3153 264
rect 3167 256 3193 264
rect 4047 256 4613 264
rect 5656 264 5664 276
rect 6827 276 6913 284
rect 5656 256 5873 264
rect 6387 256 6553 264
rect 2447 236 2613 244
rect 2707 236 3453 244
rect 5227 236 5393 244
rect 5407 236 5953 244
rect 5967 236 6293 244
rect 167 216 313 224
rect 327 216 433 224
rect 447 216 1353 224
rect 2867 216 2953 224
rect 2967 216 3433 224
rect 3927 216 4473 224
rect 4527 216 4653 224
rect 4947 216 5053 224
rect 6367 216 6473 224
rect 567 196 733 204
rect 2467 196 2513 204
rect 3287 196 3513 204
rect 3527 196 3593 204
rect 4267 196 4373 204
rect 4647 196 4673 204
rect 4687 196 4713 204
rect 6787 196 6833 204
rect 707 176 793 184
rect 807 176 973 184
rect 1207 176 1273 184
rect 1287 177 1553 185
rect 2456 184 2464 193
rect 1727 176 2464 184
rect 2707 176 2793 184
rect 3227 176 3653 184
rect 3707 176 3793 184
rect 1907 155 1993 163
rect 2147 155 2273 163
rect 2487 157 2513 165
rect 3656 164 3664 174
rect 4087 177 4173 185
rect 4307 177 4333 185
rect 3996 164 4004 174
rect 3656 156 4004 164
rect 4036 164 4044 174
rect 4447 176 4533 184
rect 4627 176 4704 184
rect 4036 156 4284 164
rect -24 136 113 144
rect 367 135 553 143
rect 567 135 613 143
rect 667 135 693 143
rect 747 135 833 143
rect 927 135 953 143
rect 1447 136 1553 144
rect 2627 135 2673 143
rect 2727 135 2953 143
rect 3167 135 3193 143
rect 3407 136 3533 144
rect 3807 135 3833 143
rect 4027 136 4073 144
rect 4207 135 4253 143
rect 4276 144 4284 156
rect 4696 146 4704 176
rect 4807 176 4873 184
rect 5027 176 5173 184
rect 6427 176 6513 184
rect 6567 176 6673 184
rect 5707 156 5833 164
rect 6127 156 6144 164
rect 4276 136 4353 144
rect 4367 135 4433 143
rect 4487 135 4513 143
rect 4567 135 4633 143
rect 4747 135 4793 143
rect 4867 136 5073 144
rect 5087 136 5313 144
rect 6136 144 6144 156
rect 6407 156 6504 164
rect 6136 136 6413 144
rect 6496 146 6504 156
rect 6867 135 6933 143
rect 2067 116 2113 124
rect 2127 115 2413 123
rect 3607 116 3673 124
rect 4887 116 4933 124
rect 5687 116 5733 124
rect 3087 96 3233 104
rect 3247 96 3353 104
rect 3547 96 3693 104
rect 1387 76 2473 84
rect 3716 84 3724 113
rect 5747 116 5913 124
rect 5927 115 5953 123
rect 6267 116 6533 124
rect 3747 96 4153 104
rect 4407 96 4693 104
rect 4787 96 5573 104
rect 2807 76 4293 84
rect 5847 76 6013 84
rect 6027 76 6453 84
rect 2487 36 3613 44
rect 3627 36 4893 44
rect 4907 36 5033 44
use INVX1  _828_
timestamp 0
transform 1 0 890 0 1 5470
box -6 -8 46 268
use INVX1  _829_
timestamp 0
transform 1 0 1570 0 1 5470
box -6 -8 46 268
use NOR2X1  _830_
timestamp 0
transform -1 0 2470 0 1 5470
box -6 -8 66 268
use NAND3X1  _831_
timestamp 0
transform -1 0 1470 0 1 5470
box -6 -8 86 268
use INVX1  _832_
timestamp 0
transform 1 0 2330 0 1 5990
box -6 -8 46 268
use INVX1  _833_
timestamp 0
transform 1 0 2030 0 -1 5990
box -6 -8 46 268
use NOR2X1  _834_
timestamp 0
transform -1 0 1690 0 1 4950
box -6 -8 66 268
use NAND3X1  _835_
timestamp 0
transform -1 0 1790 0 1 5470
box -6 -8 86 268
use OAI22X1  _836_
timestamp 0
transform -1 0 1130 0 1 5470
box -6 -8 106 268
use NAND2X1  _837_
timestamp 0
transform 1 0 910 0 -1 5470
box -6 -8 66 268
use INVX1  _838_
timestamp 0
transform -1 0 790 0 -1 4950
box -6 -8 46 268
use OAI21X1  _839_
timestamp 0
transform -1 0 1030 0 1 4950
box -6 -8 86 268
use INVX1  _840_
timestamp 0
transform 1 0 110 0 -1 3390
box -6 -8 46 268
use NOR2X1  _841_
timestamp 0
transform -1 0 170 0 -1 2870
box -6 -8 66 268
use NAND3X1  _842_
timestamp 0
transform 1 0 110 0 -1 3910
box -6 -8 86 268
use OAI21X1  _843_
timestamp 0
transform -1 0 350 0 1 3910
box -6 -8 86 268
use INVX1  _844_
timestamp 0
transform 1 0 750 0 1 3390
box -6 -8 46 268
use AOI21X1  _845_
timestamp 0
transform 1 0 290 0 -1 3910
box -6 -8 86 268
use NOR2X1  _846_
timestamp 0
transform -1 0 850 0 -1 3910
box -6 -8 66 268
use NOR2X1  _847_
timestamp 0
transform -1 0 1010 0 -1 3910
box -6 -8 66 268
use AOI21X1  _848_
timestamp 0
transform -1 0 690 0 -1 3910
box -6 -8 86 268
use OAI21X1  _849_
timestamp 0
transform 1 0 270 0 -1 4430
box -6 -8 86 268
use NOR3X1  _850_
timestamp 0
transform -1 0 430 0 1 4950
box -6 -8 166 268
use NAND2X1  _851_
timestamp 0
transform -1 0 970 0 -1 5990
box -6 -8 66 268
use OR2X2  _852_
timestamp 0
transform -1 0 810 0 -1 5990
box -6 -8 86 268
use NOR2X1  _853_
timestamp 0
transform 1 0 630 0 1 5990
box -6 -8 66 268
use NOR2X1  _854_
timestamp 0
transform -1 0 170 0 -1 4430
box -6 -8 66 268
use NAND2X1  _855_
timestamp 0
transform -1 0 650 0 -1 4950
box -6 -8 66 268
use NOR2X1  _856_
timestamp 0
transform -1 0 850 0 1 4950
box -6 -8 66 268
use INVX2  _857_
timestamp 0
transform 1 0 1070 0 -1 5990
box -6 -8 46 268
use NOR3X1  _858_
timestamp 0
transform -1 0 690 0 1 4950
box -6 -8 166 268
use INVX8  _859_
timestamp 0
transform 1 0 110 0 1 5990
box -6 -8 106 268
use INVX1  _860_
timestamp 0
transform 1 0 1130 0 1 4950
box -6 -8 46 268
use NOR2X1  _861_
timestamp 0
transform 1 0 890 0 -1 4950
box -6 -8 66 268
use NAND3X1  _862_
timestamp 0
transform -1 0 830 0 -1 5470
box -6 -8 86 268
use OAI21X1  _863_
timestamp 0
transform -1 0 650 0 -1 5470
box -6 -8 86 268
use OAI21X1  _864_
timestamp 0
transform 1 0 890 0 1 4430
box -6 -8 86 268
use INVX1  _865_
timestamp 0
transform 1 0 470 0 -1 3910
box -6 -8 46 268
use INVX1  _866_
timestamp 0
transform -1 0 1450 0 1 4430
box -6 -8 46 268
use OAI21X1  _867_
timestamp 0
transform 1 0 1050 0 -1 4950
box -6 -8 86 268
use NAND3X1  _868_
timestamp 0
transform 1 0 1070 0 1 4430
box -6 -8 86 268
use NAND2X1  _869_
timestamp 0
transform -1 0 1310 0 1 4430
box -6 -8 66 268
use NOR2X1  _870_
timestamp 0
transform 1 0 1190 0 -1 4430
box -6 -8 66 268
use INVX2  _871_
timestamp 0
transform -1 0 1510 0 -1 3390
box -6 -8 46 268
use OAI21X1  _872_
timestamp 0
transform -1 0 990 0 1 3910
box -6 -8 86 268
use AOI21X1  _873_
timestamp 0
transform 1 0 1090 0 1 3910
box -6 -8 86 268
use INVX1  _874_
timestamp 0
transform 1 0 1070 0 1 3390
box -6 -8 46 268
use NOR2X1  _875_
timestamp 0
transform 1 0 1310 0 -1 3390
box -6 -8 66 268
use NAND2X1  _876_
timestamp 0
transform -1 0 1270 0 1 3390
box -6 -8 66 268
use OAI21X1  _877_
timestamp 0
transform 1 0 1370 0 1 3390
box -6 -8 86 268
use AOI21X1  _878_
timestamp 0
transform -1 0 970 0 1 3390
box -6 -8 86 268
use INVX1  _879_
timestamp 0
transform -1 0 150 0 1 2350
box -6 -8 46 268
use NAND2X1  _880_
timestamp 0
transform 1 0 1230 0 1 2870
box -6 -8 66 268
use OAI21X1  _881_
timestamp 0
transform 1 0 270 0 -1 2870
box -6 -8 86 268
use AOI21X1  _882_
timestamp 0
transform -1 0 330 0 1 2350
box -6 -8 86 268
use INVX1  _883_
timestamp 0
transform 1 0 910 0 -1 2870
box -6 -8 46 268
use OAI21X1  _884_
timestamp 0
transform -1 0 1130 0 1 2870
box -6 -8 86 268
use NOR3X1  _885_
timestamp 0
transform -1 0 1210 0 -1 3390
box -6 -8 166 268
use NOR2X1  _886_
timestamp 0
transform -1 0 950 0 1 2870
box -6 -8 66 268
use NAND2X1  _887_
timestamp 0
transform 1 0 910 0 -1 3390
box -6 -8 66 268
use NAND3X1  _888_
timestamp 0
transform -1 0 790 0 1 2870
box -6 -8 86 268
use INVX1  _889_
timestamp 0
transform 1 0 570 0 1 2870
box -6 -8 46 268
use NAND3X1  _890_
timestamp 0
transform -1 0 810 0 -1 3390
box -6 -8 86 268
use NAND2X1  _891_
timestamp 0
transform 1 0 390 0 -1 3390
box -6 -8 66 268
use NAND3X1  _892_
timestamp 0
transform -1 0 630 0 -1 3390
box -6 -8 86 268
use INVX1  _893_
timestamp 0
transform -1 0 290 0 -1 3390
box -6 -8 46 268
use AOI21X1  _894_
timestamp 0
transform -1 0 650 0 1 3390
box -6 -8 86 268
use NOR2X1  _895_
timestamp 0
transform -1 0 790 0 1 4430
box -6 -8 66 268
use INVX1  _896_
timestamp 0
transform 1 0 1870 0 -1 4950
box -6 -8 46 268
use INVX1  _897_
timestamp 0
transform -1 0 2610 0 1 5470
box -6 -8 46 268
use OAI21X1  _898_
timestamp 0
transform -1 0 2310 0 1 5470
box -6 -8 86 268
use NOR2X1  _899_
timestamp 0
transform 1 0 2190 0 -1 5470
box -6 -8 66 268
use AOI21X1  _900_
timestamp 0
transform -1 0 1870 0 1 4950
box -6 -8 86 268
use AOI21X1  _901_
timestamp 0
transform 1 0 1690 0 -1 4950
box -6 -8 86 268
use INVX1  _902_
timestamp 0
transform -1 0 1750 0 -1 5470
box -6 -8 46 268
use NAND2X1  _903_
timestamp 0
transform -1 0 1910 0 -1 5470
box -6 -8 66 268
use NAND3X1  _904_
timestamp 0
transform -1 0 1610 0 -1 5470
box -6 -8 86 268
use OAI21X1  _905_
timestamp 0
transform -1 0 1530 0 1 4950
box -6 -8 86 268
use OAI21X1  _906_
timestamp 0
transform 1 0 1270 0 1 4950
box -6 -8 86 268
use OAI21X1  _907_
timestamp 0
transform 1 0 1850 0 -1 5990
box -6 -8 86 268
use NAND3X1  _908_
timestamp 0
transform 1 0 2350 0 -1 5470
box -6 -8 86 268
use NAND2X1  _909_
timestamp 0
transform 1 0 2070 0 1 5470
box -6 -8 66 268
use NAND3X1  _910_
timestamp 0
transform -1 0 1970 0 1 5470
box -6 -8 86 268
use OAI21X1  _911_
timestamp 0
transform 1 0 1670 0 -1 5990
box -6 -8 86 268
use OAI21X1  _912_
timestamp 0
transform -1 0 1870 0 1 5990
box -6 -8 86 268
use INVX1  _913_
timestamp 0
transform 1 0 2910 0 1 5990
box -6 -8 46 268
use NAND2X1  _914_
timestamp 0
transform -1 0 3290 0 1 5990
box -6 -8 66 268
use OAI21X1  _915_
timestamp 0
transform 1 0 2170 0 -1 5990
box -6 -8 86 268
use NAND3X1  _916_
timestamp 0
transform -1 0 2230 0 1 5990
box -6 -8 86 268
use OAI21X1  _917_
timestamp 0
transform 1 0 1610 0 1 5990
box -6 -8 86 268
use OAI21X1  _918_
timestamp 0
transform 1 0 2010 0 -1 5470
box -6 -8 86 268
use NAND3X1  _919_
timestamp 0
transform -1 0 3130 0 1 5990
box -6 -8 86 268
use INVX1  _920_
timestamp 0
transform -1 0 3350 0 -1 6510
box -6 -8 46 268
use OAI21X1  _921_
timestamp 0
transform 1 0 2710 0 -1 5990
box -6 -8 86 268
use NAND3X1  _922_
timestamp 0
transform -1 0 2610 0 -1 5990
box -6 -8 86 268
use OAI21X1  _923_
timestamp 0
transform -1 0 2430 0 -1 5990
box -6 -8 86 268
use OAI21X1  _924_
timestamp 0
transform 1 0 1970 0 1 5990
box -6 -8 86 268
use NOR3X1  _925_
timestamp 0
transform 1 0 2650 0 1 5990
box -6 -8 166 268
use NAND2X1  _926_
timestamp 0
transform -1 0 2850 0 -1 6510
box -6 -8 66 268
use INVX1  _927_
timestamp 0
transform -1 0 3490 0 -1 6510
box -6 -8 46 268
use OAI21X1  _928_
timestamp 0
transform -1 0 3210 0 -1 6510
box -6 -8 86 268
use NAND3X1  _929_
timestamp 0
transform -1 0 2690 0 -1 6510
box -6 -8 86 268
use OAI21X1  _930_
timestamp 0
transform -1 0 2510 0 -1 6510
box -6 -8 86 268
use OAI21X1  _931_
timestamp 0
transform -1 0 1050 0 1 5990
box -6 -8 86 268
use NAND3X1  _932_
timestamp 0
transform -1 0 3030 0 -1 6510
box -6 -8 86 268
use OAI21X1  _933_
timestamp 0
transform -1 0 2950 0 -1 5990
box -6 -8 86 268
use NAND3X1  _934_
timestamp 0
transform -1 0 2550 0 1 5990
box -6 -8 86 268
use OAI21X1  _935_
timestamp 0
transform -1 0 870 0 1 5990
box -6 -8 86 268
use NOR2X1  _936_
timestamp 0
transform -1 0 1290 0 1 5470
box -6 -8 66 268
use NOR2X1  _937_
timestamp 0
transform -1 0 790 0 1 5470
box -6 -8 66 268
use DFFSR  _938_
timestamp 0
transform 1 0 170 0 -1 5990
box -6 -8 466 268
use DFFSR  _939_
timestamp 0
transform 1 0 10 0 -1 5470
box -6 -8 466 268
use DFFSR  _940_
timestamp 0
transform 1 0 630 0 -1 4430
box -6 -8 466 268
use DFFSR  _941_
timestamp 0
transform 1 0 1010 0 -1 3910
box -6 -8 466 268
use DFFSR  _942_
timestamp 0
transform 1 0 10 0 1 3390
box -6 -8 466 268
use DFFSR  _943_
timestamp 0
transform 1 0 10 0 -1 2350
box -6 -8 466 268
use DFFSR  _944_
timestamp 0
transform 1 0 350 0 -1 2870
box -6 -8 466 268
use DFFSR  _945_
timestamp 0
transform 1 0 10 0 1 2870
box -6 -8 466 268
use DFFSR  _946_
timestamp 0
transform 1 0 350 0 1 3910
box -6 -8 466 268
use DFFSR  _947_
timestamp 0
transform 1 0 170 0 1 4430
box -6 -8 466 268
use DFFSR  _948_
timestamp 0
transform 1 0 1130 0 -1 4950
box -6 -8 466 268
use DFFSR  _949_
timestamp 0
transform 1 0 970 0 -1 5470
box -6 -8 466 268
use DFFSR  _950_
timestamp 0
transform 1 0 1410 0 -1 6510
box -6 -8 466 268
use DFFSR  _951_
timestamp 0
transform 1 0 1050 0 1 5990
box -6 -8 466 268
use DFFSR  _952_
timestamp 0
transform 1 0 950 0 -1 6510
box -6 -8 466 268
use DFFSR  _953_
timestamp 0
transform 1 0 1870 0 -1 6510
box -6 -8 466 268
use DFFSR  _954_
timestamp 0
transform 1 0 490 0 -1 6510
box -6 -8 466 268
use DFFSR  _955_
timestamp 0
transform 1 0 1110 0 -1 5990
box -6 -8 466 268
use DFFSR  _956_
timestamp 0
transform 1 0 170 0 1 5470
box -6 -8 466 268
use INVX1  _957_
timestamp 0
transform 1 0 1890 0 -1 2870
box -6 -8 46 268
use INVX1  _958_
timestamp 0
transform -1 0 1310 0 1 2350
box -6 -8 46 268
use NOR2X1  _959_
timestamp 0
transform -1 0 1790 0 -1 2870
box -6 -8 66 268
use NAND3X1  _960_
timestamp 0
transform 1 0 1550 0 -1 2870
box -6 -8 86 268
use NOR2X1  _961_
timestamp 0
transform 1 0 1050 0 -1 2870
box -6 -8 66 268
use NOR2X1  _962_
timestamp 0
transform -1 0 490 0 1 2350
box -6 -8 66 268
use NAND2X1  _963_
timestamp 0
transform -1 0 1270 0 -1 2870
box -6 -8 66 268
use INVX2  _964_
timestamp 0
transform 1 0 2110 0 -1 3390
box -6 -8 46 268
use OAI21X1  _965_
timestamp 0
transform 1 0 1590 0 1 2870
box -6 -8 86 268
use NOR2X1  _966_
timestamp 0
transform 1 0 1770 0 1 2870
box -6 -8 66 268
use NAND2X1  _967_
timestamp 0
transform 1 0 1610 0 -1 3390
box -6 -8 66 268
use INVX1  _968_
timestamp 0
transform -1 0 3090 0 -1 5990
box -6 -8 46 268
use NOR2X1  _969_
timestamp 0
transform -1 0 6170 0 -1 4430
box -6 -8 66 268
use NOR2X1  _970_
timestamp 0
transform -1 0 6490 0 1 4430
box -6 -8 66 268
use NAND2X1  _971_
timestamp 0
transform 1 0 5950 0 -1 4430
box -6 -8 66 268
use AOI21X1  _972_
timestamp 0
transform -1 0 5850 0 -1 4430
box -6 -8 86 268
use XOR2X1  _973_
timestamp 0
transform 1 0 5450 0 -1 3910
box -6 -8 126 268
use NAND2X1  _974_
timestamp 0
transform 1 0 3290 0 1 3910
box -6 -8 66 268
use INVX1  _975_
timestamp 0
transform 1 0 2970 0 1 3910
box -6 -8 46 268
use INVX2  _976_
timestamp 0
transform -1 0 6590 0 -1 1830
box -6 -8 46 268
use NAND2X1  _977_
timestamp 0
transform 1 0 5810 0 1 3390
box -6 -8 66 268
use NOR2X1  _978_
timestamp 0
transform 1 0 5650 0 1 3390
box -6 -8 66 268
use AOI21X1  _979_
timestamp 0
transform -1 0 5550 0 1 3390
box -6 -8 86 268
use NOR2X1  _980_
timestamp 0
transform 1 0 5310 0 1 3390
box -6 -8 66 268
use NOR2X1  _981_
timestamp 0
transform 1 0 3550 0 -1 3910
box -6 -8 66 268
use INVX1  _982_
timestamp 0
transform -1 0 3590 0 -1 5470
box -6 -8 46 268
use INVX2  _983_
timestamp 0
transform -1 0 5390 0 -1 2870
box -6 -8 46 268
use NAND2X1  _984_
timestamp 0
transform 1 0 3950 0 1 4430
box -6 -8 66 268
use NAND3X1  _985_
timestamp 0
transform -1 0 4230 0 -1 4430
box -6 -8 86 268
use INVX1  _986_
timestamp 0
transform -1 0 3330 0 1 4430
box -6 -8 46 268
use NAND2X1  _987_
timestamp 0
transform -1 0 4050 0 -1 4430
box -6 -8 66 268
use INVX1  _988_
timestamp 0
transform 1 0 3690 0 -1 4430
box -6 -8 46 268
use NOR2X1  _989_
timestamp 0
transform -1 0 4570 0 -1 4430
box -6 -8 66 268
use INVX2  _990_
timestamp 0
transform 1 0 2950 0 -1 4950
box -6 -8 46 268
use INVX2  _991_
timestamp 0
transform -1 0 6430 0 1 790
box -6 -8 46 268
use NAND2X1  _992_
timestamp 0
transform -1 0 6330 0 -1 4430
box -6 -8 66 268
use OAI21X1  _993_
timestamp 0
transform 1 0 6050 0 1 3910
box -6 -8 86 268
use NAND2X1  _994_
timestamp 0
transform 1 0 6230 0 1 3910
box -6 -8 66 268
use NOR2X1  _995_
timestamp 0
transform 1 0 4270 0 1 3910
box -6 -8 66 268
use AOI21X1  _996_
timestamp 0
transform 1 0 4330 0 -1 4430
box -6 -8 86 268
use NAND2X1  _997_
timestamp 0
transform -1 0 4350 0 1 4430
box -6 -8 66 268
use INVX2  _998_
timestamp 0
transform 1 0 5610 0 -1 790
box -6 -8 46 268
use INVX2  _999_
timestamp 0
transform 1 0 6110 0 1 2350
box -6 -8 46 268
use NAND2X1  _1000_
timestamp 0
transform -1 0 6910 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1001_
timestamp 0
transform -1 0 6110 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1002_
timestamp 0
transform -1 0 5950 0 1 3910
box -6 -8 86 268
use NAND2X1  _1003_
timestamp 0
transform -1 0 5770 0 1 3910
box -6 -8 66 268
use OAI21X1  _1004_
timestamp 0
transform -1 0 4890 0 1 4430
box -6 -8 86 268
use INVX2  _1005_
timestamp 0
transform 1 0 6050 0 1 4950
box -6 -8 46 268
use AOI21X1  _1006_
timestamp 0
transform -1 0 5670 0 -1 4430
box -6 -8 86 268
use INVX1  _1007_
timestamp 0
transform -1 0 5550 0 1 4430
box -6 -8 46 268
use NAND3X1  _1008_
timestamp 0
transform -1 0 5890 0 1 4430
box -6 -8 86 268
use NAND2X1  _1009_
timestamp 0
transform -1 0 5710 0 1 4430
box -6 -8 66 268
use AOI22X1  _1010_
timestamp 0
transform -1 0 5270 0 1 4430
box -6 -8 106 268
use OAI21X1  _1011_
timestamp 0
transform 1 0 4990 0 1 4430
box -6 -8 86 268
use INVX1  _1012_
timestamp 0
transform 1 0 4750 0 -1 6510
box -6 -8 46 268
use INVX1  _1013_
timestamp 0
transform 1 0 4910 0 1 5990
box -6 -8 46 268
use INVX1  _1014_
timestamp 0
transform -1 0 5410 0 1 4430
box -6 -8 46 268
use NOR2X1  _1015_
timestamp 0
transform -1 0 5610 0 1 3910
box -6 -8 66 268
use NOR2X1  _1016_
timestamp 0
transform 1 0 5430 0 -1 4430
box -6 -8 66 268
use AOI22X1  _1017_
timestamp 0
transform -1 0 4930 0 -1 4430
box -6 -8 106 268
use NAND2X1  _1018_
timestamp 0
transform -1 0 4730 0 -1 4430
box -6 -8 66 268
use INVX1  _1019_
timestamp 0
transform -1 0 5350 0 -1 3910
box -6 -8 46 268
use OR2X2  _1020_
timestamp 0
transform -1 0 5290 0 1 3910
box -6 -8 86 268
use AOI22X1  _1021_
timestamp 0
transform -1 0 4030 0 1 3910
box -6 -8 106 268
use NAND2X1  _1022_
timestamp 0
transform 1 0 3770 0 1 3910
box -6 -8 66 268
use AOI21X1  _1023_
timestamp 0
transform -1 0 3110 0 -1 3910
box -6 -8 86 268
use INVX2  _1024_
timestamp 0
transform -1 0 2750 0 1 5470
box -6 -8 46 268
use XOR2X1  _1025_
timestamp 0
transform -1 0 4230 0 1 3390
box -6 -8 126 268
use AOI22X1  _1026_
timestamp 0
transform 1 0 3710 0 -1 3910
box -6 -8 106 268
use INVX1  _1027_
timestamp 0
transform 1 0 2970 0 1 3390
box -6 -8 46 268
use INVX2  _1028_
timestamp 0
transform 1 0 6330 0 -1 3390
box -6 -8 46 268
use XOR2X1  _1029_
timestamp 0
transform 1 0 4910 0 1 3390
box -6 -8 126 268
use NOR2X1  _1030_
timestamp 0
transform 1 0 3830 0 -1 5470
box -6 -8 66 268
use INVX1  _1031_
timestamp 0
transform -1 0 6950 0 -1 5470
box -6 -8 46 268
use NOR2X1  _1032_
timestamp 0
transform 1 0 4630 0 1 4950
box -6 -8 66 268
use NOR2X1  _1033_
timestamp 0
transform 1 0 4130 0 1 4950
box -6 -8 66 268
use NAND2X1  _1034_
timestamp 0
transform 1 0 3930 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1035_
timestamp 0
transform -1 0 4530 0 1 4950
box -6 -8 66 268
use NAND3X1  _1036_
timestamp 0
transform -1 0 4370 0 1 4950
box -6 -8 86 268
use INVX2  _1037_
timestamp 0
transform 1 0 6450 0 -1 6510
box -6 -8 46 268
use NAND2X1  _1038_
timestamp 0
transform 1 0 3990 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1039_
timestamp 0
transform -1 0 4630 0 1 5470
box -6 -8 66 268
use NOR2X1  _1040_
timestamp 0
transform -1 0 4790 0 1 5470
box -6 -8 66 268
use NOR2X1  _1041_
timestamp 0
transform 1 0 4070 0 1 5470
box -6 -8 66 268
use NOR2X1  _1042_
timestamp 0
transform -1 0 4290 0 1 5470
box -6 -8 66 268
use NAND3X1  _1043_
timestamp 0
transform -1 0 4470 0 1 5470
box -6 -8 86 268
use NOR2X1  _1044_
timestamp 0
transform 1 0 3770 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1045_
timestamp 0
transform -1 0 4530 0 1 4430
box -6 -8 86 268
use INVX1  _1046_
timestamp 0
transform -1 0 2690 0 -1 4950
box -6 -8 46 268
use OAI22X1  _1047_
timestamp 0
transform 1 0 4270 0 -1 4950
box -6 -8 106 268
use OR2X2  _1048_
timestamp 0
transform -1 0 4170 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1049_
timestamp 0
transform -1 0 3890 0 -1 4430
box -6 -8 66 268
use AOI21X1  _1050_
timestamp 0
transform 1 0 3350 0 -1 4430
box -6 -8 86 268
use NOR2X1  _1051_
timestamp 0
transform -1 0 3590 0 -1 4430
box -6 -8 66 268
use AOI21X1  _1052_
timestamp 0
transform -1 0 4710 0 1 4430
box -6 -8 86 268
use AOI21X1  _1053_
timestamp 0
transform -1 0 4190 0 1 4430
box -6 -8 86 268
use OAI21X1  _1054_
timestamp 0
transform 1 0 3770 0 1 4430
box -6 -8 86 268
use AOI21X1  _1055_
timestamp 0
transform -1 0 3970 0 1 5470
box -6 -8 86 268
use AOI21X1  _1056_
timestamp 0
transform -1 0 4030 0 1 4950
box -6 -8 86 268
use OAI21X1  _1057_
timestamp 0
transform 1 0 3770 0 1 4950
box -6 -8 86 268
use AOI21X1  _1058_
timestamp 0
transform -1 0 3670 0 1 4430
box -6 -8 86 268
use OAI21X1  _1059_
timestamp 0
transform -1 0 3190 0 1 3910
box -6 -8 86 268
use NOR2X1  _1060_
timestamp 0
transform 1 0 3450 0 1 3910
box -6 -8 66 268
use NAND2X1  _1061_
timestamp 0
transform -1 0 3670 0 1 3910
box -6 -8 66 268
use OAI21X1  _1062_
timestamp 0
transform -1 0 3550 0 1 3390
box -6 -8 86 268
use NOR2X1  _1063_
timestamp 0
transform 1 0 590 0 1 2350
box -6 -8 66 268
use NAND3X1  _1064_
timestamp 0
transform 1 0 750 0 1 2350
box -6 -8 86 268
use INVX1  _1065_
timestamp 0
transform 1 0 1150 0 -1 2350
box -6 -8 46 268
use INVX1  _1066_
timestamp 0
transform 1 0 850 0 -1 2350
box -6 -8 46 268
use NOR2X1  _1067_
timestamp 0
transform -1 0 1050 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1068_
timestamp 0
transform -1 0 1170 0 1 2350
box -6 -8 86 268
use NOR2X1  _1069_
timestamp 0
transform -1 0 990 0 1 2350
box -6 -8 66 268
use OAI21X1  _1070_
timestamp 0
transform -1 0 1450 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1071_
timestamp 0
transform 1 0 2470 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1072_
timestamp 0
transform -1 0 3370 0 1 3390
box -6 -8 86 268
use AOI21X1  _1073_
timestamp 0
transform -1 0 3190 0 1 3390
box -6 -8 86 268
use OAI21X1  _1074_
timestamp 0
transform -1 0 2870 0 1 3390
box -6 -8 86 268
use NAND3X1  _1075_
timestamp 0
transform 1 0 1550 0 1 3390
box -6 -8 86 268
use INVX1  _1076_
timestamp 0
transform -1 0 1470 0 -1 270
box -6 -8 46 268
use INVX1  _1077_
timestamp 0
transform 1 0 1270 0 1 3910
box -6 -8 46 268
use AND2X2  _1078_
timestamp 0
transform -1 0 3290 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1079_
timestamp 0
transform -1 0 2930 0 -1 3910
box -6 -8 86 268
use AOI22X1  _1080_
timestamp 0
transform 1 0 1890 0 1 3390
box -6 -8 106 268
use INVX2  _1081_
timestamp 0
transform -1 0 2770 0 -1 790
box -6 -8 46 268
use INVX2  _1082_
timestamp 0
transform 1 0 1930 0 -1 790
box -6 -8 46 268
use INVX2  _1083_
timestamp 0
transform -1 0 2430 0 1 790
box -6 -8 46 268
use NOR2X1  _1084_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 66 268
use AOI21X1  _1085_
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 86 268
use INVX1  _1086_
timestamp 0
transform 1 0 1110 0 1 270
box -6 -8 46 268
use INVX2  _1087_
timestamp 0
transform -1 0 1610 0 1 270
box -6 -8 46 268
use NOR2X1  _1088_
timestamp 0
transform -1 0 1310 0 1 270
box -6 -8 66 268
use NAND3X1  _1089_
timestamp 0
transform 1 0 1390 0 -1 790
box -6 -8 86 268
use XOR2X1  _1090_
timestamp 0
transform -1 0 1110 0 1 790
box -6 -8 126 268
use NAND2X1  _1091_
timestamp 0
transform 1 0 470 0 -1 1830
box -6 -8 66 268
use INVX2  _1092_
timestamp 0
transform 1 0 110 0 -1 1310
box -6 -8 46 268
use INVX1  _1093_
timestamp 0
transform -1 0 470 0 1 1310
box -6 -8 46 268
use NAND2X1  _1094_
timestamp 0
transform 1 0 110 0 1 1310
box -6 -8 66 268
use INVX2  _1095_
timestamp 0
transform 1 0 970 0 1 270
box -6 -8 46 268
use NAND2X1  _1096_
timestamp 0
transform -1 0 1290 0 -1 790
box -6 -8 66 268
use XOR2X1  _1097_
timestamp 0
transform 1 0 790 0 -1 790
box -6 -8 126 268
use XOR2X1  _1098_
timestamp 0
transform -1 0 230 0 -1 1830
box -6 -8 126 268
use AOI21X1  _1099_
timestamp 0
transform 1 0 110 0 1 1830
box -6 -8 86 268
use INVX1  _1100_
timestamp 0
transform -1 0 1990 0 -1 1830
box -6 -8 46 268
use INVX1  _1101_
timestamp 0
transform -1 0 2530 0 -1 1310
box -6 -8 46 268
use NAND2X1  _1102_
timestamp 0
transform 1 0 2110 0 1 1310
box -6 -8 66 268
use OAI21X1  _1103_
timestamp 0
transform -1 0 2390 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1104_
timestamp 0
transform -1 0 1290 0 1 790
box -6 -8 86 268
use AND2X2  _1105_
timestamp 0
transform -1 0 890 0 1 790
box -6 -8 86 268
use NAND2X1  _1106_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 66 268
use XOR2X1  _1107_
timestamp 0
transform -1 0 1130 0 -1 790
box -6 -8 126 268
use OR2X2  _1108_
timestamp 0
transform 1 0 1070 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1109_
timestamp 0
transform -1 0 710 0 1 790
box -6 -8 66 268
use NAND2X1  _1110_
timestamp 0
transform -1 0 810 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1111_
timestamp 0
transform -1 0 810 0 1 1310
box -6 -8 66 268
use OAI21X1  _1112_
timestamp 0
transform -1 0 650 0 1 1310
box -6 -8 86 268
use NOR2X1  _1113_
timestamp 0
transform 1 0 590 0 -1 1310
box -6 -8 66 268
use INVX1  _1114_
timestamp 0
transform -1 0 370 0 -1 1830
box -6 -8 46 268
use NAND2X1  _1115_
timestamp 0
transform -1 0 330 0 1 1310
box -6 -8 66 268
use NAND2X1  _1116_
timestamp 0
transform 1 0 430 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1117_
timestamp 0
transform 1 0 250 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1118_
timestamp 0
transform 1 0 290 0 1 1830
box -6 -8 86 268
use OAI21X1  _1119_
timestamp 0
transform 1 0 2210 0 1 790
box -6 -8 86 268
use INVX1  _1120_
timestamp 0
transform -1 0 2390 0 1 1830
box -6 -8 46 268
use NOR2X1  _1121_
timestamp 0
transform 1 0 2050 0 1 790
box -6 -8 66 268
use NAND2X1  _1122_
timestamp 0
transform -1 0 2490 0 1 1310
box -6 -8 66 268
use NAND2X1  _1123_
timestamp 0
transform 1 0 2270 0 1 1310
box -6 -8 66 268
use NAND3X1  _1124_
timestamp 0
transform 1 0 1710 0 1 790
box -6 -8 86 268
use NAND2X1  _1125_
timestamp 0
transform 1 0 1890 0 1 790
box -6 -8 66 268
use NOR2X1  _1126_
timestamp 0
transform 1 0 1790 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1127_
timestamp 0
transform 1 0 1610 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1128_
timestamp 0
transform 1 0 1550 0 1 2350
box -6 -8 86 268
use NAND2X1  _1129_
timestamp 0
transform 1 0 1590 0 1 1310
box -6 -8 66 268
use NAND3X1  _1130_
timestamp 0
transform -1 0 1830 0 1 1310
box -6 -8 86 268
use NAND2X1  _1131_
timestamp 0
transform -1 0 2150 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1132_
timestamp 0
transform -1 0 2210 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1133_
timestamp 0
transform -1 0 2030 0 -1 1310
box -6 -8 86 268
use AOI22X1  _1134_
timestamp 0
transform -1 0 1850 0 -1 1310
box -6 -8 106 268
use NAND2X1  _1135_
timestamp 0
transform 1 0 1250 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1136_
timestamp 0
transform -1 0 1490 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1137_
timestamp 0
transform -1 0 1150 0 1 1310
box -6 -8 66 268
use AOI22X1  _1138_
timestamp 0
transform -1 0 730 0 1 1830
box -6 -8 106 268
use NAND2X1  _1139_
timestamp 0
transform -1 0 530 0 1 1830
box -6 -8 66 268
use INVX2  _1140_
timestamp 0
transform -1 0 3950 0 -1 3910
box -6 -8 46 268
use INVX2  _1141_
timestamp 0
transform 1 0 4130 0 1 3910
box -6 -8 46 268
use INVX2  _1142_
timestamp 0
transform -1 0 4690 0 -1 2870
box -6 -8 46 268
use INVX1  _1143_
timestamp 0
transform 1 0 5570 0 -1 3390
box -6 -8 46 268
use NOR2X1  _1144_
timestamp 0
transform 1 0 6590 0 1 4430
box -6 -8 66 268
use AOI21X1  _1145_
timestamp 0
transform -1 0 5630 0 1 4950
box -6 -8 86 268
use AND2X2  _1146_
timestamp 0
transform 1 0 4850 0 -1 5470
box -6 -8 86 268
use NAND3X1  _1147_
timestamp 0
transform -1 0 5110 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1148_
timestamp 0
transform -1 0 4750 0 -1 5470
box -6 -8 86 268
use INVX2  _1149_
timestamp 0
transform 1 0 5730 0 1 4950
box -6 -8 46 268
use NOR2X1  _1150_
timestamp 0
transform -1 0 5290 0 1 4950
box -6 -8 66 268
use NAND3X1  _1151_
timestamp 0
transform -1 0 5290 0 -1 5470
box -6 -8 86 268
use OR2X2  _1152_
timestamp 0
transform -1 0 4570 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1153_
timestamp 0
transform -1 0 4390 0 -1 5470
box -6 -8 66 268
use INVX2  _1154_
timestamp 0
transform -1 0 6430 0 1 3910
box -6 -8 46 268
use INVX2  _1155_
timestamp 0
transform -1 0 6850 0 -1 3390
box -6 -8 46 268
use NAND2X1  _1156_
timestamp 0
transform 1 0 3270 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1157_
timestamp 0
transform 1 0 3590 0 -1 4950
box -6 -8 86 268
use NOR3X1  _1158_
timestamp 0
transform -1 0 6330 0 1 4430
box -6 -8 166 268
use NAND2X1  _1159_
timestamp 0
transform 1 0 5390 0 1 4950
box -6 -8 66 268
use NAND2X1  _1160_
timestamp 0
transform 1 0 5310 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1161_
timestamp 0
transform 1 0 4250 0 -1 6510
box -6 -8 66 268
use INVX2  _1162_
timestamp 0
transform -1 0 5130 0 1 4950
box -6 -8 46 268
use NOR3X1  _1163_
timestamp 0
transform 1 0 4890 0 1 5470
box -6 -8 166 268
use NAND3X1  _1164_
timestamp 0
transform 1 0 5130 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1165_
timestamp 0
transform 1 0 5150 0 1 5470
box -6 -8 86 268
use OAI21X1  _1166_
timestamp 0
transform -1 0 4970 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1167_
timestamp 0
transform -1 0 6070 0 1 4430
box -6 -8 86 268
use AND2X2  _1168_
timestamp 0
transform 1 0 5870 0 1 4950
box -6 -8 86 268
use NOR2X1  _1169_
timestamp 0
transform 1 0 3910 0 -1 6510
box -6 -8 66 268
use NAND2X1  _1170_
timestamp 0
transform 1 0 3190 0 -1 4430
box -6 -8 66 268
use NOR2X1  _1171_
timestamp 0
transform 1 0 2950 0 1 4430
box -6 -8 66 268
use OAI21X1  _1172_
timestamp 0
transform -1 0 3190 0 1 4430
box -6 -8 86 268
use NAND3X1  _1173_
timestamp 0
transform 1 0 3090 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1174_
timestamp 0
transform 1 0 3590 0 -1 6510
box -6 -8 66 268
use AOI21X1  _1175_
timestamp 0
transform 1 0 3730 0 -1 6510
box -6 -8 86 268
use OAI21X1  _1176_
timestamp 0
transform -1 0 4150 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1177_
timestamp 0
transform 1 0 4410 0 -1 6510
box -6 -8 86 268
use NOR2X1  _1178_
timestamp 0
transform -1 0 5130 0 -1 6510
box -6 -8 66 268
use NAND3X1  _1179_
timestamp 0
transform 1 0 5390 0 -1 5470
box -6 -8 86 268
use INVX2  _1180_
timestamp 0
transform 1 0 4790 0 1 4950
box -6 -8 46 268
use NAND3X1  _1181_
timestamp 0
transform 1 0 5330 0 1 5470
box -6 -8 86 268
use NAND2X1  _1182_
timestamp 0
transform 1 0 5230 0 1 5990
box -6 -8 66 268
use AND2X2  _1183_
timestamp 0
transform -1 0 5510 0 -1 6510
box -6 -8 86 268
use AOI22X1  _1184_
timestamp 0
transform 1 0 5230 0 -1 6510
box -6 -8 106 268
use NAND2X1  _1185_
timestamp 0
transform -1 0 4650 0 -1 6510
box -6 -8 66 268
use NAND2X1  _1186_
timestamp 0
transform -1 0 5670 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1187_
timestamp 0
transform -1 0 5270 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1188_
timestamp 0
transform -1 0 4910 0 -1 5990
box -6 -8 66 268
use AOI22X1  _1189_
timestamp 0
transform -1 0 4650 0 1 5990
box -6 -8 106 268
use OAI21X1  _1190_
timestamp 0
transform 1 0 5750 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1191_
timestamp 0
transform 1 0 6210 0 1 5470
box -6 -8 66 268
use OAI22X1  _1192_
timestamp 0
transform 1 0 4330 0 -1 5990
box -6 -8 106 268
use AOI21X1  _1193_
timestamp 0
transform -1 0 4450 0 1 5990
box -6 -8 86 268
use INVX1  _1194_
timestamp 0
transform -1 0 3730 0 -1 5470
box -6 -8 46 268
use NAND2X1  _1195_
timestamp 0
transform 1 0 3730 0 1 5470
box -6 -8 66 268
use OAI21X1  _1196_
timestamp 0
transform 1 0 3550 0 1 5470
box -6 -8 86 268
use OAI22X1  _1197_
timestamp 0
transform 1 0 3190 0 1 5470
box -6 -8 106 268
use NOR2X1  _1198_
timestamp 0
transform 1 0 3450 0 1 4950
box -6 -8 66 268
use NOR2X1  _1199_
timestamp 0
transform -1 0 3490 0 1 4430
box -6 -8 66 268
use OR2X2  _1200_
timestamp 0
transform -1 0 2330 0 1 4950
box -6 -8 86 268
use NOR2X1  _1201_
timestamp 0
transform 1 0 3610 0 1 4950
box -6 -8 66 268
use NOR2X1  _1202_
timestamp 0
transform 1 0 3430 0 -1 4950
box -6 -8 66 268
use OR2X2  _1203_
timestamp 0
transform -1 0 3350 0 1 4950
box -6 -8 86 268
use OR2X2  _1204_
timestamp 0
transform 1 0 2590 0 1 4950
box -6 -8 86 268
use NAND2X1  _1205_
timestamp 0
transform 1 0 2490 0 -1 4950
box -6 -8 66 268
use INVX1  _1206_
timestamp 0
transform 1 0 2170 0 -1 4950
box -6 -8 46 268
use NAND2X1  _1207_
timestamp 0
transform 1 0 2790 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1208_
timestamp 0
transform 1 0 2310 0 -1 4950
box -6 -8 86 268
use INVX1  _1209_
timestamp 0
transform -1 0 3170 0 1 4950
box -6 -8 46 268
use AOI21X1  _1210_
timestamp 0
transform -1 0 3030 0 1 4950
box -6 -8 86 268
use OAI21X1  _1211_
timestamp 0
transform 1 0 2770 0 1 4950
box -6 -8 86 268
use NOR2X1  _1212_
timestamp 0
transform 1 0 4530 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1213_
timestamp 0
transform 1 0 4690 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1214_
timestamp 0
transform 1 0 4170 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1215_
timestamp 0
transform -1 0 4110 0 1 5990
box -6 -8 66 268
use NOR2X1  _1216_
timestamp 0
transform 1 0 4750 0 1 5990
box -6 -8 66 268
use NOR2X1  _1217_
timestamp 0
transform 1 0 4210 0 1 5990
box -6 -8 66 268
use NAND2X1  _1218_
timestamp 0
transform -1 0 3950 0 1 5990
box -6 -8 66 268
use NAND2X1  _1219_
timestamp 0
transform -1 0 3250 0 -1 5990
box -6 -8 66 268
use NAND2X1  _1220_
timestamp 0
transform 1 0 3830 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1221_
timestamp 0
transform -1 0 3450 0 1 5470
box -6 -8 66 268
use NOR2X1  _1222_
timestamp 0
transform 1 0 3390 0 -1 3910
box -6 -8 66 268
use NOR2X1  _1223_
timestamp 0
transform -1 0 3550 0 -1 5990
box -6 -8 66 268
use NAND3X1  _1224_
timestamp 0
transform 1 0 3650 0 -1 5990
box -6 -8 86 268
use NOR2X1  _1225_
timestamp 0
transform -1 0 3790 0 1 5990
box -6 -8 66 268
use AOI21X1  _1226_
timestamp 0
transform -1 0 4070 0 -1 5990
box -6 -8 86 268
use NOR2X1  _1227_
timestamp 0
transform 1 0 3350 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1228_
timestamp 0
transform -1 0 3450 0 1 5990
box -6 -8 66 268
use OAI21X1  _1229_
timestamp 0
transform -1 0 3630 0 1 5990
box -6 -8 86 268
use AOI21X1  _1230_
timestamp 0
transform 1 0 2850 0 1 5470
box -6 -8 86 268
use NOR2X1  _1231_
timestamp 0
transform 1 0 2430 0 1 4950
box -6 -8 66 268
use NAND2X1  _1232_
timestamp 0
transform 1 0 2010 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1233_
timestamp 0
transform -1 0 1970 0 1 4430
box -6 -8 66 268
use AND2X2  _1234_
timestamp 0
transform -1 0 2330 0 1 4430
box -6 -8 86 268
use NAND3X1  _1235_
timestamp 0
transform 1 0 2530 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1236_
timestamp 0
transform -1 0 2790 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1237_
timestamp 0
transform 1 0 2890 0 -1 5470
box -6 -8 66 268
use INVX1  _1238_
timestamp 0
transform -1 0 1690 0 -1 1830
box -6 -8 46 268
use NOR2X1  _1239_
timestamp 0
transform -1 0 1910 0 1 1830
box -6 -8 66 268
use NOR2X1  _1240_
timestamp 0
transform 1 0 1930 0 1 2870
box -6 -8 66 268
use NOR2X1  _1241_
timestamp 0
transform -1 0 2490 0 1 4430
box -6 -8 66 268
use AOI21X1  _1242_
timestamp 0
transform -1 0 2110 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1243_
timestamp 0
transform 1 0 2210 0 -1 4430
box -6 -8 86 268
use INVX1  _1244_
timestamp 0
transform 1 0 1350 0 -1 4430
box -6 -8 46 268
use XOR2X1  _1245_
timestamp 0
transform -1 0 1810 0 1 4430
box -6 -8 126 268
use OAI21X1  _1246_
timestamp 0
transform 1 0 1670 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1247_
timestamp 0
transform -1 0 2850 0 1 4430
box -6 -8 86 268
use OAI21X1  _1248_
timestamp 0
transform 1 0 2590 0 1 4430
box -6 -8 86 268
use INVX1  _1249_
timestamp 0
transform -1 0 1590 0 1 4430
box -6 -8 46 268
use NAND3X1  _1250_
timestamp 0
transform -1 0 1570 0 -1 4430
box -6 -8 86 268
use AOI21X1  _1251_
timestamp 0
transform 1 0 1750 0 1 3910
box -6 -8 86 268
use AOI21X1  _1252_
timestamp 0
transform -1 0 2150 0 1 4430
box -6 -8 86 268
use NAND3X1  _1253_
timestamp 0
transform -1 0 2190 0 1 3910
box -6 -8 86 268
use OAI21X1  _1254_
timestamp 0
transform 1 0 1850 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1255_
timestamp 0
transform 1 0 1930 0 1 3910
box -6 -8 86 268
use NAND2X1  _1256_
timestamp 0
transform -1 0 1790 0 1 2350
box -6 -8 66 268
use NAND2X1  _1257_
timestamp 0
transform 1 0 2290 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1258_
timestamp 0
transform 1 0 2130 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1259_
timestamp 0
transform 1 0 1890 0 1 2350
box -6 -8 86 268
use NAND2X1  _1260_
timestamp 0
transform -1 0 1550 0 -1 1830
box -6 -8 66 268
use INVX1  _1261_
timestamp 0
transform -1 0 1450 0 1 2350
box -6 -8 46 268
use XOR2X1  _1262_
timestamp 0
transform 1 0 2030 0 -1 2870
box -6 -8 126 268
use XOR2X1  _1263_
timestamp 0
transform -1 0 2370 0 -1 2870
box -6 -8 126 268
use NAND3X1  _1264_
timestamp 0
transform -1 0 2170 0 1 3390
box -6 -8 86 268
use INVX1  _1265_
timestamp 0
transform -1 0 1970 0 -1 3910
box -6 -8 46 268
use AOI21X1  _1266_
timestamp 0
transform 1 0 1750 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1267_
timestamp 0
transform 1 0 2070 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1268_
timestamp 0
transform -1 0 2330 0 1 3390
box -6 -8 66 268
use NAND2X1  _1269_
timestamp 0
transform 1 0 2250 0 -1 3910
box -6 -8 66 268
use OAI22X1  _1270_
timestamp 0
transform -1 0 2510 0 -1 3910
box -6 -8 106 268
use INVX1  _1271_
timestamp 0
transform 1 0 2430 0 -1 2350
box -6 -8 46 268
use NAND2X1  _1272_
timestamp 0
transform 1 0 2070 0 1 2350
box -6 -8 66 268
use AOI22X1  _1273_
timestamp 0
transform -1 0 2750 0 -1 2870
box -6 -8 106 268
use NAND2X1  _1274_
timestamp 0
transform -1 0 370 0 1 790
box -6 -8 66 268
use OAI21X1  _1275_
timestamp 0
transform -1 0 550 0 1 790
box -6 -8 86 268
use OAI22X1  _1276_
timestamp 0
transform 1 0 110 0 1 790
box -6 -8 106 268
use NOR2X1  _1277_
timestamp 0
transform 1 0 450 0 -1 790
box -6 -8 66 268
use NOR2X1  _1278_
timestamp 0
transform -1 0 870 0 1 270
box -6 -8 66 268
use AOI21X1  _1279_
timestamp 0
transform 1 0 450 0 1 270
box -6 -8 86 268
use OR2X2  _1280_
timestamp 0
transform 1 0 270 0 1 270
box -6 -8 86 268
use NAND2X1  _1281_
timestamp 0
transform -1 0 1010 0 -1 270
box -6 -8 66 268
use AND2X2  _1282_
timestamp 0
transform -1 0 850 0 -1 270
box -6 -8 86 268
use NAND3X1  _1283_
timestamp 0
transform 1 0 630 0 1 270
box -6 -8 86 268
use NAND2X1  _1284_
timestamp 0
transform 1 0 1590 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1285_
timestamp 0
transform -1 0 1310 0 1 1310
box -6 -8 66 268
use NAND2X1  _1286_
timestamp 0
transform -1 0 1390 0 -1 1830
box -6 -8 66 268
use NOR2X1  _1287_
timestamp 0
transform -1 0 1410 0 1 1830
box -6 -8 66 268
use OAI21X1  _1288_
timestamp 0
transform 1 0 1950 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1289_
timestamp 0
transform -1 0 1230 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1290_
timestamp 0
transform -1 0 1250 0 1 1830
box -6 -8 86 268
use OAI21X1  _1291_
timestamp 0
transform 1 0 590 0 -1 270
box -6 -8 86 268
use NAND2X1  _1292_
timestamp 0
transform -1 0 170 0 1 270
box -6 -8 66 268
use NOR2X1  _1293_
timestamp 0
transform -1 0 170 0 -1 790
box -6 -8 66 268
use OAI21X1  _1294_
timestamp 0
transform -1 0 350 0 -1 790
box -6 -8 86 268
use AOI21X1  _1295_
timestamp 0
transform 1 0 610 0 -1 790
box -6 -8 86 268
use OAI21X1  _1296_
timestamp 0
transform -1 0 910 0 1 1830
box -6 -8 86 268
use NOR2X1  _1297_
timestamp 0
transform 1 0 1790 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1298_
timestamp 0
transform -1 0 1590 0 1 1830
box -6 -8 86 268
use NOR2X1  _1299_
timestamp 0
transform -1 0 1070 0 1 1830
box -6 -8 66 268
use NAND2X1  _1300_
timestamp 0
transform -1 0 1750 0 1 1830
box -6 -8 66 268
use NAND2X1  _1301_
timestamp 0
transform 1 0 2190 0 1 1830
box -6 -8 66 268
use NAND3X1  _1302_
timestamp 0
transform 1 0 2010 0 1 1830
box -6 -8 86 268
use NAND3X1  _1303_
timestamp 0
transform 1 0 2230 0 1 2350
box -6 -8 86 268
use NOR3X1  _1304_
timestamp 0
transform -1 0 2770 0 -1 3910
box -6 -8 166 268
use NAND3X1  _1305_
timestamp 0
transform -1 0 1650 0 -1 3910
box -6 -8 86 268
use AOI21X1  _1306_
timestamp 0
transform -1 0 1490 0 1 3910
box -6 -8 86 268
use NOR2X1  _1307_
timestamp 0
transform 1 0 1410 0 1 270
box -6 -8 66 268
use INVX8  _1308_
timestamp 0
transform 1 0 1390 0 1 2870
box -6 -8 106 268
use INVX1  _1309_
timestamp 0
transform -1 0 5310 0 -1 1310
box -6 -8 46 268
use NOR2X1  _1310_
timestamp 0
transform 1 0 2990 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1311_
timestamp 0
transform 1 0 2630 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1312_
timestamp 0
transform 1 0 1710 0 1 270
box -6 -8 66 268
use NAND3X1  _1313_
timestamp 0
transform 1 0 1750 0 -1 790
box -6 -8 86 268
use AOI21X1  _1314_
timestamp 0
transform 1 0 2810 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1315_
timestamp 0
transform -1 0 5090 0 -1 5990
box -6 -8 86 268
use NOR2X1  _1316_
timestamp 0
transform 1 0 5690 0 1 5470
box -6 -8 66 268
use AOI21X1  _1317_
timestamp 0
transform 1 0 5570 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1318_
timestamp 0
transform 1 0 5850 0 1 5470
box -6 -8 86 268
use NAND2X1  _1319_
timestamp 0
transform -1 0 5770 0 -1 5990
box -6 -8 66 268
use NAND3X1  _1320_
timestamp 0
transform -1 0 6490 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1321_
timestamp 0
transform -1 0 6770 0 1 5470
box -6 -8 66 268
use NAND2X1  _1322_
timestamp 0
transform -1 0 6830 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1323_
timestamp 0
transform 1 0 6790 0 1 5990
box -6 -8 66 268
use OAI21X1  _1324_
timestamp 0
transform 1 0 5050 0 1 5990
box -6 -8 86 268
use OAI21X1  _1325_
timestamp 0
transform -1 0 5590 0 1 5470
box -6 -8 86 268
use NAND3X1  _1326_
timestamp 0
transform 1 0 5370 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1327_
timestamp 0
transform 1 0 5570 0 1 5990
box -6 -8 86 268
use NAND3X1  _1328_
timestamp 0
transform 1 0 5750 0 1 5990
box -6 -8 86 268
use AOI21X1  _1329_
timestamp 0
transform 1 0 5930 0 1 5990
box -6 -8 86 268
use NAND3X1  _1330_
timestamp 0
transform 1 0 5470 0 -1 4950
box -6 -8 86 268
use INVX1  _1331_
timestamp 0
transform 1 0 6470 0 -1 4950
box -6 -8 46 268
use NAND2X1  _1332_
timestamp 0
transform -1 0 5870 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1333_
timestamp 0
transform 1 0 5970 0 -1 4950
box -6 -8 66 268
use AOI21X1  _1334_
timestamp 0
transform -1 0 6270 0 1 4950
box -6 -8 86 268
use NOR2X1  _1335_
timestamp 0
transform 1 0 6430 0 -1 4430
box -6 -8 66 268
use NOR2X1  _1336_
timestamp 0
transform 1 0 6590 0 -1 4430
box -6 -8 66 268
use NAND2X1  _1337_
timestamp 0
transform -1 0 6810 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1338_
timestamp 0
transform -1 0 6830 0 -1 5470
box -6 -8 86 268
use INVX1  _1339_
timestamp 0
transform -1 0 6890 0 1 3910
box -6 -8 46 268
use NOR2X1  _1340_
timestamp 0
transform 1 0 6530 0 1 3910
box -6 -8 66 268
use OAI21X1  _1341_
timestamp 0
transform -1 0 6950 0 1 5470
box -6 -8 86 268
use NOR2X1  _1342_
timestamp 0
transform 1 0 5650 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1343_
timestamp 0
transform 1 0 6610 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1344_
timestamp 0
transform -1 0 6830 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1345_
timestamp 0
transform 1 0 6670 0 1 4950
box -6 -8 86 268
use NAND3X1  _1346_
timestamp 0
transform 1 0 6610 0 1 5990
box -6 -8 86 268
use AND2X2  _1347_
timestamp 0
transform 1 0 5870 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1348_
timestamp 0
transform 1 0 6370 0 1 5470
box -6 -8 86 268
use NAND2X1  _1349_
timestamp 0
transform -1 0 6650 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1350_
timestamp 0
transform 1 0 6550 0 1 5470
box -6 -8 66 268
use AOI21X1  _1351_
timestamp 0
transform 1 0 5550 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1352_
timestamp 0
transform 1 0 5770 0 -1 6510
box -6 -8 66 268
use OAI21X1  _1353_
timestamp 0
transform -1 0 6010 0 -1 6510
box -6 -8 86 268
use NAND3X1  _1354_
timestamp 0
transform 1 0 6110 0 1 5990
box -6 -8 86 268
use NAND3X1  _1355_
timestamp 0
transform 1 0 6410 0 -1 5990
box -6 -8 86 268
use AND2X2  _1356_
timestamp 0
transform 1 0 6590 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1357_
timestamp 0
transform -1 0 6310 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1358_
timestamp 0
transform 1 0 6050 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1359_
timestamp 0
transform 1 0 6510 0 1 4950
box -6 -8 66 268
use NOR2X1  _1360_
timestamp 0
transform 1 0 6130 0 -1 4950
box -6 -8 66 268
use NAND3X1  _1361_
timestamp 0
transform -1 0 6370 0 -1 4950
box -6 -8 86 268
use NOR2X1  _1362_
timestamp 0
transform -1 0 6790 0 -1 3910
box -6 -8 66 268
use NOR2X1  _1363_
timestamp 0
transform 1 0 6690 0 1 3910
box -6 -8 66 268
use NAND3X1  _1364_
timestamp 0
transform -1 0 6830 0 1 4430
box -6 -8 86 268
use OR2X2  _1365_
timestamp 0
transform -1 0 6930 0 1 4950
box -6 -8 86 268
use NAND2X1  _1366_
timestamp 0
transform -1 0 6150 0 -1 5470
box -6 -8 66 268
use OAI21X1  _1367_
timestamp 0
transform -1 0 6310 0 -1 5470
box -6 -8 86 268
use INVX1  _1368_
timestamp 0
transform -1 0 5410 0 1 2870
box -6 -8 46 268
use NAND2X1  _1369_
timestamp 0
transform -1 0 4630 0 1 2870
box -6 -8 66 268
use NOR2X1  _1370_
timestamp 0
transform 1 0 3910 0 1 2870
box -6 -8 66 268
use INVX1  _1371_
timestamp 0
transform 1 0 4250 0 1 2870
box -6 -8 46 268
use OR2X2  _1372_
timestamp 0
transform -1 0 5210 0 1 3390
box -6 -8 86 268
use OAI22X1  _1373_
timestamp 0
transform -1 0 4810 0 1 3390
box -6 -8 106 268
use NAND3X1  _1374_
timestamp 0
transform 1 0 5850 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1375_
timestamp 0
transform -1 0 5450 0 1 3910
box -6 -8 66 268
use NAND2X1  _1376_
timestamp 0
transform 1 0 6570 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1377_
timestamp 0
transform -1 0 6930 0 1 3390
box -6 -8 66 268
use OAI21X1  _1378_
timestamp 0
transform -1 0 6710 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1379_
timestamp 0
transform -1 0 6770 0 1 3390
box -6 -8 86 268
use NAND3X1  _1380_
timestamp 0
transform 1 0 6210 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1381_
timestamp 0
transform -1 0 6470 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1382_
timestamp 0
transform -1 0 5750 0 -1 3910
box -6 -8 86 268
use AOI22X1  _1383_
timestamp 0
transform 1 0 4830 0 1 3910
box -6 -8 106 268
use NAND2X1  _1384_
timestamp 0
transform -1 0 5050 0 -1 3910
box -6 -8 66 268
use AOI22X1  _1385_
timestamp 0
transform -1 0 5330 0 -1 4430
box -6 -8 106 268
use OAI22X1  _1386_
timestamp 0
transform -1 0 5130 0 -1 4430
box -6 -8 106 268
use AOI21X1  _1387_
timestamp 0
transform -1 0 5110 0 1 3910
box -6 -8 86 268
use AOI22X1  _1388_
timestamp 0
transform 1 0 4330 0 1 3390
box -6 -8 106 268
use OAI21X1  _1389_
timestamp 0
transform -1 0 4610 0 1 3390
box -6 -8 86 268
use OAI21X1  _1390_
timestamp 0
transform -1 0 2010 0 1 1310
box -6 -8 86 268
use NOR2X1  _1391_
timestamp 0
transform -1 0 1450 0 1 790
box -6 -8 66 268
use AND2X2  _1392_
timestamp 0
transform -1 0 1490 0 1 1310
box -6 -8 86 268
use NAND3X1  _1393_
timestamp 0
transform -1 0 990 0 1 1310
box -6 -8 86 268
use NOR2X1  _1394_
timestamp 0
transform 1 0 990 0 -1 1830
box -6 -8 66 268
use AOI21X1  _1395_
timestamp 0
transform -1 0 4230 0 -1 5470
box -6 -8 86 268
use INVX1  _1396_
timestamp 0
transform -1 0 3070 0 -1 2870
box -6 -8 46 268
use NAND3X1  _1397_
timestamp 0
transform 1 0 2850 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1398_
timestamp 0
transform 1 0 4390 0 1 2870
box -6 -8 86 268
use AOI22X1  _1399_
timestamp 0
transform 1 0 4530 0 1 1310
box -6 -8 106 268
use OAI21X1  _1400_
timestamp 0
transform 1 0 6030 0 1 5470
box -6 -8 86 268
use NOR2X1  _1401_
timestamp 0
transform -1 0 5990 0 -1 5470
box -6 -8 66 268
use NAND2X1  _1402_
timestamp 0
transform -1 0 4530 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1403_
timestamp 0
transform 1 0 4790 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1404_
timestamp 0
transform 1 0 4630 0 -1 4950
box -6 -8 66 268
use NOR2X1  _1405_
timestamp 0
transform 1 0 4930 0 1 4950
box -6 -8 66 268
use NAND3X1  _1406_
timestamp 0
transform -1 0 5030 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1407_
timestamp 0
transform -1 0 5210 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1408_
timestamp 0
transform 1 0 5090 0 -1 1310
box -6 -8 86 268
use INVX1  _1409_
timestamp 0
transform -1 0 5130 0 1 270
box -6 -8 46 268
use NAND2X1  _1410_
timestamp 0
transform 1 0 4370 0 1 1310
box -6 -8 66 268
use NAND2X1  _1411_
timestamp 0
transform -1 0 6170 0 -1 6510
box -6 -8 66 268
use AND2X2  _1412_
timestamp 0
transform 1 0 5390 0 1 5990
box -6 -8 86 268
use NAND3X1  _1413_
timestamp 0
transform 1 0 6270 0 -1 6510
box -6 -8 86 268
use NOR3X1  _1414_
timestamp 0
transform -1 0 6750 0 -1 6510
box -6 -8 166 268
use NAND2X1  _1415_
timestamp 0
transform -1 0 6330 0 1 5990
box -6 -8 66 268
use AOI21X1  _1416_
timestamp 0
transform -1 0 6510 0 1 5990
box -6 -8 86 268
use OAI21X1  _1417_
timestamp 0
transform -1 0 5590 0 1 2870
box -6 -8 86 268
use AOI21X1  _1418_
timestamp 0
transform -1 0 5130 0 1 1310
box -6 -8 86 268
use AOI22X1  _1419_
timestamp 0
transform -1 0 4530 0 -1 3910
box -6 -8 106 268
use AND2X2  _1420_
timestamp 0
transform -1 0 4890 0 -1 3910
box -6 -8 86 268
use OAI22X1  _1421_
timestamp 0
transform -1 0 4730 0 1 3910
box -6 -8 106 268
use AOI22X1  _1422_
timestamp 0
transform 1 0 4430 0 1 3910
box -6 -8 106 268
use OAI21X1  _1423_
timestamp 0
transform -1 0 4710 0 -1 3910
box -6 -8 86 268
use OAI22X1  _1424_
timestamp 0
transform 1 0 4050 0 -1 3910
box -6 -8 106 268
use AOI21X1  _1425_
timestamp 0
transform -1 0 4330 0 -1 3910
box -6 -8 86 268
use AND2X2  _1426_
timestamp 0
transform 1 0 810 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1427_
timestamp 0
transform 1 0 630 0 -1 1830
box -6 -8 86 268
use NOR3X1  _1428_
timestamp 0
transform 1 0 2410 0 1 2350
box -6 -8 166 268
use OAI21X1  _1429_
timestamp 0
transform -1 0 4150 0 1 2870
box -6 -8 86 268
use AOI21X1  _1430_
timestamp 0
transform -1 0 4810 0 1 2870
box -6 -8 86 268
use INVX1  _1431_
timestamp 0
transform -1 0 4950 0 1 1310
box -6 -8 46 268
use NAND3X1  _1432_
timestamp 0
transform -1 0 4810 0 1 1310
box -6 -8 86 268
use OAI21X1  _1433_
timestamp 0
transform -1 0 4990 0 1 270
box -6 -8 86 268
use INVX2  _1434_
timestamp 0
transform 1 0 2430 0 1 270
box -6 -8 46 268
use OAI21X1  _1435_
timestamp 0
transform 1 0 4730 0 1 270
box -6 -8 86 268
use NOR2X1  _1436_
timestamp 0
transform -1 0 2350 0 1 3910
box -6 -8 66 268
use NOR2X1  _1437_
timestamp 0
transform 1 0 2390 0 -1 4430
box -6 -8 66 268
use AND2X2  _1438_
timestamp 0
transform 1 0 2450 0 1 3910
box -6 -8 86 268
use NAND2X1  _1439_
timestamp 0
transform 1 0 2710 0 -1 4430
box -6 -8 66 268
use NAND2X1  _1440_
timestamp 0
transform 1 0 3030 0 -1 4430
box -6 -8 66 268
use NOR2X1  _1441_
timestamp 0
transform -1 0 2930 0 -1 4430
box -6 -8 66 268
use NAND3X1  _1442_
timestamp 0
transform 1 0 2790 0 1 3910
box -6 -8 86 268
use INVX1  _1443_
timestamp 0
transform 1 0 2250 0 1 2870
box -6 -8 46 268
use NOR2X1  _1444_
timestamp 0
transform 1 0 1730 0 1 3390
box -6 -8 66 268
use NOR2X1  _1445_
timestamp 0
transform 1 0 1770 0 -1 3390
box -6 -8 66 268
use AND2X2  _1446_
timestamp 0
transform 1 0 2430 0 1 3390
box -6 -8 86 268
use NAND3X1  _1447_
timestamp 0
transform 1 0 2550 0 1 2870
box -6 -8 86 268
use NOR2X1  _1448_
timestamp 0
transform 1 0 2930 0 1 1830
box -6 -8 66 268
use INVX2  _1449_
timestamp 0
transform 1 0 4410 0 -1 1310
box -6 -8 46 268
use OAI21X1  _1450_
timestamp 0
transform -1 0 4310 0 -1 1830
box -6 -8 86 268
use XOR2X1  _1451_
timestamp 0
transform 1 0 4870 0 -1 1310
box -6 -8 126 268
use NOR2X1  _1452_
timestamp 0
transform 1 0 2870 0 -1 790
box -6 -8 66 268
use NOR2X1  _1453_
timestamp 0
transform 1 0 2690 0 1 790
box -6 -8 66 268
use INVX1  _1454_
timestamp 0
transform -1 0 2890 0 1 790
box -6 -8 46 268
use NAND2X1  _1455_
timestamp 0
transform -1 0 5350 0 -1 790
box -6 -8 66 268
use NAND2X1  _1456_
timestamp 0
transform 1 0 5310 0 1 790
box -6 -8 66 268
use NOR2X1  _1457_
timestamp 0
transform -1 0 5510 0 -1 790
box -6 -8 66 268
use OAI21X1  _1458_
timestamp 0
transform -1 0 5550 0 1 790
box -6 -8 86 268
use XOR2X1  _1459_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 126 268
use NAND2X1  _1460_
timestamp 0
transform 1 0 4470 0 1 790
box -6 -8 66 268
use OAI21X1  _1461_
timestamp 0
transform 1 0 3530 0 1 790
box -6 -8 86 268
use AOI21X1  _1462_
timestamp 0
transform -1 0 3210 0 1 790
box -6 -8 86 268
use XOR2X1  _1463_
timestamp 0
transform 1 0 2830 0 -1 270
box -6 -8 126 268
use NAND2X1  _1464_
timestamp 0
transform 1 0 2270 0 1 270
box -6 -8 66 268
use NAND2X1  _1465_
timestamp 0
transform 1 0 2570 0 1 270
box -6 -8 66 268
use NAND2X1  _1466_
timestamp 0
transform -1 0 2790 0 1 270
box -6 -8 66 268
use INVX1  _1467_
timestamp 0
transform 1 0 3050 0 -1 270
box -6 -8 46 268
use NAND2X1  _1468_
timestamp 0
transform 1 0 3190 0 -1 270
box -6 -8 66 268
use OAI21X1  _1469_
timestamp 0
transform 1 0 2650 0 -1 270
box -6 -8 86 268
use OAI21X1  _1470_
timestamp 0
transform 1 0 3650 0 -1 270
box -6 -8 86 268
use XOR2X1  _1471_
timestamp 0
transform -1 0 3990 0 1 270
box -6 -8 126 268
use NAND2X1  _1472_
timestamp 0
transform -1 0 3890 0 -1 270
box -6 -8 66 268
use OAI21X1  _1473_
timestamp 0
transform 1 0 4090 0 1 270
box -6 -8 86 268
use XNOR2X1  _1474_
timestamp 0
transform 1 0 5190 0 -1 270
box -6 -8 126 268
use NAND2X1  _1475_
timestamp 0
transform -1 0 4330 0 1 270
box -6 -8 66 268
use NAND2X1  _1476_
timestamp 0
transform -1 0 4910 0 -1 270
box -6 -8 66 268
use INVX1  _1477_
timestamp 0
transform 1 0 4590 0 1 270
box -6 -8 46 268
use NAND3X1  _1478_
timestamp 0
transform -1 0 4750 0 -1 270
box -6 -8 86 268
use NAND2X1  _1479_
timestamp 0
transform -1 0 4490 0 1 270
box -6 -8 66 268
use INVX1  _1480_
timestamp 0
transform 1 0 6030 0 1 790
box -6 -8 46 268
use NAND2X1  _1481_
timestamp 0
transform 1 0 5870 0 1 790
box -6 -8 66 268
use XOR2X1  _1482_
timestamp 0
transform -1 0 5770 0 1 790
box -6 -8 126 268
use XNOR2X1  _1483_
timestamp 0
transform 1 0 3650 0 1 270
box -6 -8 126 268
use OAI21X1  _1484_
timestamp 0
transform -1 0 2970 0 1 270
box -6 -8 86 268
use XNOR2X1  _1485_
timestamp 0
transform 1 0 3070 0 1 270
box -6 -8 126 268
use INVX1  _1486_
timestamp 0
transform 1 0 3510 0 -1 270
box -6 -8 46 268
use NAND2X1  _1487_
timestamp 0
transform 1 0 3350 0 -1 270
box -6 -8 66 268
use NAND2X1  _1488_
timestamp 0
transform 1 0 3030 0 -1 790
box -6 -8 66 268
use NOR2X1  _1489_
timestamp 0
transform 1 0 2990 0 1 790
box -6 -8 66 268
use XNOR2X1  _1490_
timestamp 0
transform -1 0 3430 0 1 790
box -6 -8 126 268
use INVX1  _1491_
timestamp 0
transform -1 0 4770 0 -1 1310
box -6 -8 46 268
use XNOR2X1  _1492_
timestamp 0
transform -1 0 4750 0 1 790
box -6 -8 126 268
use NAND3X1  _1493_
timestamp 0
transform -1 0 4150 0 1 790
box -6 -8 86 268
use AOI21X1  _1494_
timestamp 0
transform 1 0 3570 0 -1 790
box -6 -8 86 268
use NAND3X1  _1495_
timestamp 0
transform 1 0 3750 0 -1 790
box -6 -8 86 268
use OAI21X1  _1496_
timestamp 0
transform -1 0 4550 0 -1 790
box -6 -8 86 268
use OAI21X1  _1497_
timestamp 0
transform 1 0 5010 0 -1 270
box -6 -8 86 268
use NAND2X1  _1498_
timestamp 0
transform 1 0 4510 0 -1 270
box -6 -8 66 268
use OAI21X1  _1499_
timestamp 0
transform 1 0 4330 0 -1 270
box -6 -8 86 268
use NOR2X1  _1500_
timestamp 0
transform -1 0 4050 0 -1 270
box -6 -8 66 268
use AOI21X1  _1501_
timestamp 0
transform 1 0 4150 0 -1 270
box -6 -8 86 268
use XOR2X1  _1502_
timestamp 0
transform 1 0 4250 0 1 790
box -6 -8 126 268
use XOR2X1  _1503_
timestamp 0
transform 1 0 4250 0 -1 790
box -6 -8 126 268
use NAND3X1  _1504_
timestamp 0
transform -1 0 4630 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1505_
timestamp 0
transform -1 0 4270 0 1 1310
box -6 -8 86 268
use OAI21X1  _1506_
timestamp 0
transform 1 0 4410 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1507_
timestamp 0
transform 1 0 4650 0 -1 790
box -6 -8 86 268
use OAI21X1  _1508_
timestamp 0
transform 1 0 4850 0 1 790
box -6 -8 86 268
use NAND3X1  _1509_
timestamp 0
transform 1 0 2250 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1510_
timestamp 0
transform -1 0 2690 0 1 3910
box -6 -8 86 268
use OR2X2  _1511_
timestamp 0
transform 1 0 2430 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1512_
timestamp 0
transform 1 0 2550 0 -1 4430
box -6 -8 66 268
use NAND3X1  _1513_
timestamp 0
transform -1 0 2690 0 1 3390
box -6 -8 86 268
use NOR2X1  _1514_
timestamp 0
transform -1 0 2670 0 -1 3390
box -6 -8 66 268
use NAND2X1  _1515_
timestamp 0
transform 1 0 2730 0 1 2870
box -6 -8 66 268
use NOR2X1  _1516_
timestamp 0
transform -1 0 2950 0 1 2870
box -6 -8 66 268
use INVX1  _1517_
timestamp 0
transform 1 0 3790 0 -1 1830
box -6 -8 46 268
use NOR2X1  _1518_
timestamp 0
transform 1 0 4070 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1519_
timestamp 0
transform -1 0 4310 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1520_
timestamp 0
transform 1 0 3230 0 1 1310
box -6 -8 86 268
use NOR2X1  _1521_
timestamp 0
transform -1 0 4090 0 1 1310
box -6 -8 66 268
use NAND3X1  _1522_
timestamp 0
transform -1 0 3970 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1523_
timestamp 0
transform 1 0 3050 0 1 1310
box -6 -8 86 268
use NAND2X1  _1524_
timestamp 0
transform -1 0 4150 0 -1 790
box -6 -8 66 268
use NOR2X1  _1525_
timestamp 0
transform 1 0 3230 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1526_
timestamp 0
transform 1 0 3390 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1527_
timestamp 0
transform 1 0 3030 0 1 5470
box -6 -8 66 268
use NAND3X1  _1528_
timestamp 0
transform -1 0 3130 0 -1 5470
box -6 -8 86 268
use NOR2X1  _1529_
timestamp 0
transform -1 0 1350 0 -1 2350
box -6 -8 66 268
use NAND3X1  _1530_
timestamp 0
transform 1 0 1450 0 -1 2350
box -6 -8 86 268
use NOR2X1  _1531_
timestamp 0
transform 1 0 1590 0 1 3910
box -6 -8 66 268
use NAND3X1  _1532_
timestamp 0
transform -1 0 2010 0 -1 3390
box -6 -8 86 268
use NOR2X1  _1533_
timestamp 0
transform -1 0 2150 0 1 2870
box -6 -8 66 268
use NAND2X1  _1534_
timestamp 0
transform -1 0 2450 0 1 2870
box -6 -8 66 268
use NOR2X1  _1535_
timestamp 0
transform -1 0 2830 0 -1 3390
box -6 -8 66 268
use NAND3X1  _1536_
timestamp 0
transform -1 0 3470 0 -1 790
box -6 -8 86 268
use OAI22X1  _1537_
timestamp 0
transform 1 0 2530 0 -1 790
box -6 -8 106 268
use INVX1  _1538_
timestamp 0
transform 1 0 3930 0 1 790
box -6 -8 46 268
use OR2X2  _1539_
timestamp 0
transform -1 0 3370 0 1 270
box -6 -8 86 268
use OAI22X1  _1540_
timestamp 0
transform 1 0 1870 0 1 270
box -6 -8 106 268
use OR2X2  _1541_
timestamp 0
transform -1 0 3550 0 1 270
box -6 -8 86 268
use OAI22X1  _1542_
timestamp 0
transform 1 0 2070 0 1 270
box -6 -8 106 268
use NAND2X1  _1543_
timestamp 0
transform 1 0 3930 0 -1 790
box -6 -8 66 268
use OAI22X1  _1544_
timestamp 0
transform 1 0 3190 0 -1 790
box -6 -8 106 268
use NOR2X1  _1545_
timestamp 0
transform 1 0 2490 0 1 1830
box -6 -8 66 268
use NAND2X1  _1546_
timestamp 0
transform 1 0 3630 0 -1 1830
box -6 -8 66 268
use XOR2X1  _1547_
timestamp 0
transform 1 0 4790 0 -1 2870
box -6 -8 126 268
use INVX1  _1548_
timestamp 0
transform 1 0 3930 0 -1 1830
box -6 -8 46 268
use NOR2X1  _1549_
timestamp 0
transform -1 0 4970 0 1 1830
box -6 -8 66 268
use XOR2X1  _1550_
timestamp 0
transform 1 0 5050 0 -1 1830
box -6 -8 126 268
use XNOR2X1  _1551_
timestamp 0
transform -1 0 5350 0 1 1830
box -6 -8 126 268
use OAI21X1  _1552_
timestamp 0
transform 1 0 4490 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1553_
timestamp 0
transform -1 0 4630 0 1 1830
box -6 -8 86 268
use INVX1  _1554_
timestamp 0
transform 1 0 5270 0 -1 1830
box -6 -8 46 268
use NAND2X1  _1555_
timestamp 0
transform 1 0 5070 0 1 1830
box -6 -8 66 268
use OAI21X1  _1556_
timestamp 0
transform -1 0 5150 0 -1 2350
box -6 -8 86 268
use NOR2X1  _1557_
timestamp 0
transform -1 0 4930 0 1 2350
box -6 -8 66 268
use INVX2  _1558_
timestamp 0
transform -1 0 3870 0 -1 2870
box -6 -8 46 268
use NOR2X1  _1559_
timestamp 0
transform 1 0 5010 0 -1 2870
box -6 -8 66 268
use NOR2X1  _1560_
timestamp 0
transform -1 0 5090 0 1 2350
box -6 -8 66 268
use XNOR2X1  _1561_
timestamp 0
transform -1 0 4790 0 -1 2350
box -6 -8 126 268
use OAI21X1  _1562_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 86 268
use OAI21X1  _1563_
timestamp 0
transform -1 0 4270 0 1 1830
box -6 -8 86 268
use AOI21X1  _1564_
timestamp 0
transform -1 0 4970 0 -1 2350
box -6 -8 86 268
use INVX1  _1565_
timestamp 0
transform 1 0 3590 0 -1 2350
box -6 -8 46 268
use NOR2X1  _1566_
timestamp 0
transform 1 0 3530 0 -1 2870
box -6 -8 66 268
use INVX1  _1567_
timestamp 0
transform -1 0 3070 0 1 2350
box -6 -8 46 268
use NOR2X1  _1568_
timestamp 0
transform 1 0 3690 0 -1 2870
box -6 -8 66 268
use INVX1  _1569_
timestamp 0
transform -1 0 3370 0 1 2350
box -6 -8 46 268
use NAND2X1  _1570_
timestamp 0
transform 1 0 3170 0 1 2350
box -6 -8 66 268
use OAI21X1  _1571_
timestamp 0
transform 1 0 3230 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1572_
timestamp 0
transform 1 0 3410 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1573_
timestamp 0
transform 1 0 3970 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1574_
timestamp 0
transform -1 0 4550 0 1 2350
box -6 -8 66 268
use NOR2X1  _1575_
timestamp 0
transform -1 0 4050 0 1 2350
box -6 -8 66 268
use NOR2X1  _1576_
timestamp 0
transform -1 0 4210 0 1 2350
box -6 -8 66 268
use OAI21X1  _1577_
timestamp 0
transform -1 0 3550 0 1 2350
box -6 -8 86 268
use NAND2X1  _1578_
timestamp 0
transform -1 0 3890 0 1 2350
box -6 -8 66 268
use OR2X2  _1579_
timestamp 0
transform 1 0 3650 0 1 2350
box -6 -8 86 268
use NAND3X1  _1580_
timestamp 0
transform 1 0 3730 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1581_
timestamp 0
transform -1 0 3990 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1582_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 86 268
use OAI21X1  _1583_
timestamp 0
transform -1 0 4170 0 -1 2350
box -6 -8 86 268
use XOR2X1  _1584_
timestamp 0
transform -1 0 4770 0 1 2350
box -6 -8 126 268
use XNOR2X1  _1585_
timestamp 0
transform 1 0 4270 0 -1 2350
box -6 -8 126 268
use OAI21X1  _1586_
timestamp 0
transform -1 0 4810 0 1 1830
box -6 -8 86 268
use XOR2X1  _1587_
timestamp 0
transform -1 0 3430 0 -1 2870
box -6 -8 126 268
use INVX1  _1588_
timestamp 0
transform -1 0 3210 0 -1 2870
box -6 -8 46 268
use OAI21X1  _1589_
timestamp 0
transform -1 0 4550 0 -1 2870
box -6 -8 86 268
use INVX1  _1590_
timestamp 0
transform -1 0 4370 0 -1 2870
box -6 -8 46 268
use AND2X2  _1591_
timestamp 0
transform 1 0 4310 0 1 2350
box -6 -8 86 268
use AOI21X1  _1592_
timestamp 0
transform 1 0 4150 0 -1 2870
box -6 -8 86 268
use AND2X2  _1593_
timestamp 0
transform 1 0 2670 0 1 2350
box -6 -8 86 268
use OAI21X1  _1594_
timestamp 0
transform 1 0 2850 0 1 2350
box -6 -8 86 268
use OAI22X1  _1595_
timestamp 0
transform -1 0 3130 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1596_
timestamp 0
transform -1 0 3290 0 1 2870
box -6 -8 66 268
use OAI21X1  _1597_
timestamp 0
transform 1 0 3050 0 1 2870
box -6 -8 86 268
use NAND2X1  _1598_
timestamp 0
transform -1 0 3450 0 1 2870
box -6 -8 66 268
use OAI21X1  _1599_
timestamp 0
transform -1 0 3810 0 1 2870
box -6 -8 86 268
use NAND3X1  _1600_
timestamp 0
transform 1 0 3550 0 1 2870
box -6 -8 86 268
use XOR2X1  _1601_
timestamp 0
transform -1 0 3590 0 -1 3390
box -6 -8 126 268
use OAI21X1  _1602_
timestamp 0
transform -1 0 3010 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1603_
timestamp 0
transform -1 0 3190 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1604_
timestamp 0
transform -1 0 3370 0 -1 3390
box -6 -8 86 268
use XOR2X1  _1605_
timestamp 0
transform 1 0 4150 0 -1 3390
box -6 -8 126 268
use NOR2X1  _1606_
timestamp 0
transform 1 0 6350 0 1 4950
box -6 -8 66 268
use NAND3X1  _1607_
timestamp 0
transform 1 0 6310 0 -1 2350
box -6 -8 86 268
use NOR2X1  _1608_
timestamp 0
transform -1 0 6530 0 -1 3390
box -6 -8 66 268
use NAND3X1  _1609_
timestamp 0
transform 1 0 6250 0 1 2350
box -6 -8 86 268
use OAI21X1  _1610_
timestamp 0
transform 1 0 6650 0 -1 2350
box -6 -8 86 268
use INVX1  _1611_
timestamp 0
transform 1 0 5690 0 1 1310
box -6 -8 46 268
use INVX1  _1612_
timestamp 0
transform -1 0 6930 0 -1 3910
box -6 -8 46 268
use NAND3X1  _1613_
timestamp 0
transform -1 0 6590 0 1 3390
box -6 -8 86 268
use OAI21X1  _1614_
timestamp 0
transform -1 0 6410 0 1 3390
box -6 -8 86 268
use NAND3X1  _1615_
timestamp 0
transform -1 0 6230 0 1 3390
box -6 -8 86 268
use NAND3X1  _1616_
timestamp 0
transform 1 0 5970 0 1 3390
box -6 -8 86 268
use NOR2X1  _1617_
timestamp 0
transform 1 0 5710 0 -1 3390
box -6 -8 66 268
use AOI21X1  _1618_
timestamp 0
transform -1 0 5570 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1619_
timestamp 0
transform 1 0 5410 0 -1 1830
box -6 -8 66 268
use XOR2X1  _1620_
timestamp 0
transform -1 0 6290 0 1 790
box -6 -8 126 268
use NOR2X1  _1621_
timestamp 0
transform 1 0 5410 0 -1 1310
box -6 -8 66 268
use INVX1  _1622_
timestamp 0
transform 1 0 6830 0 -1 2350
box -6 -8 46 268
use NOR2X1  _1623_
timestamp 0
transform 1 0 6490 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1624_
timestamp 0
transform -1 0 6950 0 -1 1830
box -6 -8 86 268
use INVX1  _1625_
timestamp 0
transform -1 0 6650 0 -1 1310
box -6 -8 46 268
use NOR2X1  _1626_
timestamp 0
transform 1 0 6610 0 1 1310
box -6 -8 66 268
use NOR2X1  _1627_
timestamp 0
transform 1 0 6450 0 -1 1310
box -6 -8 66 268
use XOR2X1  _1628_
timestamp 0
transform -1 0 6350 0 -1 1310
box -6 -8 126 268
use MUX2X1  _1629_
timestamp 0
transform 1 0 6030 0 -1 1310
box -6 -8 106 268
use AOI21X1  _1630_
timestamp 0
transform 1 0 6750 0 -1 1310
box -6 -8 86 268
use INVX1  _1631_
timestamp 0
transform -1 0 6830 0 -1 790
box -6 -8 46 268
use XOR2X1  _1632_
timestamp 0
transform -1 0 6790 0 -1 270
box -6 -8 126 268
use NAND2X1  _1633_
timestamp 0
transform -1 0 6750 0 1 270
box -6 -8 66 268
use OR2X2  _1634_
timestamp 0
transform -1 0 6590 0 1 270
box -6 -8 86 268
use NAND3X1  _1635_
timestamp 0
transform 1 0 6330 0 1 270
box -6 -8 86 268
use OAI21X1  _1636_
timestamp 0
transform -1 0 6570 0 -1 270
box -6 -8 86 268
use OAI21X1  _1637_
timestamp 0
transform 1 0 6150 0 1 270
box -6 -8 86 268
use XOR2X1  _1638_
timestamp 0
transform -1 0 6650 0 1 790
box -6 -8 126 268
use XNOR2X1  _1639_
timestamp 0
transform 1 0 6410 0 -1 790
box -6 -8 126 268
use MUX2X1  _1640_
timestamp 0
transform 1 0 5750 0 -1 790
box -6 -8 106 268
use OAI21X1  _1641_
timestamp 0
transform -1 0 6870 0 1 2350
box -6 -8 86 268
use NAND2X1  _1642_
timestamp 0
transform -1 0 6350 0 -1 2870
box -6 -8 66 268
use NAND2X1  _1643_
timestamp 0
transform -1 0 6650 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1644_
timestamp 0
transform -1 0 6370 0 1 1310
box -6 -8 86 268
use NAND2X1  _1645_
timestamp 0
transform 1 0 6630 0 -1 790
box -6 -8 66 268
use OAI21X1  _1646_
timestamp 0
transform -1 0 6830 0 1 790
box -6 -8 86 268
use XOR2X1  _1647_
timestamp 0
transform -1 0 6190 0 -1 2870
box -6 -8 126 268
use MUX2X1  _1648_
timestamp 0
transform 1 0 5870 0 -1 2870
box -6 -8 106 268
use NAND3X1  _1649_
timestamp 0
transform -1 0 6830 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1650_
timestamp 0
transform -1 0 6830 0 1 2870
box -6 -8 86 268
use XOR2X1  _1651_
timestamp 0
transform -1 0 6430 0 1 2870
box -6 -8 126 268
use XOR2X1  _1652_
timestamp 0
transform -1 0 6650 0 1 2870
box -6 -8 126 268
use MUX2X1  _1653_
timestamp 0
transform 1 0 5670 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1654_
timestamp 0
transform 1 0 6430 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1655_
timestamp 0
transform 1 0 6430 0 1 2350
box -6 -8 86 268
use AOI21X1  _1656_
timestamp 0
transform 1 0 6610 0 1 2350
box -6 -8 86 268
use OAI21X1  _1657_
timestamp 0
transform -1 0 6930 0 1 270
box -6 -8 86 268
use NAND2X1  _1658_
timestamp 0
transform 1 0 6210 0 -1 1830
box -6 -8 66 268
use NAND2X1  _1659_
timestamp 0
transform -1 0 6950 0 -1 270
box -6 -8 66 268
use OR2X2  _1660_
timestamp 0
transform -1 0 6750 0 1 1830
box -6 -8 86 268
use NAND2X1  _1661_
timestamp 0
transform -1 0 6910 0 1 1830
box -6 -8 66 268
use NAND3X1  _1662_
timestamp 0
transform -1 0 6570 0 1 1830
box -6 -8 86 268
use OAI21X1  _1663_
timestamp 0
transform 1 0 6090 0 1 1830
box -6 -8 86 268
use XOR2X1  _1664_
timestamp 0
transform 1 0 6270 0 1 1830
box -6 -8 126 268
use NAND3X1  _1665_
timestamp 0
transform -1 0 6450 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1666_
timestamp 0
transform -1 0 6770 0 -1 1830
box -6 -8 86 268
use INVX1  _1667_
timestamp 0
transform 1 0 6470 0 1 1310
box -6 -8 46 268
use NAND2X1  _1668_
timestamp 0
transform 1 0 6770 0 1 1310
box -6 -8 66 268
use NAND3X1  _1669_
timestamp 0
transform -1 0 6110 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1670_
timestamp 0
transform 1 0 5910 0 1 1830
box -6 -8 86 268
use NAND3X1  _1671_
timestamp 0
transform 1 0 5590 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1672_
timestamp 0
transform -1 0 6210 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1673_
timestamp 0
transform 1 0 5770 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1674_
timestamp 0
transform -1 0 6030 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1675_
timestamp 0
transform 1 0 4070 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1676_
timestamp 0
transform 1 0 5250 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1677_
timestamp 0
transform 1 0 5170 0 -1 2870
box -6 -8 86 268
use DFFSR  _1678_
timestamp 0
transform -1 0 5930 0 -1 1310
box -6 -8 466 268
use DFFSR  _1679_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 466 268
use DFFSR  _1680_
timestamp 0
transform -1 0 5770 0 -1 270
box -6 -8 466 268
use DFFSR  _1681_
timestamp 0
transform 1 0 3470 0 1 1310
box -6 -8 466 268
use DFFSR  _1682_
timestamp 0
transform -1 0 5190 0 -1 790
box -6 -8 466 268
use DFFSR  _1683_
timestamp 0
transform -1 0 3070 0 -1 1830
box -6 -8 466 268
use DFFSR  _1684_
timestamp 0
transform -1 0 2950 0 1 1310
box -6 -8 466 268
use DFFSR  _1685_
timestamp 0
transform -1 0 2430 0 -1 790
box -6 -8 466 268
use DFFSR  _1686_
timestamp 0
transform -1 0 2090 0 -1 270
box -6 -8 466 268
use DFFSR  _1687_
timestamp 0
transform 1 0 2090 0 -1 270
box -6 -8 466 268
use DFFSR  _1688_
timestamp 0
transform 1 0 3050 0 -1 1310
box -6 -8 466 268
use DFFSR  _1689_
timestamp 0
transform -1 0 2610 0 -1 1830
box -6 -8 466 268
use DFFSR  _1690_
timestamp 0
transform 1 0 5010 0 -1 3390
box -6 -8 466 268
use DFFSR  _1691_
timestamp 0
transform 1 0 2990 0 1 1830
box -6 -8 466 268
use DFFSR  _1692_
timestamp 0
transform 1 0 3450 0 1 1830
box -6 -8 466 268
use DFFSR  _1693_
timestamp 0
transform 1 0 4270 0 -1 3390
box -6 -8 466 268
use DFFSR  _1694_
timestamp 0
transform -1 0 5550 0 1 2350
box -6 -8 466 268
use DFFSR  _1695_
timestamp 0
transform -1 0 4950 0 -1 1830
box -6 -8 466 268
use DFFSR  _1696_
timestamp 0
transform -1 0 2930 0 -1 2350
box -6 -8 466 268
use DFFSR  _1697_
timestamp 0
transform -1 0 4050 0 -1 3390
box -6 -8 466 268
use DFFSR  _1698_
timestamp 0
transform -1 0 4010 0 1 3390
box -6 -8 466 268
use DFFSR  _1699_
timestamp 0
transform 1 0 5850 0 -1 790
box -6 -8 466 268
use DFFSR  _1700_
timestamp 0
transform 1 0 5730 0 1 1310
box -6 -8 466 268
use DFFSR  _1701_
timestamp 0
transform 1 0 5930 0 -1 270
box -6 -8 466 268
use DFFSR  _1702_
timestamp 0
transform 1 0 5590 0 1 270
box -6 -8 466 268
use DFFSR  _1703_
timestamp 0
transform 1 0 5750 0 1 2870
box -6 -8 466 268
use DFFSR  _1704_
timestamp 0
transform 1 0 5550 0 1 2350
box -6 -8 466 268
use DFFSR  _1705_
timestamp 0
transform 1 0 5470 0 -1 1830
box -6 -8 466 268
use DFFSR  _1706_
timestamp 0
transform -1 0 5810 0 1 1830
box -6 -8 466 268
use DFFSR  _1707_
timestamp 0
transform 1 0 5770 0 -1 3390
box -6 -8 466 268
use DFFSR  _1708_
timestamp 0
transform 1 0 3070 0 -1 1830
box -6 -8 466 268
use DFFSR  _1709_
timestamp 0
transform -1 0 5590 0 1 1310
box -6 -8 466 268
use DFFSR  _1710_
timestamp 0
transform -1 0 5270 0 1 2870
box -6 -8 466 268
use BUFX2  _1711_
timestamp 0
transform -1 0 170 0 -1 4950
box -6 -8 66 268
use BUFX2  _1712_
timestamp 0
transform -1 0 170 0 1 4950
box -6 -8 66 268
use BUFX2  _1713_
timestamp 0
transform -1 0 1170 0 -1 270
box -6 -8 66 268
use BUFX2  _1714_
timestamp 0
transform 1 0 270 0 -1 6510
box -6 -8 66 268
use BUFX2  _1715_
timestamp 0
transform -1 0 170 0 -1 270
box -6 -8 66 268
use BUFX2  _1716_
timestamp 0
transform -1 0 170 0 1 4430
box -6 -8 66 268
use BUFX2  _1717_
timestamp 0
transform 1 0 430 0 -1 270
box -6 -8 66 268
use BUFX2  _1718_
timestamp 0
transform -1 0 170 0 -1 6510
box -6 -8 66 268
use BUFX2  _1719_
timestamp 0
transform 1 0 1270 0 -1 270
box -6 -8 66 268
use BUFX2  _1720_
timestamp 0
transform -1 0 170 0 1 5470
box -6 -8 66 268
use BUFX2  _1721_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 66 268
use BUFX2  _1722_
timestamp 0
transform -1 0 170 0 1 3910
box -6 -8 66 268
use BUFX2  _1723_
timestamp 0
transform 1 0 1570 0 -1 270
box -6 -8 66 268
use BUFX2  _1724_
timestamp 0
transform 1 0 430 0 -1 6510
box -6 -8 66 268
use BUFX2  _1725_
timestamp 0
transform -1 0 530 0 1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert0
timestamp 0
transform -1 0 170 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 310 0 1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 270 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 430 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 5870 0 -1 270
box -6 -8 66 268
use BUFX2  BUFX2_insert12
timestamp 0
transform -1 0 5490 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 5690 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert14
timestamp 0
transform -1 0 2590 0 1 790
box -6 -8 66 268
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 3410 0 1 1310
box -6 -8 66 268
use CLKBUF1  CLKBUF1_insert4
timestamp 0
transform 1 0 5030 0 1 790
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert5
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert6
timestamp 0
transform -1 0 5010 0 -1 3390
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert7
timestamp 0
transform 1 0 570 0 -1 2350
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 630 0 -1 4430
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform 1 0 2650 0 1 1830
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform -1 0 3790 0 -1 1310
box -6 -8 186 268
use FILL  FILL102150x62550
timestamp 0
transform -1 0 6830 0 -1 4430
box -6 -8 26 268
use FILL  FILL102450x7950
timestamp 0
transform -1 0 6850 0 -1 790
box -6 -8 26 268
use FILL  FILL102450x11850
timestamp 0
transform 1 0 6830 0 1 790
box -6 -8 26 268
use FILL  FILL102450x15750
timestamp 0
transform -1 0 6850 0 -1 1310
box -6 -8 26 268
use FILL  FILL102450x19650
timestamp 0
transform 1 0 6830 0 1 1310
box -6 -8 26 268
use FILL  FILL102450x39150
timestamp 0
transform -1 0 6850 0 -1 2870
box -6 -8 26 268
use FILL  FILL102450x43050
timestamp 0
transform 1 0 6830 0 1 2870
box -6 -8 26 268
use FILL  FILL102450x62550
timestamp 0
transform -1 0 6850 0 -1 4430
box -6 -8 26 268
use FILL  FILL102450x66450
timestamp 0
transform 1 0 6830 0 1 4430
box -6 -8 26 268
use FILL  FILL102450x70350
timestamp 0
transform -1 0 6850 0 -1 4950
box -6 -8 26 268
use FILL  FILL102450x85950
timestamp 0
transform -1 0 6850 0 -1 5990
box -6 -8 26 268
use FILL  FILL102750x7950
timestamp 0
transform -1 0 6870 0 -1 790
box -6 -8 26 268
use FILL  FILL102750x11850
timestamp 0
transform 1 0 6850 0 1 790
box -6 -8 26 268
use FILL  FILL102750x15750
timestamp 0
transform -1 0 6870 0 -1 1310
box -6 -8 26 268
use FILL  FILL102750x19650
timestamp 0
transform 1 0 6850 0 1 1310
box -6 -8 26 268
use FILL  FILL102750x39150
timestamp 0
transform -1 0 6870 0 -1 2870
box -6 -8 26 268
use FILL  FILL102750x43050
timestamp 0
transform 1 0 6850 0 1 2870
box -6 -8 26 268
use FILL  FILL102750x46950
timestamp 0
transform -1 0 6870 0 -1 3390
box -6 -8 26 268
use FILL  FILL102750x62550
timestamp 0
transform -1 0 6870 0 -1 4430
box -6 -8 26 268
use FILL  FILL102750x66450
timestamp 0
transform 1 0 6850 0 1 4430
box -6 -8 26 268
use FILL  FILL102750x70350
timestamp 0
transform -1 0 6870 0 -1 4950
box -6 -8 26 268
use FILL  FILL102750x85950
timestamp 0
transform -1 0 6870 0 -1 5990
box -6 -8 26 268
use FILL  FILL102750x89850
timestamp 0
transform 1 0 6850 0 1 5990
box -6 -8 26 268
use FILL  FILL103050x7950
timestamp 0
transform -1 0 6890 0 -1 790
box -6 -8 26 268
use FILL  FILL103050x11850
timestamp 0
transform 1 0 6870 0 1 790
box -6 -8 26 268
use FILL  FILL103050x15750
timestamp 0
transform -1 0 6890 0 -1 1310
box -6 -8 26 268
use FILL  FILL103050x19650
timestamp 0
transform 1 0 6870 0 1 1310
box -6 -8 26 268
use FILL  FILL103050x31350
timestamp 0
transform -1 0 6890 0 -1 2350
box -6 -8 26 268
use FILL  FILL103050x35250
timestamp 0
transform 1 0 6870 0 1 2350
box -6 -8 26 268
use FILL  FILL103050x39150
timestamp 0
transform -1 0 6890 0 -1 2870
box -6 -8 26 268
use FILL  FILL103050x43050
timestamp 0
transform 1 0 6870 0 1 2870
box -6 -8 26 268
use FILL  FILL103050x46950
timestamp 0
transform -1 0 6890 0 -1 3390
box -6 -8 26 268
use FILL  FILL103050x62550
timestamp 0
transform -1 0 6890 0 -1 4430
box -6 -8 26 268
use FILL  FILL103050x66450
timestamp 0
transform 1 0 6870 0 1 4430
box -6 -8 26 268
use FILL  FILL103050x70350
timestamp 0
transform -1 0 6890 0 -1 4950
box -6 -8 26 268
use FILL  FILL103050x85950
timestamp 0
transform -1 0 6890 0 -1 5990
box -6 -8 26 268
use FILL  FILL103050x89850
timestamp 0
transform 1 0 6870 0 1 5990
box -6 -8 26 268
use FILL  FILL103350x7950
timestamp 0
transform -1 0 6910 0 -1 790
box -6 -8 26 268
use FILL  FILL103350x11850
timestamp 0
transform 1 0 6890 0 1 790
box -6 -8 26 268
use FILL  FILL103350x15750
timestamp 0
transform -1 0 6910 0 -1 1310
box -6 -8 26 268
use FILL  FILL103350x19650
timestamp 0
transform 1 0 6890 0 1 1310
box -6 -8 26 268
use FILL  FILL103350x31350
timestamp 0
transform -1 0 6910 0 -1 2350
box -6 -8 26 268
use FILL  FILL103350x35250
timestamp 0
transform 1 0 6890 0 1 2350
box -6 -8 26 268
use FILL  FILL103350x39150
timestamp 0
transform -1 0 6910 0 -1 2870
box -6 -8 26 268
use FILL  FILL103350x43050
timestamp 0
transform 1 0 6890 0 1 2870
box -6 -8 26 268
use FILL  FILL103350x46950
timestamp 0
transform -1 0 6910 0 -1 3390
box -6 -8 26 268
use FILL  FILL103350x58650
timestamp 0
transform 1 0 6890 0 1 3910
box -6 -8 26 268
use FILL  FILL103350x62550
timestamp 0
transform -1 0 6910 0 -1 4430
box -6 -8 26 268
use FILL  FILL103350x66450
timestamp 0
transform 1 0 6890 0 1 4430
box -6 -8 26 268
use FILL  FILL103350x70350
timestamp 0
transform -1 0 6910 0 -1 4950
box -6 -8 26 268
use FILL  FILL103350x85950
timestamp 0
transform -1 0 6910 0 -1 5990
box -6 -8 26 268
use FILL  FILL103350x89850
timestamp 0
transform 1 0 6890 0 1 5990
box -6 -8 26 268
use FILL  FILL103650x7950
timestamp 0
transform -1 0 6930 0 -1 790
box -6 -8 26 268
use FILL  FILL103650x11850
timestamp 0
transform 1 0 6910 0 1 790
box -6 -8 26 268
use FILL  FILL103650x15750
timestamp 0
transform -1 0 6930 0 -1 1310
box -6 -8 26 268
use FILL  FILL103650x19650
timestamp 0
transform 1 0 6910 0 1 1310
box -6 -8 26 268
use FILL  FILL103650x27450
timestamp 0
transform 1 0 6910 0 1 1830
box -6 -8 26 268
use FILL  FILL103650x31350
timestamp 0
transform -1 0 6930 0 -1 2350
box -6 -8 26 268
use FILL  FILL103650x35250
timestamp 0
transform 1 0 6910 0 1 2350
box -6 -8 26 268
use FILL  FILL103650x39150
timestamp 0
transform -1 0 6930 0 -1 2870
box -6 -8 26 268
use FILL  FILL103650x43050
timestamp 0
transform 1 0 6910 0 1 2870
box -6 -8 26 268
use FILL  FILL103650x46950
timestamp 0
transform -1 0 6930 0 -1 3390
box -6 -8 26 268
use FILL  FILL103650x58650
timestamp 0
transform 1 0 6910 0 1 3910
box -6 -8 26 268
use FILL  FILL103650x62550
timestamp 0
transform -1 0 6930 0 -1 4430
box -6 -8 26 268
use FILL  FILL103650x66450
timestamp 0
transform 1 0 6910 0 1 4430
box -6 -8 26 268
use FILL  FILL103650x70350
timestamp 0
transform -1 0 6930 0 -1 4950
box -6 -8 26 268
use FILL  FILL103650x85950
timestamp 0
transform -1 0 6930 0 -1 5990
box -6 -8 26 268
use FILL  FILL103650x89850
timestamp 0
transform 1 0 6910 0 1 5990
box -6 -8 26 268
use FILL  FILL103650x93750
timestamp 0
transform -1 0 6930 0 -1 6510
box -6 -8 26 268
use FILL  FILL103950x4050
timestamp 0
transform 1 0 6930 0 1 270
box -6 -8 26 268
use FILL  FILL103950x7950
timestamp 0
transform -1 0 6950 0 -1 790
box -6 -8 26 268
use FILL  FILL103950x11850
timestamp 0
transform 1 0 6930 0 1 790
box -6 -8 26 268
use FILL  FILL103950x15750
timestamp 0
transform -1 0 6950 0 -1 1310
box -6 -8 26 268
use FILL  FILL103950x19650
timestamp 0
transform 1 0 6930 0 1 1310
box -6 -8 26 268
use FILL  FILL103950x27450
timestamp 0
transform 1 0 6930 0 1 1830
box -6 -8 26 268
use FILL  FILL103950x31350
timestamp 0
transform -1 0 6950 0 -1 2350
box -6 -8 26 268
use FILL  FILL103950x35250
timestamp 0
transform 1 0 6930 0 1 2350
box -6 -8 26 268
use FILL  FILL103950x39150
timestamp 0
transform -1 0 6950 0 -1 2870
box -6 -8 26 268
use FILL  FILL103950x43050
timestamp 0
transform 1 0 6930 0 1 2870
box -6 -8 26 268
use FILL  FILL103950x46950
timestamp 0
transform -1 0 6950 0 -1 3390
box -6 -8 26 268
use FILL  FILL103950x50850
timestamp 0
transform 1 0 6930 0 1 3390
box -6 -8 26 268
use FILL  FILL103950x54750
timestamp 0
transform -1 0 6950 0 -1 3910
box -6 -8 26 268
use FILL  FILL103950x58650
timestamp 0
transform 1 0 6930 0 1 3910
box -6 -8 26 268
use FILL  FILL103950x62550
timestamp 0
transform -1 0 6950 0 -1 4430
box -6 -8 26 268
use FILL  FILL103950x66450
timestamp 0
transform 1 0 6930 0 1 4430
box -6 -8 26 268
use FILL  FILL103950x70350
timestamp 0
transform -1 0 6950 0 -1 4950
box -6 -8 26 268
use FILL  FILL103950x74250
timestamp 0
transform 1 0 6930 0 1 4950
box -6 -8 26 268
use FILL  FILL103950x85950
timestamp 0
transform -1 0 6950 0 -1 5990
box -6 -8 26 268
use FILL  FILL103950x89850
timestamp 0
transform 1 0 6930 0 1 5990
box -6 -8 26 268
use FILL  FILL103950x93750
timestamp 0
transform -1 0 6950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__828_
timestamp 0
transform 1 0 790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__829_
timestamp 0
transform 1 0 1470 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__830_
timestamp 0
transform -1 0 2330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__831_
timestamp 0
transform -1 0 1310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__832_
timestamp 0
transform 1 0 2230 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__833_
timestamp 0
transform 1 0 1930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__834_
timestamp 0
transform -1 0 1550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__835_
timestamp 0
transform -1 0 1630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__836_
timestamp 0
transform -1 0 950 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__837_
timestamp 0
transform 1 0 830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__838_
timestamp 0
transform -1 0 670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__839_
timestamp 0
transform -1 0 870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__840_
timestamp 0
transform 1 0 10 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__841_
timestamp 0
transform -1 0 30 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__842_
timestamp 0
transform 1 0 10 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__843_
timestamp 0
transform -1 0 190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__844_
timestamp 0
transform 1 0 650 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__845_
timestamp 0
transform 1 0 190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__846_
timestamp 0
transform -1 0 710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__847_
timestamp 0
transform -1 0 870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__848_
timestamp 0
transform -1 0 530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__849_
timestamp 0
transform 1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__850_
timestamp 0
transform -1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__851_
timestamp 0
transform -1 0 830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__852_
timestamp 0
transform -1 0 650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__853_
timestamp 0
transform 1 0 530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__854_
timestamp 0
transform -1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__855_
timestamp 0
transform -1 0 510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__856_
timestamp 0
transform -1 0 710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__857_
timestamp 0
transform 1 0 970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__858_
timestamp 0
transform -1 0 450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__859_
timestamp 0
transform 1 0 10 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__860_
timestamp 0
transform 1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__861_
timestamp 0
transform 1 0 790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__862_
timestamp 0
transform -1 0 670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__863_
timestamp 0
transform -1 0 490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__864_
timestamp 0
transform 1 0 790 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__865_
timestamp 0
transform 1 0 370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__866_
timestamp 0
transform -1 0 1330 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__867_
timestamp 0
transform 1 0 950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__868_
timestamp 0
transform 1 0 970 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__869_
timestamp 0
transform -1 0 1170 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__870_
timestamp 0
transform 1 0 1090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__871_
timestamp 0
transform -1 0 1390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__872_
timestamp 0
transform -1 0 830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__873_
timestamp 0
transform 1 0 990 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__874_
timestamp 0
transform 1 0 970 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__875_
timestamp 0
transform 1 0 1210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__876_
timestamp 0
transform -1 0 1130 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__877_
timestamp 0
transform 1 0 1270 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__878_
timestamp 0
transform -1 0 810 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__879_
timestamp 0
transform -1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__880_
timestamp 0
transform 1 0 1130 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__881_
timestamp 0
transform 1 0 170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__882_
timestamp 0
transform -1 0 170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__883_
timestamp 0
transform 1 0 810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__884_
timestamp 0
transform -1 0 970 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__885_
timestamp 0
transform -1 0 990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__886_
timestamp 0
transform -1 0 810 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__887_
timestamp 0
transform 1 0 810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__888_
timestamp 0
transform -1 0 630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__889_
timestamp 0
transform 1 0 470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__890_
timestamp 0
transform -1 0 650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__891_
timestamp 0
transform 1 0 290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__892_
timestamp 0
transform -1 0 470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__893_
timestamp 0
transform -1 0 170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__894_
timestamp 0
transform -1 0 490 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__895_
timestamp 0
transform -1 0 650 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__896_
timestamp 0
transform 1 0 1770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__897_
timestamp 0
transform -1 0 2490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__898_
timestamp 0
transform -1 0 2150 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__899_
timestamp 0
transform 1 0 2090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__900_
timestamp 0
transform -1 0 1710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__901_
timestamp 0
transform 1 0 1590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__902_
timestamp 0
transform -1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__903_
timestamp 0
transform -1 0 1770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__904_
timestamp 0
transform -1 0 1450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__905_
timestamp 0
transform -1 0 1370 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__906_
timestamp 0
transform 1 0 1170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__907_
timestamp 0
transform 1 0 1750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__908_
timestamp 0
transform 1 0 2250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__909_
timestamp 0
transform 1 0 1970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__910_
timestamp 0
transform -1 0 1810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__911_
timestamp 0
transform 1 0 1570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__912_
timestamp 0
transform -1 0 1710 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__913_
timestamp 0
transform 1 0 2810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__914_
timestamp 0
transform -1 0 3150 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__915_
timestamp 0
transform 1 0 2070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__916_
timestamp 0
transform -1 0 2070 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__917_
timestamp 0
transform 1 0 1510 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__918_
timestamp 0
transform 1 0 1910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__919_
timestamp 0
transform -1 0 2970 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__920_
timestamp 0
transform -1 0 3230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__921_
timestamp 0
transform 1 0 2610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform -1 0 2450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform -1 0 2270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform 1 0 1870 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform 1 0 2550 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform -1 0 2710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform -1 0 3370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform -1 0 3050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform -1 0 2530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform -1 0 2350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform -1 0 890 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform -1 0 2870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform -1 0 2810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform -1 0 2390 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform -1 0 710 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform -1 0 1150 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform -1 0 650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform 1 0 1790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform -1 0 1190 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 1650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform 1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform 1 0 950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform -1 0 350 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform -1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform 1 0 2010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform 1 0 1490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform 1 0 1670 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform 1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform -1 0 2970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform -1 0 6030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform -1 0 6350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform 1 0 5850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform -1 0 5690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform 1 0 5350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform 1 0 3190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform 1 0 2870 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform -1 0 6470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform 1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform 1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform -1 0 5390 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform 1 0 5210 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform 1 0 3450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform -1 0 3470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform -1 0 5270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform 1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform -1 0 4070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform -1 0 3210 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform -1 0 3910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform 1 0 3590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform -1 0 4430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform 1 0 2850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform -1 0 6310 0 1 790
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform -1 0 6190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform 1 0 5950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform 1 0 6130 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform 1 0 4170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform 1 0 4230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform -1 0 4210 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform 1 0 5510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform 1 0 6010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform -1 0 6770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 5950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform -1 0 5790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform -1 0 5630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform -1 0 4730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform 1 0 5950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 5510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform -1 0 5430 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform -1 0 5730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform -1 0 5570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 5090 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform 1 0 4890 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform 1 0 4650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 4810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform -1 0 5290 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 5470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform 1 0 5330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform -1 0 4750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 4590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 5230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform -1 0 5130 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 3850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform 1 0 3670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 2950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform -1 0 2630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform -1 0 4030 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform 1 0 3610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 2870 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform 1 0 6230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 4810 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform 1 0 3730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 6850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 4530 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform 1 0 4030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 3830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform -1 0 4390 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform -1 0 4210 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform 1 0 6350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform 1 0 3890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform -1 0 4490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform -1 0 4650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 3970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform -1 0 4150 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 4310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform 1 0 3670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform -1 0 4370 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform -1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 4170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform -1 0 4010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 3750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform -1 0 3450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 4550 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform -1 0 4030 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 3670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform -1 0 3810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 3870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 3670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 3510 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 3030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform 1 0 3350 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 3530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform -1 0 3390 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform 1 0 490 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform 1 0 1050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform -1 0 910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform -1 0 1010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform -1 0 850 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform -1 0 1290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform 1 0 2370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 3210 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform -1 0 3030 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform -1 0 2710 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform 1 0 1450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 1350 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 1170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform -1 0 3130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform -1 0 2790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform -1 0 2650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 1830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform -1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform 1 0 1450 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 1490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform 1 0 1010 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 1490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 1170 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 1290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 910 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 10 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform -1 0 350 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 10 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 870 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 1150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform 1 0 690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform -1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform 1 0 10 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform -1 0 1870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 2410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform 1 0 2010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform -1 0 2230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 1130 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform -1 0 830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform 1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 570 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform -1 0 670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 490 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform -1 0 250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform -1 0 190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform 1 0 150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform 1 0 2110 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform -1 0 2270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform 1 0 1950 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 2170 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 1610 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform 1 0 1790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 1690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform 1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 1450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform 1 0 1490 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform -1 0 1670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform -1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform -1 0 2050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform -1 0 1870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform -1 0 1670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 1150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform -1 0 1330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform -1 0 1010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform -1 0 550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform -1 0 390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform -1 0 3830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 4030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform 1 0 5470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform 1 0 6490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform -1 0 5470 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 4750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 4950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform -1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform 1 0 5630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform -1 0 5150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform -1 0 5130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 4410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform -1 0 4250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform -1 0 6310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform -1 0 6730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform 1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform 1 0 3490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 6090 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform 1 0 5290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform 1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform 1 0 4150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform 1 0 4790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform 1 0 5030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform 1 0 5050 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform -1 0 4810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform -1 0 5910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform 1 0 5770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 3810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 3090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 2850 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform -1 0 3030 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 3490 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 3650 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform -1 0 3990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform 1 0 4310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 4990 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform 1 0 5290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform 1 0 4690 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 5230 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform 1 0 5130 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform -1 0 5350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 5130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform -1 0 4510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform -1 0 5530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 5110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform -1 0 4770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 4470 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform 1 0 5650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform 1 0 6110 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform 1 0 4230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 4290 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform -1 0 3610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform 1 0 3630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform 1 0 3450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 3090 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform 1 0 3350 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform -1 0 3350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform -1 0 2170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 3510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 3330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 3190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform 1 0 2490 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform 1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 2070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform 1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform 1 0 2210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 3050 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 2870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform 1 0 4430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 4590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform 1 0 4070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform -1 0 3970 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform 1 0 4650 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 4110 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform -1 0 3810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform -1 0 3110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 3730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform -1 0 3310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 3290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform -1 0 3430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 3550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform -1 0 3650 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform -1 0 3910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 3250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform -1 0 3310 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 3470 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 2750 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 2330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform 1 0 1910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 1830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform -1 0 2170 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform 1 0 2430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform -1 0 2630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 2790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform -1 0 1570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 1770 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 1830 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform -1 0 2350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform -1 0 1950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform 1 0 2110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 1250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform -1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 1570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform -1 0 2690 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 2490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 1470 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform -1 0 1410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 1650 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 1990 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 2030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform 1 0 1750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform 1 0 1830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform -1 0 1650 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 2190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 2030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform 1 0 1790 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform -1 0 1410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform -1 0 1330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform 1 0 1930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 2170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform -1 0 2010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 1650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 1970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform -1 0 2190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform 1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform -1 0 2330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 2350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform 1 0 1970 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform -1 0 2570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform -1 0 230 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform 1 0 10 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 350 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform -1 0 730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform 1 0 350 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 170 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 870 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 690 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 1490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 1170 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 1250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 1270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform 1 0 1850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 1070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform -1 0 1090 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 490 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform -1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform -1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform 1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform -1 0 750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 1690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 1430 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform -1 0 930 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 1610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 2090 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform 1 0 1910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform 1 0 2130 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform -1 0 2530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform -1 0 1490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform -1 0 1330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform 1 0 1310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 1290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform -1 0 5190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform 1 0 2890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform 1 0 2530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform 1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 1650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform 1 0 2710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform -1 0 4930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 5590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 5470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 5750 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform -1 0 5650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 6330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 6630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 6690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 6690 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform 1 0 4950 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform -1 0 5430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform 1 0 5470 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform 1 0 5650 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform 1 0 5830 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 5370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 6370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform -1 0 5730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 5870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform -1 0 6110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform 1 0 6330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform 1 0 6490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform -1 0 6670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform -1 0 6670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform -1 0 6770 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform 1 0 6430 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 6790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 5550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 6510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 6690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 6570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform 1 0 6510 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 5770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform 1 0 6270 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform -1 0 6510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform 1 0 6450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 5450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform 1 0 5670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform -1 0 5850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform 1 0 6010 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 6310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform 1 0 6490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 6150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 5950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 6410 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 6030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform -1 0 6210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform -1 0 6650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform 1 0 6590 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 6670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 6770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 6010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform -1 0 6170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 5290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform -1 0 4490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform 1 0 3810 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform 1 0 4150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 4630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform 1 0 5750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 5310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 6470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 6790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 6550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 6610 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform 1 0 6110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform -1 0 6310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 5590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform 1 0 4730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform -1 0 4910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform -1 0 5150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform -1 0 4950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform -1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 4230 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform -1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform -1 0 1850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform -1 0 1310 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform -1 0 1330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform -1 0 830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform 1 0 890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform -1 0 4070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 2950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform 1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 4290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 4430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform 1 0 5930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 5850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 4390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform 1 0 4690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform 1 0 4530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform 1 0 4830 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 4870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform -1 0 5070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 4990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform -1 0 5010 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform 1 0 4270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform -1 0 6030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 5290 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 6170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform -1 0 6510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform -1 0 6210 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform -1 0 6350 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform -1 0 5430 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 4970 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform -1 0 4350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform -1 0 4730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 4550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform -1 0 4550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform 1 0 3950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform -1 0 4170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform 1 0 530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform 1 0 2310 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform -1 0 3990 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform -1 0 4650 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 4830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform -1 0 4650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 4830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 2330 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform 1 0 4630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform -1 0 2210 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 2290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform 1 0 2350 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform 1 0 2610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform 1 0 2930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 2790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform 1 0 2690 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 2150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 1630 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform 1 0 1670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform 1 0 2330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform 1 0 2450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 2830 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform 1 0 4310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform 1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1452_
timestamp 0
transform 1 0 2770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1453_
timestamp 0
transform 1 0 2590 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1454_
timestamp 0
transform -1 0 2770 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1455_
timestamp 0
transform -1 0 5210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1456_
timestamp 0
transform 1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1457_
timestamp 0
transform -1 0 5370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1458_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1459_
timestamp 0
transform 1 0 3610 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 4370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 3430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1462_
timestamp 0
transform -1 0 3070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1463_
timestamp 0
transform 1 0 2730 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1464_
timestamp 0
transform 1 0 2170 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 2470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1466_
timestamp 0
transform -1 0 2650 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1467_
timestamp 0
transform 1 0 2950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1468_
timestamp 0
transform 1 0 3090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1469_
timestamp 0
transform 1 0 2550 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1470_
timestamp 0
transform 1 0 3550 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1471_
timestamp 0
transform -1 0 3790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1472_
timestamp 0
transform -1 0 3750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1473_
timestamp 0
transform 1 0 3990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1474_
timestamp 0
transform 1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1475_
timestamp 0
transform -1 0 4190 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1476_
timestamp 0
transform -1 0 4770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1477_
timestamp 0
transform 1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1478_
timestamp 0
transform -1 0 4590 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1479_
timestamp 0
transform -1 0 4350 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1480_
timestamp 0
transform 1 0 5930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 5770 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1482_
timestamp 0
transform -1 0 5570 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1483_
timestamp 0
transform 1 0 3550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 2810 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1485_
timestamp 0
transform 1 0 2970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1486_
timestamp 0
transform 1 0 3410 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1487_
timestamp 0
transform 1 0 3250 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 2930 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 2890 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1490_
timestamp 0
transform -1 0 3230 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 4650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1492_
timestamp 0
transform -1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1493_
timestamp 0
transform -1 0 3990 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1494_
timestamp 0
transform 1 0 3470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1495_
timestamp 0
transform 1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1496_
timestamp 0
transform -1 0 4390 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1497_
timestamp 0
transform 1 0 4910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 4410 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1499_
timestamp 0
transform 1 0 4230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1500_
timestamp 0
transform -1 0 3910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1501_
timestamp 0
transform 1 0 4050 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1502_
timestamp 0
transform 1 0 4150 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1503_
timestamp 0
transform 1 0 4150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1504_
timestamp 0
transform -1 0 4470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1505_
timestamp 0
transform -1 0 4110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1506_
timestamp 0
transform 1 0 4310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 4550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1508_
timestamp 0
transform 1 0 4750 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1509_
timestamp 0
transform 1 0 2150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1510_
timestamp 0
transform -1 0 2550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1511_
timestamp 0
transform 1 0 2330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1512_
timestamp 0
transform 1 0 2450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1513_
timestamp 0
transform -1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1514_
timestamp 0
transform -1 0 2530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1515_
timestamp 0
transform 1 0 2630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1516_
timestamp 0
transform -1 0 2810 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1517_
timestamp 0
transform 1 0 3690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1518_
timestamp 0
transform 1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1519_
timestamp 0
transform -1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1520_
timestamp 0
transform 1 0 3130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1521_
timestamp 0
transform -1 0 3950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1522_
timestamp 0
transform -1 0 3810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 2950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1524_
timestamp 0
transform -1 0 4010 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1525_
timestamp 0
transform 1 0 3130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1526_
timestamp 0
transform 1 0 3290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 2930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1528_
timestamp 0
transform -1 0 2970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1529_
timestamp 0
transform -1 0 1210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 1350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 1490 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1532_
timestamp 0
transform -1 0 1850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 2010 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 2310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 2690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1536_
timestamp 0
transform -1 0 3310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1537_
timestamp 0
transform 1 0 2430 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1538_
timestamp 0
transform 1 0 3830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1539_
timestamp 0
transform -1 0 3210 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1540_
timestamp 0
transform 1 0 1770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1541_
timestamp 0
transform -1 0 3390 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1542_
timestamp 0
transform 1 0 1970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1543_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1544_
timestamp 0
transform 1 0 3090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1545_
timestamp 0
transform 1 0 2390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 3530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1547_
timestamp 0
transform 1 0 4690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1548_
timestamp 0
transform 1 0 3830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1549_
timestamp 0
transform -1 0 4830 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1550_
timestamp 0
transform 1 0 4950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1551_
timestamp 0
transform -1 0 5150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1552_
timestamp 0
transform 1 0 4390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1553_
timestamp 0
transform -1 0 4470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1554_
timestamp 0
transform 1 0 5170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1555_
timestamp 0
transform 1 0 4970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1556_
timestamp 0
transform -1 0 4990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1557_
timestamp 0
transform -1 0 4790 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1558_
timestamp 0
transform -1 0 3770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1559_
timestamp 0
transform 1 0 4910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1560_
timestamp 0
transform -1 0 4950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1561_
timestamp 0
transform -1 0 4590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1562_
timestamp 0
transform 1 0 3910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 4110 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1564_
timestamp 0
transform -1 0 4810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 3490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1566_
timestamp 0
transform 1 0 3430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1567_
timestamp 0
transform -1 0 2950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1568_
timestamp 0
transform 1 0 3590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 3250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1570_
timestamp 0
transform 1 0 3070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1571_
timestamp 0
transform 1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1572_
timestamp 0
transform 1 0 3310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1573_
timestamp 0
transform 1 0 3870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1574_
timestamp 0
transform -1 0 4410 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1575_
timestamp 0
transform -1 0 3910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1576_
timestamp 0
transform -1 0 4070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1577_
timestamp 0
transform -1 0 3390 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1578_
timestamp 0
transform -1 0 3750 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1579_
timestamp 0
transform 1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 3630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 3830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1582_
timestamp 0
transform 1 0 4270 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 4010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1584_
timestamp 0
transform -1 0 4570 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1585_
timestamp 0
transform 1 0 4170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1586_
timestamp 0
transform -1 0 4650 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1587_
timestamp 0
transform -1 0 3230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1588_
timestamp 0
transform -1 0 3090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 4390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1590_
timestamp 0
transform -1 0 4250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1591_
timestamp 0
transform 1 0 4210 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1592_
timestamp 0
transform 1 0 4050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1593_
timestamp 0
transform 1 0 2570 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1594_
timestamp 0
transform 1 0 2750 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1595_
timestamp 0
transform -1 0 2950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1596_
timestamp 0
transform -1 0 3150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1597_
timestamp 0
transform 1 0 2950 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1598_
timestamp 0
transform -1 0 3310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1599_
timestamp 0
transform -1 0 3650 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1600_
timestamp 0
transform 1 0 3450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1601_
timestamp 0
transform -1 0 3390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1602_
timestamp 0
transform -1 0 2850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1603_
timestamp 0
transform -1 0 3030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1604_
timestamp 0
transform -1 0 3210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 4050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1606_
timestamp 0
transform 1 0 6270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1607_
timestamp 0
transform 1 0 6210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1608_
timestamp 0
transform -1 0 6390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1609_
timestamp 0
transform 1 0 6150 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1610_
timestamp 0
transform 1 0 6550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1611_
timestamp 0
transform 1 0 5590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1612_
timestamp 0
transform -1 0 6810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1613_
timestamp 0
transform -1 0 6430 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1614_
timestamp 0
transform -1 0 6250 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1615_
timestamp 0
transform -1 0 6070 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1616_
timestamp 0
transform 1 0 5870 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1617_
timestamp 0
transform 1 0 5610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1618_
timestamp 0
transform -1 0 5410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1619_
timestamp 0
transform 1 0 5310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1620_
timestamp 0
transform -1 0 6090 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1621_
timestamp 0
transform 1 0 5310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1622_
timestamp 0
transform 1 0 6730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1623_
timestamp 0
transform 1 0 6390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1624_
timestamp 0
transform -1 0 6790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1625_
timestamp 0
transform -1 0 6530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1626_
timestamp 0
transform 1 0 6510 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1627_
timestamp 0
transform 1 0 6350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1628_
timestamp 0
transform -1 0 6150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1629_
timestamp 0
transform 1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1630_
timestamp 0
transform 1 0 6650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1631_
timestamp 0
transform -1 0 6710 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1632_
timestamp 0
transform -1 0 6590 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1633_
timestamp 0
transform -1 0 6610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1634_
timestamp 0
transform -1 0 6430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1635_
timestamp 0
transform 1 0 6230 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1636_
timestamp 0
transform -1 0 6410 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1637_
timestamp 0
transform 1 0 6050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1638_
timestamp 0
transform -1 0 6450 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1639_
timestamp 0
transform 1 0 6310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 5650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1641_
timestamp 0
transform -1 0 6710 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1642_
timestamp 0
transform -1 0 6210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1643_
timestamp 0
transform -1 0 6510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1644_
timestamp 0
transform -1 0 6210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1645_
timestamp 0
transform 1 0 6530 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1646_
timestamp 0
transform -1 0 6670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1647_
timestamp 0
transform -1 0 5990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1648_
timestamp 0
transform 1 0 5770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1649_
timestamp 0
transform -1 0 6670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1650_
timestamp 0
transform -1 0 6670 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1651_
timestamp 0
transform -1 0 6230 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1652_
timestamp 0
transform -1 0 6450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1653_
timestamp 0
transform 1 0 5570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1654_
timestamp 0
transform 1 0 6350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1655_
timestamp 0
transform 1 0 6330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1656_
timestamp 0
transform 1 0 6510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1657_
timestamp 0
transform -1 0 6770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 6110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1659_
timestamp 0
transform -1 0 6810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1660_
timestamp 0
transform -1 0 6590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1661_
timestamp 0
transform -1 0 6770 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1662_
timestamp 0
transform -1 0 6410 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1663_
timestamp 0
transform 1 0 5990 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1664_
timestamp 0
transform 1 0 6170 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1665_
timestamp 0
transform -1 0 6290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1666_
timestamp 0
transform -1 0 6610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1667_
timestamp 0
transform 1 0 6370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1668_
timestamp 0
transform 1 0 6670 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1669_
timestamp 0
transform -1 0 5950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1670_
timestamp 0
transform 1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1671_
timestamp 0
transform 1 0 5490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1672_
timestamp 0
transform -1 0 6050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1673_
timestamp 0
transform 1 0 5670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1674_
timestamp 0
transform -1 0 5870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1675_
timestamp 0
transform 1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1676_
timestamp 0
transform 1 0 5150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1677_
timestamp 0
transform 1 0 5070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1711_
timestamp 0
transform -1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1712_
timestamp 0
transform -1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 1030 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1714_
timestamp 0
transform 1 0 170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1715_
timestamp 0
transform -1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1716_
timestamp 0
transform -1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1717_
timestamp 0
transform 1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1718_
timestamp 0
transform -1 0 30 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1719_
timestamp 0
transform 1 0 1170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1721_
timestamp 0
transform -1 0 190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1722_
timestamp 0
transform -1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 1470 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1724_
timestamp 0
transform 1 0 330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_0__1725_
timestamp 0
transform -1 0 390 0 1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform -1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 210 0 1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 5770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform -1 0 5350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 5590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform -1 0 2450 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 3310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert4
timestamp 0
transform 1 0 4930 0 1 790
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert5
timestamp 0
transform -1 0 1890 0 1 4950
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert6
timestamp 0
transform -1 0 4750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert7
timestamp 0
transform 1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert8
timestamp 0
transform -1 0 370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert9
timestamp 0
transform 1 0 2550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert10
timestamp 0
transform -1 0 3530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__828_
timestamp 0
transform 1 0 810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__829_
timestamp 0
transform 1 0 1490 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__830_
timestamp 0
transform -1 0 2350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__831_
timestamp 0
transform -1 0 1330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__832_
timestamp 0
transform 1 0 2250 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__833_
timestamp 0
transform 1 0 1950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__834_
timestamp 0
transform -1 0 1570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__835_
timestamp 0
transform -1 0 1650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__836_
timestamp 0
transform -1 0 970 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__837_
timestamp 0
transform 1 0 850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__838_
timestamp 0
transform -1 0 690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__839_
timestamp 0
transform -1 0 890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__840_
timestamp 0
transform 1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__841_
timestamp 0
transform -1 0 50 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__842_
timestamp 0
transform 1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__843_
timestamp 0
transform -1 0 210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__844_
timestamp 0
transform 1 0 670 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__845_
timestamp 0
transform 1 0 210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__846_
timestamp 0
transform -1 0 730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__847_
timestamp 0
transform -1 0 890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__848_
timestamp 0
transform -1 0 550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__849_
timestamp 0
transform 1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__850_
timestamp 0
transform -1 0 210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__851_
timestamp 0
transform -1 0 850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__852_
timestamp 0
transform -1 0 670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__853_
timestamp 0
transform 1 0 550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__854_
timestamp 0
transform -1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__855_
timestamp 0
transform -1 0 530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__856_
timestamp 0
transform -1 0 730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__857_
timestamp 0
transform 1 0 990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__858_
timestamp 0
transform -1 0 470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__859_
timestamp 0
transform 1 0 30 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__860_
timestamp 0
transform 1 0 1050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__861_
timestamp 0
transform 1 0 810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__862_
timestamp 0
transform -1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__863_
timestamp 0
transform -1 0 510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__864_
timestamp 0
transform 1 0 810 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__865_
timestamp 0
transform 1 0 390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__866_
timestamp 0
transform -1 0 1350 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__867_
timestamp 0
transform 1 0 970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__868_
timestamp 0
transform 1 0 990 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__869_
timestamp 0
transform -1 0 1190 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__870_
timestamp 0
transform 1 0 1110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__871_
timestamp 0
transform -1 0 1410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__872_
timestamp 0
transform -1 0 850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__873_
timestamp 0
transform 1 0 1010 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__874_
timestamp 0
transform 1 0 990 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__875_
timestamp 0
transform 1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__876_
timestamp 0
transform -1 0 1150 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__877_
timestamp 0
transform 1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__878_
timestamp 0
transform -1 0 830 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__879_
timestamp 0
transform -1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__880_
timestamp 0
transform 1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__881_
timestamp 0
transform 1 0 190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__882_
timestamp 0
transform -1 0 190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__883_
timestamp 0
transform 1 0 830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__884_
timestamp 0
transform -1 0 990 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__885_
timestamp 0
transform -1 0 1010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__886_
timestamp 0
transform -1 0 830 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__887_
timestamp 0
transform 1 0 830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__888_
timestamp 0
transform -1 0 650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__889_
timestamp 0
transform 1 0 490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__890_
timestamp 0
transform -1 0 670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__891_
timestamp 0
transform 1 0 310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__892_
timestamp 0
transform -1 0 490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__893_
timestamp 0
transform -1 0 190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__894_
timestamp 0
transform -1 0 510 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__895_
timestamp 0
transform -1 0 670 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__896_
timestamp 0
transform 1 0 1790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__897_
timestamp 0
transform -1 0 2510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__898_
timestamp 0
transform -1 0 2170 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__899_
timestamp 0
transform 1 0 2110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__900_
timestamp 0
transform -1 0 1730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__901_
timestamp 0
transform 1 0 1610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__902_
timestamp 0
transform -1 0 1650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__903_
timestamp 0
transform -1 0 1790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__904_
timestamp 0
transform -1 0 1470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__905_
timestamp 0
transform -1 0 1390 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__906_
timestamp 0
transform 1 0 1190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__907_
timestamp 0
transform 1 0 1770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__908_
timestamp 0
transform 1 0 2270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__909_
timestamp 0
transform 1 0 1990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__910_
timestamp 0
transform -1 0 1830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__911_
timestamp 0
transform 1 0 1590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__912_
timestamp 0
transform -1 0 1730 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__913_
timestamp 0
transform 1 0 2830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__914_
timestamp 0
transform -1 0 3170 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__915_
timestamp 0
transform 1 0 2090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__916_
timestamp 0
transform -1 0 2090 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__917_
timestamp 0
transform 1 0 1530 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__918_
timestamp 0
transform 1 0 1930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__919_
timestamp 0
transform -1 0 2990 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__920_
timestamp 0
transform -1 0 3250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__921_
timestamp 0
transform 1 0 2630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform -1 0 2470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform -1 0 2290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform 1 0 1890 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform 1 0 2570 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform -1 0 2730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform -1 0 3390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform -1 0 3070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform -1 0 2550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform -1 0 2370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform -1 0 910 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform -1 0 2890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform -1 0 2830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform -1 0 2410 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform -1 0 730 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform -1 0 1170 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform -1 0 670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform 1 0 1810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform -1 0 1210 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 1670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform 1 0 1470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform 1 0 970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform -1 0 370 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform -1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform 1 0 2030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform 1 0 1510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform 1 0 1690 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform 1 0 1530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform -1 0 2990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform -1 0 6050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform -1 0 6370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform 1 0 5870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform -1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform 1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform 1 0 3210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform 1 0 2890 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform -1 0 6490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform 1 0 5730 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform 1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform -1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform 1 0 5230 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform 1 0 3470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform -1 0 3490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform -1 0 5290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform 1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform -1 0 4090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform -1 0 3230 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform -1 0 3930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform 1 0 3610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform -1 0 4450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform 1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform -1 0 6330 0 1 790
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform -1 0 6210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform 1 0 5970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform 1 0 6150 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform 1 0 4190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform 1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform -1 0 4230 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform 1 0 5530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform 1 0 6030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform -1 0 6790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 5970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform -1 0 5810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform -1 0 5650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform -1 0 4750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform 1 0 5970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 5530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform -1 0 5450 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform -1 0 5750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform -1 0 5590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 5110 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform 1 0 4910 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform 1 0 4670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 4830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform -1 0 5310 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 5490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform 1 0 5350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform -1 0 4770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 4610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 5250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform -1 0 5150 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 3870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform 1 0 3690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 2970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform -1 0 2650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform -1 0 4050 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform 1 0 3630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 2890 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform 1 0 6250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 4830 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform 1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 6870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 4550 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform 1 0 4050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 3850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform -1 0 4410 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform -1 0 4230 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform 1 0 6370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform 1 0 3910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform -1 0 4510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform -1 0 4670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 3990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform -1 0 4170 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 4330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform 1 0 3690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform -1 0 4390 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform -1 0 2590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 4190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform -1 0 4030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 3770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 3270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform -1 0 3470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 4570 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform -1 0 4050 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 3690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform -1 0 3830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 3890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 3690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform -1 0 3530 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 3050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform 1 0 3370 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 3550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform -1 0 3410 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform 1 0 510 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform 1 0 1070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform -1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform -1 0 1030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform -1 0 870 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform -1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform 1 0 2390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 3230 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform -1 0 3050 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform -1 0 2730 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform 1 0 1470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 1370 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform 1 0 1190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform -1 0 3150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform -1 0 2810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform -1 0 2670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 1850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform -1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform 1 0 1470 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 1510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform 1 0 1030 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 1510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 1190 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform 1 0 1310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform -1 0 370 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 890 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform -1 0 1170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform 1 0 710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform -1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform 1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform -1 0 1890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 2430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform 1 0 2030 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform -1 0 2250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform -1 0 1150 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform -1 0 850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform 1 0 990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 590 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform -1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform -1 0 510 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform -1 0 270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform -1 0 210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform 1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform 1 0 2130 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform -1 0 2290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform 1 0 1970 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 2370 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 2190 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 1630 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform 1 0 1810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 1710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform 1 0 1550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 1470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform 1 0 1510 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform -1 0 1690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform -1 0 2030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform -1 0 2070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform -1 0 1890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform -1 0 1690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 1170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform -1 0 1350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform -1 0 1030 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform -1 0 570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform -1 0 410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform -1 0 3850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 4050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 4590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform 1 0 5490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform 1 0 6510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform -1 0 5490 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 4770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 4970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform -1 0 4610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform 1 0 5650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform -1 0 5170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform -1 0 5150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 4430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform -1 0 4270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform -1 0 6330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform -1 0 6750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform 1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform 1 0 3510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 6110 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform 1 0 5310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform 1 0 5230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform 1 0 4170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 5030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform 1 0 4810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform 1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform 1 0 5070 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform -1 0 4830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform -1 0 5930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform 1 0 5790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 3830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 3110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 2870 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform -1 0 3050 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 3010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 3510 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 3670 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform -1 0 4010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform 1 0 4330 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform -1 0 5010 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform 1 0 5310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform 1 0 4710 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 5250 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform 1 0 5150 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform -1 0 5370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 5150 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform -1 0 4530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform -1 0 5550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 5130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform -1 0 4790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 4490 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform 1 0 5670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform 1 0 6130 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform 1 0 4250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform -1 0 4310 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform -1 0 3630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform 1 0 3650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform 1 0 3470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 3110 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform 1 0 3370 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform -1 0 3370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform -1 0 2190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 3530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 3350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 3210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform 1 0 2510 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform 1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform 1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform 1 0 2230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 3070 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 2890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform 1 0 4450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 4610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform 1 0 4090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform -1 0 3990 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform 1 0 4670 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 4130 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform -1 0 3830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform -1 0 3130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 3750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform -1 0 3330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 3310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform -1 0 3450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 3570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform -1 0 3670 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform -1 0 3930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 3270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform -1 0 3330 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 3490 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 2770 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 2350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform 1 0 1930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 1850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform -1 0 2190 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform 1 0 2450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform -1 0 2650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 2810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform -1 0 1590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 1790 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform 1 0 1850 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform -1 0 2370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform -1 0 1970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform 1 0 2130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 1270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform -1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 1590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform -1 0 2710 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 2510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 1490 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform -1 0 1430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 1670 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 2010 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 2050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform 1 0 1770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform 1 0 1850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform -1 0 1670 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 2210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 2050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform 1 0 1810 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform -1 0 1430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform -1 0 1350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform 1 0 1950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 2190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform -1 0 2030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 1670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 1990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform -1 0 2210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform 1 0 2170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform -1 0 2350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 2370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform 1 0 1990 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform -1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform -1 0 250 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform 1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform -1 0 750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform 1 0 370 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 890 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform -1 0 710 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 1510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 1190 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 1270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 1290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform 1 0 1870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 1090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform -1 0 1110 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform -1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform -1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform 1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform -1 0 770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 1710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform -1 0 1450 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform -1 0 950 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 1630 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 2110 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform 1 0 1930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform 1 0 2150 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform -1 0 2550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform -1 0 1510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform -1 0 1350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform 1 0 1330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 1310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform -1 0 5210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform 1 0 2910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform 1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform 1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform 1 0 2730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform -1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 5610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 5490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 5770 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform -1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 6350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 6650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 6710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 6710 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform 1 0 4970 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform -1 0 5450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 5290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform 1 0 5490 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform 1 0 5670 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform 1 0 5850 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 5390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 6390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform -1 0 5750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform 1 0 5890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform -1 0 6130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform 1 0 6350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform 1 0 6510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform -1 0 6690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform -1 0 6690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform -1 0 6790 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform 1 0 6450 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform -1 0 6810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 5570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 6530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 6710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 6590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform 1 0 6530 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 5790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform 1 0 6290 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform -1 0 6530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform 1 0 6470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 5470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform 1 0 5690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform -1 0 5870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform 1 0 6030 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 6330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform 1 0 6510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 6170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 5970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 6430 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 6050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform -1 0 6230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform -1 0 6670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform 1 0 6610 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform -1 0 6690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 6790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 6030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform -1 0 6190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 5310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform -1 0 4510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform 1 0 3830 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform 1 0 4170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 5070 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 4650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform 1 0 5770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 5330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 6490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 6810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 6570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 6630 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform 1 0 6130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform -1 0 6330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 5610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform 1 0 4750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform -1 0 4930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform -1 0 5170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform -1 0 4970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform -1 0 4970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 4250 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform -1 0 4470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform -1 0 1870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform -1 0 1330 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform -1 0 1350 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform -1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform 1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform -1 0 4090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 2970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform 1 0 2770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 4310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 4450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform 1 0 5950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 5870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 4410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform 1 0 4710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform 1 0 4550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform 1 0 4850 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform -1 0 4890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform -1 0 5090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 5010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform -1 0 5030 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform 1 0 4290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform -1 0 6050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 5310 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 6190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform -1 0 6530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform -1 0 6230 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform -1 0 6370 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform -1 0 5450 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform -1 0 4370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform -1 0 4750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 4570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform -1 0 4570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform 1 0 3970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform -1 0 4190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform 1 0 550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform 1 0 2330 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform -1 0 4010 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform -1 0 4670 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 4850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform -1 0 4670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 4850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 2350 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform 1 0 4650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform -1 0 2230 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 2310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform 1 0 2370 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform 1 0 2630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform 1 0 2950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform -1 0 2810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform 1 0 2710 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 2170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 1650 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform 1 0 1690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform 1 0 2350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform 1 0 2470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 2850 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform 1 0 4330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 4170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform 1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1452_
timestamp 0
transform 1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1453_
timestamp 0
transform 1 0 2610 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1454_
timestamp 0
transform -1 0 2790 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1455_
timestamp 0
transform -1 0 5230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1456_
timestamp 0
transform 1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1457_
timestamp 0
transform -1 0 5390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1458_
timestamp 0
transform -1 0 5410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1459_
timestamp 0
transform 1 0 3630 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1461_
timestamp 0
transform 1 0 3450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1462_
timestamp 0
transform -1 0 3090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1463_
timestamp 0
transform 1 0 2750 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1464_
timestamp 0
transform 1 0 2190 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 2490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1466_
timestamp 0
transform -1 0 2670 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1467_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1468_
timestamp 0
transform 1 0 3110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1469_
timestamp 0
transform 1 0 2570 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1470_
timestamp 0
transform 1 0 3570 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1471_
timestamp 0
transform -1 0 3810 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1472_
timestamp 0
transform -1 0 3770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1473_
timestamp 0
transform 1 0 4010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1474_
timestamp 0
transform 1 0 5110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1475_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1476_
timestamp 0
transform -1 0 4790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1477_
timestamp 0
transform 1 0 4510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1478_
timestamp 0
transform -1 0 4610 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1479_
timestamp 0
transform -1 0 4370 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1480_
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1482_
timestamp 0
transform -1 0 5590 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1483_
timestamp 0
transform 1 0 3570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 2830 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1485_
timestamp 0
transform 1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1486_
timestamp 0
transform 1 0 3430 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1487_
timestamp 0
transform 1 0 3270 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1488_
timestamp 0
transform 1 0 2950 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 2910 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1490_
timestamp 0
transform -1 0 3250 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 4670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1492_
timestamp 0
transform -1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1493_
timestamp 0
transform -1 0 4010 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1494_
timestamp 0
transform 1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1495_
timestamp 0
transform 1 0 3670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1496_
timestamp 0
transform -1 0 4410 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1497_
timestamp 0
transform 1 0 4930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 4430 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1499_
timestamp 0
transform 1 0 4250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1500_
timestamp 0
transform -1 0 3930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1501_
timestamp 0
transform 1 0 4070 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1502_
timestamp 0
transform 1 0 4170 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1503_
timestamp 0
transform 1 0 4170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1504_
timestamp 0
transform -1 0 4490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1505_
timestamp 0
transform -1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1506_
timestamp 0
transform 1 0 4330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1507_
timestamp 0
transform 1 0 4570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1508_
timestamp 0
transform 1 0 4770 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1509_
timestamp 0
transform 1 0 2170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1510_
timestamp 0
transform -1 0 2570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1511_
timestamp 0
transform 1 0 2350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1512_
timestamp 0
transform 1 0 2470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1513_
timestamp 0
transform -1 0 2550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1514_
timestamp 0
transform -1 0 2550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1515_
timestamp 0
transform 1 0 2650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1516_
timestamp 0
transform -1 0 2830 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1517_
timestamp 0
transform 1 0 3710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1518_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1519_
timestamp 0
transform -1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1520_
timestamp 0
transform 1 0 3150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1521_
timestamp 0
transform -1 0 3970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1522_
timestamp 0
transform -1 0 3830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1523_
timestamp 0
transform 1 0 2970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1524_
timestamp 0
transform -1 0 4030 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1525_
timestamp 0
transform 1 0 3150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1526_
timestamp 0
transform 1 0 3310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 2950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1528_
timestamp 0
transform -1 0 2990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1529_
timestamp 0
transform -1 0 1230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 1370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 1510 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1532_
timestamp 0
transform -1 0 1870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 2030 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1534_
timestamp 0
transform -1 0 2330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 2710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1536_
timestamp 0
transform -1 0 3330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1537_
timestamp 0
transform 1 0 2450 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1538_
timestamp 0
transform 1 0 3850 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1539_
timestamp 0
transform -1 0 3230 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1540_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1541_
timestamp 0
transform -1 0 3410 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1542_
timestamp 0
transform 1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1543_
timestamp 0
transform 1 0 3850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1544_
timestamp 0
transform 1 0 3110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1545_
timestamp 0
transform 1 0 2410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1546_
timestamp 0
transform 1 0 3550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1547_
timestamp 0
transform 1 0 4710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1548_
timestamp 0
transform 1 0 3850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1549_
timestamp 0
transform -1 0 4850 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1550_
timestamp 0
transform 1 0 4970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1551_
timestamp 0
transform -1 0 5170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1552_
timestamp 0
transform 1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1553_
timestamp 0
transform -1 0 4490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1554_
timestamp 0
transform 1 0 5190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1555_
timestamp 0
transform 1 0 4990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1556_
timestamp 0
transform -1 0 5010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1557_
timestamp 0
transform -1 0 4810 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1558_
timestamp 0
transform -1 0 3790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1559_
timestamp 0
transform 1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1560_
timestamp 0
transform -1 0 4970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1561_
timestamp 0
transform -1 0 4610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1562_
timestamp 0
transform 1 0 3930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 4130 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1564_
timestamp 0
transform -1 0 4830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 3510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1566_
timestamp 0
transform 1 0 3450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1567_
timestamp 0
transform -1 0 2970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1568_
timestamp 0
transform 1 0 3610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1569_
timestamp 0
transform -1 0 3270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1570_
timestamp 0
transform 1 0 3090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1571_
timestamp 0
transform 1 0 3150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1572_
timestamp 0
transform 1 0 3330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1573_
timestamp 0
transform 1 0 3890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1574_
timestamp 0
transform -1 0 4430 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1575_
timestamp 0
transform -1 0 3930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1576_
timestamp 0
transform -1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1577_
timestamp 0
transform -1 0 3410 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1578_
timestamp 0
transform -1 0 3770 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1579_
timestamp 0
transform 1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 3650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1581_
timestamp 0
transform -1 0 3850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1582_
timestamp 0
transform 1 0 4290 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 4030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1584_
timestamp 0
transform -1 0 4590 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1585_
timestamp 0
transform 1 0 4190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1586_
timestamp 0
transform -1 0 4670 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1587_
timestamp 0
transform -1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1588_
timestamp 0
transform -1 0 3110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1589_
timestamp 0
transform -1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1590_
timestamp 0
transform -1 0 4270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1591_
timestamp 0
transform 1 0 4230 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1592_
timestamp 0
transform 1 0 4070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1593_
timestamp 0
transform 1 0 2590 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1594_
timestamp 0
transform 1 0 2770 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1595_
timestamp 0
transform -1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1596_
timestamp 0
transform -1 0 3170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1597_
timestamp 0
transform 1 0 2970 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1598_
timestamp 0
transform -1 0 3330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1599_
timestamp 0
transform -1 0 3670 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1600_
timestamp 0
transform 1 0 3470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1601_
timestamp 0
transform -1 0 3410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1602_
timestamp 0
transform -1 0 2870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1603_
timestamp 0
transform -1 0 3050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1604_
timestamp 0
transform -1 0 3230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 4070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1606_
timestamp 0
transform 1 0 6290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1607_
timestamp 0
transform 1 0 6230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1608_
timestamp 0
transform -1 0 6410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1609_
timestamp 0
transform 1 0 6170 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1610_
timestamp 0
transform 1 0 6570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1611_
timestamp 0
transform 1 0 5610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1612_
timestamp 0
transform -1 0 6830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1613_
timestamp 0
transform -1 0 6450 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1614_
timestamp 0
transform -1 0 6270 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1615_
timestamp 0
transform -1 0 6090 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1616_
timestamp 0
transform 1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1617_
timestamp 0
transform 1 0 5630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1618_
timestamp 0
transform -1 0 5430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1619_
timestamp 0
transform 1 0 5330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1620_
timestamp 0
transform -1 0 6110 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1621_
timestamp 0
transform 1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1622_
timestamp 0
transform 1 0 6750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1623_
timestamp 0
transform 1 0 6410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1624_
timestamp 0
transform -1 0 6810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1625_
timestamp 0
transform -1 0 6550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1626_
timestamp 0
transform 1 0 6530 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1627_
timestamp 0
transform 1 0 6370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1628_
timestamp 0
transform -1 0 6170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1629_
timestamp 0
transform 1 0 5950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1630_
timestamp 0
transform 1 0 6670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1631_
timestamp 0
transform -1 0 6730 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1632_
timestamp 0
transform -1 0 6610 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1633_
timestamp 0
transform -1 0 6630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1634_
timestamp 0
transform -1 0 6450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1635_
timestamp 0
transform 1 0 6250 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1636_
timestamp 0
transform -1 0 6430 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1637_
timestamp 0
transform 1 0 6070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1638_
timestamp 0
transform -1 0 6470 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1639_
timestamp 0
transform 1 0 6330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 5670 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1641_
timestamp 0
transform -1 0 6730 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1642_
timestamp 0
transform -1 0 6230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1643_
timestamp 0
transform -1 0 6530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1644_
timestamp 0
transform -1 0 6230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1645_
timestamp 0
transform 1 0 6550 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1646_
timestamp 0
transform -1 0 6690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1647_
timestamp 0
transform -1 0 6010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1648_
timestamp 0
transform 1 0 5790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1649_
timestamp 0
transform -1 0 6690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1650_
timestamp 0
transform -1 0 6690 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1651_
timestamp 0
transform -1 0 6250 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1652_
timestamp 0
transform -1 0 6470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1653_
timestamp 0
transform 1 0 5590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1654_
timestamp 0
transform 1 0 6370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1655_
timestamp 0
transform 1 0 6350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1656_
timestamp 0
transform 1 0 6530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1657_
timestamp 0
transform -1 0 6790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1658_
timestamp 0
transform 1 0 6130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1659_
timestamp 0
transform -1 0 6830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1660_
timestamp 0
transform -1 0 6610 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1661_
timestamp 0
transform -1 0 6790 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1662_
timestamp 0
transform -1 0 6430 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1663_
timestamp 0
transform 1 0 6010 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1664_
timestamp 0
transform 1 0 6190 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1665_
timestamp 0
transform -1 0 6310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1666_
timestamp 0
transform -1 0 6630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1667_
timestamp 0
transform 1 0 6390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1668_
timestamp 0
transform 1 0 6690 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1669_
timestamp 0
transform -1 0 5970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1670_
timestamp 0
transform 1 0 5830 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1671_
timestamp 0
transform 1 0 5510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1672_
timestamp 0
transform -1 0 6070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1673_
timestamp 0
transform 1 0 5690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1674_
timestamp 0
transform -1 0 5890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1675_
timestamp 0
transform 1 0 3990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1676_
timestamp 0
transform 1 0 5170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1677_
timestamp 0
transform 1 0 5090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1711_
timestamp 0
transform -1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1712_
timestamp 0
transform -1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 1050 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1714_
timestamp 0
transform 1 0 190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1715_
timestamp 0
transform -1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1716_
timestamp 0
transform -1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1717_
timestamp 0
transform 1 0 350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1718_
timestamp 0
transform -1 0 50 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1719_
timestamp 0
transform 1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1721_
timestamp 0
transform -1 0 210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1722_
timestamp 0
transform -1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 1490 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1724_
timestamp 0
transform 1 0 350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_1__1725_
timestamp 0
transform -1 0 410 0 1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform -1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 230 0 1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 5790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform -1 0 5370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 5610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform -1 0 2470 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 3330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert4
timestamp 0
transform 1 0 4950 0 1 790
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert5
timestamp 0
transform -1 0 1910 0 1 4950
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert6
timestamp 0
transform -1 0 4770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert7
timestamp 0
transform 1 0 490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert8
timestamp 0
transform -1 0 390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert9
timestamp 0
transform 1 0 2570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert10
timestamp 0
transform -1 0 3550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__828_
timestamp 0
transform 1 0 830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__829_
timestamp 0
transform 1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__830_
timestamp 0
transform -1 0 2370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__831_
timestamp 0
transform -1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__832_
timestamp 0
transform 1 0 2270 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__833_
timestamp 0
transform 1 0 1970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__834_
timestamp 0
transform -1 0 1590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__835_
timestamp 0
transform -1 0 1670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__836_
timestamp 0
transform -1 0 990 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__837_
timestamp 0
transform 1 0 870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__838_
timestamp 0
transform -1 0 710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__839_
timestamp 0
transform -1 0 910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__840_
timestamp 0
transform 1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__841_
timestamp 0
transform -1 0 70 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__842_
timestamp 0
transform 1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__843_
timestamp 0
transform -1 0 230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__844_
timestamp 0
transform 1 0 690 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__845_
timestamp 0
transform 1 0 230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__846_
timestamp 0
transform -1 0 750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__847_
timestamp 0
transform -1 0 910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__848_
timestamp 0
transform -1 0 570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__849_
timestamp 0
transform 1 0 210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__850_
timestamp 0
transform -1 0 230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__851_
timestamp 0
transform -1 0 870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__852_
timestamp 0
transform -1 0 690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__853_
timestamp 0
transform 1 0 570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__854_
timestamp 0
transform -1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__855_
timestamp 0
transform -1 0 550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__856_
timestamp 0
transform -1 0 750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__857_
timestamp 0
transform 1 0 1010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__858_
timestamp 0
transform -1 0 490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__859_
timestamp 0
transform 1 0 50 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__860_
timestamp 0
transform 1 0 1070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__861_
timestamp 0
transform 1 0 830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__862_
timestamp 0
transform -1 0 710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__863_
timestamp 0
transform -1 0 530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__864_
timestamp 0
transform 1 0 830 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__865_
timestamp 0
transform 1 0 410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__866_
timestamp 0
transform -1 0 1370 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__867_
timestamp 0
transform 1 0 990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__868_
timestamp 0
transform 1 0 1010 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__869_
timestamp 0
transform -1 0 1210 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__870_
timestamp 0
transform 1 0 1130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__871_
timestamp 0
transform -1 0 1430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__872_
timestamp 0
transform -1 0 870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__873_
timestamp 0
transform 1 0 1030 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__874_
timestamp 0
transform 1 0 1010 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__875_
timestamp 0
transform 1 0 1250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__876_
timestamp 0
transform -1 0 1170 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__877_
timestamp 0
transform 1 0 1310 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__878_
timestamp 0
transform -1 0 850 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__879_
timestamp 0
transform -1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__880_
timestamp 0
transform 1 0 1170 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__881_
timestamp 0
transform 1 0 210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__882_
timestamp 0
transform -1 0 210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__883_
timestamp 0
transform 1 0 850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__884_
timestamp 0
transform -1 0 1010 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__885_
timestamp 0
transform -1 0 1030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__886_
timestamp 0
transform -1 0 850 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__887_
timestamp 0
transform 1 0 850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__888_
timestamp 0
transform -1 0 670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__889_
timestamp 0
transform 1 0 510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__890_
timestamp 0
transform -1 0 690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__891_
timestamp 0
transform 1 0 330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__892_
timestamp 0
transform -1 0 510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__893_
timestamp 0
transform -1 0 210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__894_
timestamp 0
transform -1 0 530 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__895_
timestamp 0
transform -1 0 690 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__896_
timestamp 0
transform 1 0 1810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__897_
timestamp 0
transform -1 0 2530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__898_
timestamp 0
transform -1 0 2190 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__899_
timestamp 0
transform 1 0 2130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__900_
timestamp 0
transform -1 0 1750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__901_
timestamp 0
transform 1 0 1630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__902_
timestamp 0
transform -1 0 1670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__903_
timestamp 0
transform -1 0 1810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__904_
timestamp 0
transform -1 0 1490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__905_
timestamp 0
transform -1 0 1410 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__906_
timestamp 0
transform 1 0 1210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__907_
timestamp 0
transform 1 0 1790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__908_
timestamp 0
transform 1 0 2290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__909_
timestamp 0
transform 1 0 2010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__910_
timestamp 0
transform -1 0 1850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__911_
timestamp 0
transform 1 0 1610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__912_
timestamp 0
transform -1 0 1750 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__913_
timestamp 0
transform 1 0 2850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__914_
timestamp 0
transform -1 0 3190 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__915_
timestamp 0
transform 1 0 2110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__916_
timestamp 0
transform -1 0 2110 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__917_
timestamp 0
transform 1 0 1550 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__918_
timestamp 0
transform 1 0 1950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__919_
timestamp 0
transform -1 0 3010 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__920_
timestamp 0
transform -1 0 3270 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__921_
timestamp 0
transform 1 0 2650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform -1 0 2490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform -1 0 2310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform 1 0 1910 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform 1 0 2590 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform -1 0 2750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform -1 0 3410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform -1 0 3090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform -1 0 2570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform -1 0 2390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform -1 0 930 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform -1 0 2910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform -1 0 2850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform -1 0 2430 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform -1 0 750 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform -1 0 1190 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform -1 0 690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform 1 0 1830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform -1 0 1230 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 1690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform 1 0 1490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform 1 0 990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform -1 0 390 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform -1 0 1170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform 1 0 2050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform 1 0 1530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform 1 0 1710 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform 1 0 1550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform -1 0 3010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform -1 0 6070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform -1 0 6390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform 1 0 5890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform -1 0 5730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform 1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform 1 0 3230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform 1 0 2910 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform -1 0 6510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform 1 0 5750 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform 1 0 5590 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform -1 0 5430 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform 1 0 5250 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform 1 0 3490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform -1 0 3510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform -1 0 5310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform 1 0 3890 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform -1 0 4110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform -1 0 3250 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform -1 0 3950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform 1 0 3630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform -1 0 4470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform 1 0 2890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform -1 0 6350 0 1 790
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform -1 0 6230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform 1 0 5990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform 1 0 6170 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform 1 0 4210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform 1 0 4270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform -1 0 4250 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform 1 0 5550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform 1 0 6050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform -1 0 6810 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform -1 0 5990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform -1 0 5830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform -1 0 5670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform -1 0 4770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform 1 0 5990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform -1 0 5550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform -1 0 5470 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform -1 0 5770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform -1 0 5610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 5130 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform 1 0 4930 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform 1 0 4690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 4850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform -1 0 5330 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform -1 0 5510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform 1 0 5370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform -1 0 4790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform -1 0 4630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform -1 0 5270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform -1 0 5170 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform -1 0 3890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform 1 0 3710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform -1 0 2990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform -1 0 2670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform -1 0 4070 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform 1 0 3650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 2910 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform 1 0 6270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform 1 0 4850 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform 1 0 3770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform -1 0 6890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform 1 0 4570 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform 1 0 4070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform 1 0 3870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform -1 0 4430 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform -1 0 4250 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform 1 0 6390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform 1 0 3930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform -1 0 4530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform -1 0 4690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform 1 0 4010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform -1 0 4190 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 4350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform 1 0 3710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform -1 0 4410 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform -1 0 2610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform 1 0 4210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform -1 0 4050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform -1 0 3790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform 1 0 3290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform -1 0 3490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform -1 0 4590 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform -1 0 4070 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform 1 0 3710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform -1 0 3850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform -1 0 3910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform 1 0 3710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform -1 0 3550 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform -1 0 3070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform 1 0 3390 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform -1 0 3570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform -1 0 3430 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform 1 0 530 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform 1 0 690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform 1 0 1090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform 1 0 790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform -1 0 950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform -1 0 1050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform -1 0 890 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform -1 0 1330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform 1 0 2410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform -1 0 3250 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform -1 0 3070 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform -1 0 2750 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform 1 0 1490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform -1 0 1390 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform 1 0 1210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform -1 0 3170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform -1 0 2830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform -1 0 2690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 1870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform -1 0 2350 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform 1 0 1490 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform -1 0 1530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform 1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform -1 0 1530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform -1 0 1210 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform 1 0 1330 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform -1 0 950 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform 1 0 410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform 1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform -1 0 390 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform 1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 910 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform -1 0 1190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform 1 0 730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform -1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform 1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform -1 0 1910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 2450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform 1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform -1 0 2270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform -1 0 1170 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform -1 0 770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform -1 0 870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform 1 0 1010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform -1 0 610 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform -1 0 710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform -1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform -1 0 530 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform 1 0 530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform -1 0 290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform -1 0 230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform 1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform 1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform 1 0 230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform 1 0 2150 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform -1 0 2310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform 1 0 1990 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform -1 0 2390 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform 1 0 2210 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform 1 0 1650 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform 1 0 1830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform 1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform 1 0 1570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform 1 0 1490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform 1 0 1530 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform -1 0 1710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform -1 0 2050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform -1 0 2090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform -1 0 1910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 1190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform -1 0 1370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform -1 0 1050 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform -1 0 590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform -1 0 430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform -1 0 3870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 4070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform -1 0 4610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform 1 0 5510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform 1 0 6530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform -1 0 5510 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 4790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform -1 0 4990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform -1 0 4630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform 1 0 5670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform -1 0 5190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform -1 0 5170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform -1 0 4450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform -1 0 4290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform -1 0 6350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform -1 0 6770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform 1 0 3210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform 1 0 3530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform -1 0 6130 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform 1 0 5330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform 1 0 5250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform 1 0 4190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform -1 0 5050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform 1 0 4830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform 1 0 5070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform 1 0 5090 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform -1 0 4850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform -1 0 5950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform 1 0 5810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform 1 0 3850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform 1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform 1 0 2890 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform -1 0 3070 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform 1 0 3030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 3530 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform 1 0 3690 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform -1 0 4030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform 1 0 4350 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform -1 0 5030 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform 1 0 5330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform 1 0 4730 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform 1 0 5270 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform 1 0 5170 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform -1 0 5390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform 1 0 5170 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform -1 0 4550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform -1 0 5570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 5150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform -1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform -1 0 4510 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform 1 0 5690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform 1 0 6150 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform 1 0 4270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform -1 0 4330 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform -1 0 3650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform 1 0 3670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform 1 0 3490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform 1 0 3130 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform 1 0 3390 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform -1 0 3390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform -1 0 2210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform 1 0 3550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 3370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform -1 0 3230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform 1 0 2530 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform 1 0 2430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform 1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform 1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform 1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform -1 0 3090 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform 1 0 2710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform 1 0 4470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 4630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform 1 0 4110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform -1 0 4010 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform 1 0 4690 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform 1 0 4150 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform -1 0 3850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform -1 0 3150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform 1 0 3770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform -1 0 3350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform 1 0 3330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform -1 0 3470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform 1 0 3590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform -1 0 3690 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform -1 0 3950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform 1 0 3290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform -1 0 3350 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform -1 0 3510 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 2790 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform 1 0 2370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform 1 0 1950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform -1 0 1870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform -1 0 2210 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform 1 0 2470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform -1 0 2670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform 1 0 2830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform -1 0 1610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 1810 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform 1 0 1870 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform -1 0 2390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform -1 0 1990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform 1 0 2150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 1290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform -1 0 1650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 1610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform -1 0 2730 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 2530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform -1 0 1510 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform -1 0 1450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform 1 0 1690 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform -1 0 2030 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform -1 0 2070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform 1 0 1790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform 1 0 1870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform -1 0 1690 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform 1 0 2230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 2070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform 1 0 1830 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform -1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform -1 0 1370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform 1 0 1970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform -1 0 2210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform -1 0 2050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform -1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform 1 0 1690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform 1 0 2010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform -1 0 2230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform 1 0 2190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform -1 0 2370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 2390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform 1 0 2010 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform -1 0 2610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform -1 0 270 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform -1 0 430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform 1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 390 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform -1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform 1 0 390 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform -1 0 910 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform -1 0 730 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform 1 0 570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform 1 0 1530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 1210 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform -1 0 1290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform -1 0 1310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform 1 0 1890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform -1 0 1110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform -1 0 1130 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform -1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform -1 0 70 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform -1 0 230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform 1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform -1 0 790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform 1 0 1730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform -1 0 1470 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform -1 0 970 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform -1 0 1650 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform 1 0 2130 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform 1 0 1950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform 1 0 2170 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform -1 0 2570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform -1 0 1530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform -1 0 1370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform 1 0 1350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform 1 0 1330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform -1 0 5230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform 1 0 2930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform 1 0 2570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform 1 0 1650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform 1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform 1 0 2750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform -1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 5630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform 1 0 5510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 5790 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform -1 0 5690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform -1 0 6370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform -1 0 6670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform -1 0 6730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 6730 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform 1 0 4990 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform -1 0 5470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 5310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform 1 0 5510 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform 1 0 5690 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform 1 0 5870 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 5410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform 1 0 6410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform -1 0 5770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform 1 0 5910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform -1 0 6150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform 1 0 6370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform 1 0 6530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform -1 0 6710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform -1 0 6710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform -1 0 6810 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform 1 0 6470 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform -1 0 6830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 5590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform 1 0 6550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 6730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform 1 0 6610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform 1 0 6550 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 5810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform 1 0 6310 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform -1 0 6550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform 1 0 6490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform 1 0 5490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform 1 0 5710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform -1 0 5890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform 1 0 6050 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform 1 0 6350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform 1 0 6530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 6190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform 1 0 5990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform 1 0 6450 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform 1 0 6070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform -1 0 6250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform -1 0 6690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform 1 0 6630 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform -1 0 6710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform -1 0 6810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform -1 0 6050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform -1 0 6210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform -1 0 5330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform -1 0 4530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform 1 0 3850 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform 1 0 4190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform -1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform -1 0 4670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform 1 0 5790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform -1 0 5350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform 1 0 6510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform -1 0 6830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform -1 0 6590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform -1 0 6650 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform 1 0 6150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform -1 0 6350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform -1 0 5630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform 1 0 4770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform -1 0 4950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform -1 0 5190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform -1 0 4990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform -1 0 4990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 4270 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform -1 0 4490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform -1 0 1350 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform -1 0 1370 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform -1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform 1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform -1 0 4110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform -1 0 2990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform 1 0 2790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform 1 0 4330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform 1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform 1 0 5970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform -1 0 5890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 4430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform 1 0 4730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform 1 0 4570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform 1 0 4870 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform -1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform -1 0 5110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 5030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform -1 0 5050 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform 1 0 4310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform -1 0 6070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 5330 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform 1 0 6210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform -1 0 6550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform -1 0 6250 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform -1 0 6390 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform -1 0 5470 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform -1 0 5010 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform -1 0 4390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform -1 0 4770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform -1 0 4590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 4370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform -1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform 1 0 3990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform -1 0 4210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform 1 0 750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform 1 0 570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform 1 0 2350 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform -1 0 4030 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform -1 0 4690 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform -1 0 4870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform -1 0 4690 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 4870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform 1 0 2370 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform 1 0 4670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform -1 0 2250 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform 1 0 2330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform 1 0 2390 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform 1 0 2650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform 1 0 2970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform -1 0 2830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform 1 0 2730 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform 1 0 2190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform 1 0 1670 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform 1 0 1710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform 1 0 2370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform 1 0 2490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform 1 0 4350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform -1 0 4190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform 1 0 4810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1452_
timestamp 0
transform 1 0 2810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1453_
timestamp 0
transform 1 0 2630 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1454_
timestamp 0
transform -1 0 2810 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1455_
timestamp 0
transform -1 0 5250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1456_
timestamp 0
transform 1 0 5250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1457_
timestamp 0
transform -1 0 5410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1458_
timestamp 0
transform -1 0 5430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1459_
timestamp 0
transform 1 0 3650 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1460_
timestamp 0
transform 1 0 4410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1461_
timestamp 0
transform 1 0 3470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1462_
timestamp 0
transform -1 0 3110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1463_
timestamp 0
transform 1 0 2770 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1464_
timestamp 0
transform 1 0 2210 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1465_
timestamp 0
transform 1 0 2510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1466_
timestamp 0
transform -1 0 2690 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1467_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1468_
timestamp 0
transform 1 0 3130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1469_
timestamp 0
transform 1 0 2590 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1470_
timestamp 0
transform 1 0 3590 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1471_
timestamp 0
transform -1 0 3830 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1472_
timestamp 0
transform -1 0 3790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1473_
timestamp 0
transform 1 0 4030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1474_
timestamp 0
transform 1 0 5130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1475_
timestamp 0
transform -1 0 4230 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1476_
timestamp 0
transform -1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1477_
timestamp 0
transform 1 0 4530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1478_
timestamp 0
transform -1 0 4630 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1479_
timestamp 0
transform -1 0 4390 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1480_
timestamp 0
transform 1 0 5970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1481_
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1482_
timestamp 0
transform -1 0 5610 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1483_
timestamp 0
transform 1 0 3590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1484_
timestamp 0
transform -1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1485_
timestamp 0
transform 1 0 3010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1486_
timestamp 0
transform 1 0 3450 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1487_
timestamp 0
transform 1 0 3290 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1488_
timestamp 0
transform 1 0 2970 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1489_
timestamp 0
transform 1 0 2930 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1490_
timestamp 0
transform -1 0 3270 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1491_
timestamp 0
transform -1 0 4690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1492_
timestamp 0
transform -1 0 4590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1493_
timestamp 0
transform -1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1494_
timestamp 0
transform 1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1495_
timestamp 0
transform 1 0 3690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1496_
timestamp 0
transform -1 0 4430 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1497_
timestamp 0
transform 1 0 4950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1498_
timestamp 0
transform 1 0 4450 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1499_
timestamp 0
transform 1 0 4270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1500_
timestamp 0
transform -1 0 3950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1501_
timestamp 0
transform 1 0 4090 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1502_
timestamp 0
transform 1 0 4190 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1503_
timestamp 0
transform 1 0 4190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1504_
timestamp 0
transform -1 0 4510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1505_
timestamp 0
transform -1 0 4150 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1506_
timestamp 0
transform 1 0 4350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1507_
timestamp 0
transform 1 0 4590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1508_
timestamp 0
transform 1 0 4790 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1509_
timestamp 0
transform 1 0 2190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1510_
timestamp 0
transform -1 0 2590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1511_
timestamp 0
transform 1 0 2370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1512_
timestamp 0
transform 1 0 2490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1513_
timestamp 0
transform -1 0 2570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1514_
timestamp 0
transform -1 0 2570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1515_
timestamp 0
transform 1 0 2670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1516_
timestamp 0
transform -1 0 2850 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1517_
timestamp 0
transform 1 0 3730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1518_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1519_
timestamp 0
transform -1 0 4190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1520_
timestamp 0
transform 1 0 3170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1521_
timestamp 0
transform -1 0 3990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1522_
timestamp 0
transform -1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1523_
timestamp 0
transform 1 0 2990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1524_
timestamp 0
transform -1 0 4050 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1525_
timestamp 0
transform 1 0 3170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1526_
timestamp 0
transform 1 0 3330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1527_
timestamp 0
transform 1 0 2970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1528_
timestamp 0
transform -1 0 3010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1529_
timestamp 0
transform -1 0 1250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 1390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1531_
timestamp 0
transform 1 0 1530 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1532_
timestamp 0
transform -1 0 1890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1533_
timestamp 0
transform -1 0 2050 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1534_
timestamp 0
transform -1 0 2350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1535_
timestamp 0
transform -1 0 2730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1536_
timestamp 0
transform -1 0 3350 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1537_
timestamp 0
transform 1 0 2470 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1538_
timestamp 0
transform 1 0 3870 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1539_
timestamp 0
transform -1 0 3250 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1540_
timestamp 0
transform 1 0 1810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1541_
timestamp 0
transform -1 0 3430 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1542_
timestamp 0
transform 1 0 2010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1543_
timestamp 0
transform 1 0 3870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1544_
timestamp 0
transform 1 0 3130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1545_
timestamp 0
transform 1 0 2430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1546_
timestamp 0
transform 1 0 3570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1547_
timestamp 0
transform 1 0 4730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1548_
timestamp 0
transform 1 0 3870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1549_
timestamp 0
transform -1 0 4870 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1550_
timestamp 0
transform 1 0 4990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1551_
timestamp 0
transform -1 0 5190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1552_
timestamp 0
transform 1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1553_
timestamp 0
transform -1 0 4510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1554_
timestamp 0
transform 1 0 5210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1555_
timestamp 0
transform 1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1556_
timestamp 0
transform -1 0 5030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1557_
timestamp 0
transform -1 0 4830 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1558_
timestamp 0
transform -1 0 3810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1559_
timestamp 0
transform 1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1560_
timestamp 0
transform -1 0 4990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1561_
timestamp 0
transform -1 0 4630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1562_
timestamp 0
transform 1 0 3950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1563_
timestamp 0
transform -1 0 4150 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1564_
timestamp 0
transform -1 0 4850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1565_
timestamp 0
transform 1 0 3530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1566_
timestamp 0
transform 1 0 3470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1567_
timestamp 0
transform -1 0 2990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1568_
timestamp 0
transform 1 0 3630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1569_
timestamp 0
transform -1 0 3290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1570_
timestamp 0
transform 1 0 3110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1571_
timestamp 0
transform 1 0 3170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1572_
timestamp 0
transform 1 0 3350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1573_
timestamp 0
transform 1 0 3910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1574_
timestamp 0
transform -1 0 4450 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1575_
timestamp 0
transform -1 0 3950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1576_
timestamp 0
transform -1 0 4110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1577_
timestamp 0
transform -1 0 3430 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1578_
timestamp 0
transform -1 0 3790 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1579_
timestamp 0
transform 1 0 3590 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1580_
timestamp 0
transform 1 0 3670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1581_
timestamp 0
transform -1 0 3870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1582_
timestamp 0
transform 1 0 4310 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1583_
timestamp 0
transform -1 0 4050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1584_
timestamp 0
transform -1 0 4610 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1585_
timestamp 0
transform 1 0 4210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1586_
timestamp 0
transform -1 0 4690 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1587_
timestamp 0
transform -1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1588_
timestamp 0
transform -1 0 3130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1589_
timestamp 0
transform -1 0 4430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1590_
timestamp 0
transform -1 0 4290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1591_
timestamp 0
transform 1 0 4250 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1592_
timestamp 0
transform 1 0 4090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1593_
timestamp 0
transform 1 0 2610 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1594_
timestamp 0
transform 1 0 2790 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1595_
timestamp 0
transform -1 0 2990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1596_
timestamp 0
transform -1 0 3190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1597_
timestamp 0
transform 1 0 2990 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1598_
timestamp 0
transform -1 0 3350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1599_
timestamp 0
transform -1 0 3690 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1600_
timestamp 0
transform 1 0 3490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1601_
timestamp 0
transform -1 0 3430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1602_
timestamp 0
transform -1 0 2890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1603_
timestamp 0
transform -1 0 3070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1604_
timestamp 0
transform -1 0 3250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1605_
timestamp 0
transform 1 0 4090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1606_
timestamp 0
transform 1 0 6310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1607_
timestamp 0
transform 1 0 6250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1608_
timestamp 0
transform -1 0 6430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1609_
timestamp 0
transform 1 0 6190 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1610_
timestamp 0
transform 1 0 6590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1611_
timestamp 0
transform 1 0 5630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1612_
timestamp 0
transform -1 0 6850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1613_
timestamp 0
transform -1 0 6470 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1614_
timestamp 0
transform -1 0 6290 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1615_
timestamp 0
transform -1 0 6110 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1616_
timestamp 0
transform 1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1617_
timestamp 0
transform 1 0 5650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1618_
timestamp 0
transform -1 0 5450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1619_
timestamp 0
transform 1 0 5350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1620_
timestamp 0
transform -1 0 6130 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1621_
timestamp 0
transform 1 0 5350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1622_
timestamp 0
transform 1 0 6770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1623_
timestamp 0
transform 1 0 6430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1624_
timestamp 0
transform -1 0 6830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1625_
timestamp 0
transform -1 0 6570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1626_
timestamp 0
transform 1 0 6550 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1627_
timestamp 0
transform 1 0 6390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1628_
timestamp 0
transform -1 0 6190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1629_
timestamp 0
transform 1 0 5970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1630_
timestamp 0
transform 1 0 6690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1631_
timestamp 0
transform -1 0 6750 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1632_
timestamp 0
transform -1 0 6630 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1633_
timestamp 0
transform -1 0 6650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1634_
timestamp 0
transform -1 0 6470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1635_
timestamp 0
transform 1 0 6270 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1636_
timestamp 0
transform -1 0 6450 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1637_
timestamp 0
transform 1 0 6090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1638_
timestamp 0
transform -1 0 6490 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1639_
timestamp 0
transform 1 0 6350 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1640_
timestamp 0
transform 1 0 5690 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1641_
timestamp 0
transform -1 0 6750 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1642_
timestamp 0
transform -1 0 6250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1643_
timestamp 0
transform -1 0 6550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1644_
timestamp 0
transform -1 0 6250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1645_
timestamp 0
transform 1 0 6570 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1646_
timestamp 0
transform -1 0 6710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1647_
timestamp 0
transform -1 0 6030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1648_
timestamp 0
transform 1 0 5810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1649_
timestamp 0
transform -1 0 6710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1650_
timestamp 0
transform -1 0 6710 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1651_
timestamp 0
transform -1 0 6270 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1652_
timestamp 0
transform -1 0 6490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1653_
timestamp 0
transform 1 0 5610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1654_
timestamp 0
transform 1 0 6390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1655_
timestamp 0
transform 1 0 6370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1656_
timestamp 0
transform 1 0 6550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1657_
timestamp 0
transform -1 0 6810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1658_
timestamp 0
transform 1 0 6150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1659_
timestamp 0
transform -1 0 6850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1660_
timestamp 0
transform -1 0 6630 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1661_
timestamp 0
transform -1 0 6810 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1662_
timestamp 0
transform -1 0 6450 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1663_
timestamp 0
transform 1 0 6030 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1664_
timestamp 0
transform 1 0 6210 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1665_
timestamp 0
transform -1 0 6330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1666_
timestamp 0
transform -1 0 6650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1667_
timestamp 0
transform 1 0 6410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1668_
timestamp 0
transform 1 0 6710 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1669_
timestamp 0
transform -1 0 5990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1670_
timestamp 0
transform 1 0 5850 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1671_
timestamp 0
transform 1 0 5530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1672_
timestamp 0
transform -1 0 6090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1673_
timestamp 0
transform 1 0 5710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1674_
timestamp 0
transform -1 0 5910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1675_
timestamp 0
transform 1 0 4010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1676_
timestamp 0
transform 1 0 5190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1677_
timestamp 0
transform 1 0 5110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1711_
timestamp 0
transform -1 0 70 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1712_
timestamp 0
transform -1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1713_
timestamp 0
transform -1 0 1070 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1714_
timestamp 0
transform 1 0 210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1715_
timestamp 0
transform -1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1716_
timestamp 0
transform -1 0 70 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1717_
timestamp 0
transform 1 0 370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1718_
timestamp 0
transform -1 0 70 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1719_
timestamp 0
transform 1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1720_
timestamp 0
transform -1 0 70 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1721_
timestamp 0
transform -1 0 230 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1722_
timestamp 0
transform -1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1723_
timestamp 0
transform 1 0 1510 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1724_
timestamp 0
transform 1 0 370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_2__1725_
timestamp 0
transform -1 0 430 0 1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform -1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 250 0 1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform 1 0 210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform 1 0 370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform 1 0 5810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform -1 0 5390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 5630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform -1 0 2490 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 3350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert4
timestamp 0
transform 1 0 4970 0 1 790
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert5
timestamp 0
transform -1 0 1930 0 1 4950
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert6
timestamp 0
transform -1 0 4790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert7
timestamp 0
transform 1 0 510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert8
timestamp 0
transform -1 0 410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert9
timestamp 0
transform 1 0 2590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert10
timestamp 0
transform -1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__828_
timestamp 0
transform 1 0 850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__829_
timestamp 0
transform 1 0 1530 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__830_
timestamp 0
transform -1 0 2390 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__831_
timestamp 0
transform -1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__832_
timestamp 0
transform 1 0 2290 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__833_
timestamp 0
transform 1 0 1990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__834_
timestamp 0
transform -1 0 1610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__835_
timestamp 0
transform -1 0 1690 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__836_
timestamp 0
transform -1 0 1010 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__837_
timestamp 0
transform 1 0 890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__838_
timestamp 0
transform -1 0 730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__839_
timestamp 0
transform -1 0 930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__840_
timestamp 0
transform 1 0 70 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__841_
timestamp 0
transform -1 0 90 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__842_
timestamp 0
transform 1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__843_
timestamp 0
transform -1 0 250 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__844_
timestamp 0
transform 1 0 710 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__845_
timestamp 0
transform 1 0 250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__846_
timestamp 0
transform -1 0 770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__847_
timestamp 0
transform -1 0 930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__848_
timestamp 0
transform -1 0 590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__849_
timestamp 0
transform 1 0 230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__850_
timestamp 0
transform -1 0 250 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__851_
timestamp 0
transform -1 0 890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__852_
timestamp 0
transform -1 0 710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__853_
timestamp 0
transform 1 0 590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__854_
timestamp 0
transform -1 0 90 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__855_
timestamp 0
transform -1 0 570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__856_
timestamp 0
transform -1 0 770 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__857_
timestamp 0
transform 1 0 1030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__858_
timestamp 0
transform -1 0 510 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__859_
timestamp 0
transform 1 0 70 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__860_
timestamp 0
transform 1 0 1090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__861_
timestamp 0
transform 1 0 850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__862_
timestamp 0
transform -1 0 730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__863_
timestamp 0
transform -1 0 550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__864_
timestamp 0
transform 1 0 850 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__865_
timestamp 0
transform 1 0 430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__866_
timestamp 0
transform -1 0 1390 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__867_
timestamp 0
transform 1 0 1010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__868_
timestamp 0
transform 1 0 1030 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__869_
timestamp 0
transform -1 0 1230 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__870_
timestamp 0
transform 1 0 1150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__871_
timestamp 0
transform -1 0 1450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__872_
timestamp 0
transform -1 0 890 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__873_
timestamp 0
transform 1 0 1050 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__874_
timestamp 0
transform 1 0 1030 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__875_
timestamp 0
transform 1 0 1270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__876_
timestamp 0
transform -1 0 1190 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__877_
timestamp 0
transform 1 0 1330 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__878_
timestamp 0
transform -1 0 870 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__879_
timestamp 0
transform -1 0 90 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__880_
timestamp 0
transform 1 0 1190 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__881_
timestamp 0
transform 1 0 230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__882_
timestamp 0
transform -1 0 230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__883_
timestamp 0
transform 1 0 870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__884_
timestamp 0
transform -1 0 1030 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__885_
timestamp 0
transform -1 0 1050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__886_
timestamp 0
transform -1 0 870 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__887_
timestamp 0
transform 1 0 870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__888_
timestamp 0
transform -1 0 690 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__889_
timestamp 0
transform 1 0 530 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__890_
timestamp 0
transform -1 0 710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__891_
timestamp 0
transform 1 0 350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__892_
timestamp 0
transform -1 0 530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__893_
timestamp 0
transform -1 0 230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__894_
timestamp 0
transform -1 0 550 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__895_
timestamp 0
transform -1 0 710 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__896_
timestamp 0
transform 1 0 1830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__897_
timestamp 0
transform -1 0 2550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__898_
timestamp 0
transform -1 0 2210 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__899_
timestamp 0
transform 1 0 2150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__900_
timestamp 0
transform -1 0 1770 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__901_
timestamp 0
transform 1 0 1650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__902_
timestamp 0
transform -1 0 1690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__903_
timestamp 0
transform -1 0 1830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__904_
timestamp 0
transform -1 0 1510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__905_
timestamp 0
transform -1 0 1430 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__906_
timestamp 0
transform 1 0 1230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__907_
timestamp 0
transform 1 0 1810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__908_
timestamp 0
transform 1 0 2310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__909_
timestamp 0
transform 1 0 2030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__910_
timestamp 0
transform -1 0 1870 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__911_
timestamp 0
transform 1 0 1630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__912_
timestamp 0
transform -1 0 1770 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__913_
timestamp 0
transform 1 0 2870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__914_
timestamp 0
transform -1 0 3210 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__915_
timestamp 0
transform 1 0 2130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__916_
timestamp 0
transform -1 0 2130 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__917_
timestamp 0
transform 1 0 1570 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__918_
timestamp 0
transform 1 0 1970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__919_
timestamp 0
transform -1 0 3030 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__920_
timestamp 0
transform -1 0 3290 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__921_
timestamp 0
transform 1 0 2670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__922_
timestamp 0
transform -1 0 2510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__923_
timestamp 0
transform -1 0 2330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__924_
timestamp 0
transform 1 0 1930 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__925_
timestamp 0
transform 1 0 2610 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__926_
timestamp 0
transform -1 0 2770 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__927_
timestamp 0
transform -1 0 3430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__928_
timestamp 0
transform -1 0 3110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__929_
timestamp 0
transform -1 0 2590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__930_
timestamp 0
transform -1 0 2410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform -1 0 950 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__932_
timestamp 0
transform -1 0 2930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__933_
timestamp 0
transform -1 0 2870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__934_
timestamp 0
transform -1 0 2450 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__935_
timestamp 0
transform -1 0 770 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__936_
timestamp 0
transform -1 0 1210 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__937_
timestamp 0
transform -1 0 710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__957_
timestamp 0
transform 1 0 1850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__958_
timestamp 0
transform -1 0 1250 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__959_
timestamp 0
transform -1 0 1710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__960_
timestamp 0
transform 1 0 1510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__961_
timestamp 0
transform 1 0 1010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__962_
timestamp 0
transform -1 0 410 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__963_
timestamp 0
transform -1 0 1190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__964_
timestamp 0
transform 1 0 2070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__965_
timestamp 0
transform 1 0 1550 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__966_
timestamp 0
transform 1 0 1730 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__967_
timestamp 0
transform 1 0 1570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__968_
timestamp 0
transform -1 0 3030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__969_
timestamp 0
transform -1 0 6090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__970_
timestamp 0
transform -1 0 6410 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__971_
timestamp 0
transform 1 0 5910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__972_
timestamp 0
transform -1 0 5750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__973_
timestamp 0
transform 1 0 5410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__974_
timestamp 0
transform 1 0 3250 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__975_
timestamp 0
transform 1 0 2930 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__976_
timestamp 0
transform -1 0 6530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__977_
timestamp 0
transform 1 0 5770 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__978_
timestamp 0
transform 1 0 5610 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__979_
timestamp 0
transform -1 0 5450 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__980_
timestamp 0
transform 1 0 5270 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__981_
timestamp 0
transform 1 0 3510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__982_
timestamp 0
transform -1 0 3530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__983_
timestamp 0
transform -1 0 5330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__984_
timestamp 0
transform 1 0 3910 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__985_
timestamp 0
transform -1 0 4130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__986_
timestamp 0
transform -1 0 3270 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__987_
timestamp 0
transform -1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__988_
timestamp 0
transform 1 0 3650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__989_
timestamp 0
transform -1 0 4490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__990_
timestamp 0
transform 1 0 2910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__991_
timestamp 0
transform -1 0 6370 0 1 790
box -6 -8 26 268
use FILL  FILL_3__992_
timestamp 0
transform -1 0 6250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__993_
timestamp 0
transform 1 0 6010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__994_
timestamp 0
transform 1 0 6190 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__995_
timestamp 0
transform 1 0 4230 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__996_
timestamp 0
transform 1 0 4290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__997_
timestamp 0
transform -1 0 4270 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__998_
timestamp 0
transform 1 0 5570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__999_
timestamp 0
transform 1 0 6070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1000_
timestamp 0
transform -1 0 6830 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1001_
timestamp 0
transform -1 0 6010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1002_
timestamp 0
transform -1 0 5850 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1003_
timestamp 0
transform -1 0 5690 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1004_
timestamp 0
transform -1 0 4790 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1005_
timestamp 0
transform 1 0 6010 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1006_
timestamp 0
transform -1 0 5570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1007_
timestamp 0
transform -1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1008_
timestamp 0
transform -1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1009_
timestamp 0
transform -1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1010_
timestamp 0
transform -1 0 5150 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1011_
timestamp 0
transform 1 0 4950 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1012_
timestamp 0
transform 1 0 4710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1013_
timestamp 0
transform 1 0 4870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1014_
timestamp 0
transform -1 0 5350 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1015_
timestamp 0
transform -1 0 5530 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1016_
timestamp 0
transform 1 0 5390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1017_
timestamp 0
transform -1 0 4810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1018_
timestamp 0
transform -1 0 4650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1019_
timestamp 0
transform -1 0 5290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1020_
timestamp 0
transform -1 0 5190 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1021_
timestamp 0
transform -1 0 3910 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1022_
timestamp 0
transform 1 0 3730 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1023_
timestamp 0
transform -1 0 3010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1024_
timestamp 0
transform -1 0 2690 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1025_
timestamp 0
transform -1 0 4090 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1026_
timestamp 0
transform 1 0 3670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1027_
timestamp 0
transform 1 0 2930 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1028_
timestamp 0
transform 1 0 6290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1029_
timestamp 0
transform 1 0 4870 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1030_
timestamp 0
transform 1 0 3790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1031_
timestamp 0
transform -1 0 6910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1032_
timestamp 0
transform 1 0 4590 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1033_
timestamp 0
transform 1 0 4090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1034_
timestamp 0
transform 1 0 3890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1035_
timestamp 0
transform -1 0 4450 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1036_
timestamp 0
transform -1 0 4270 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1037_
timestamp 0
transform 1 0 6410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1038_
timestamp 0
transform 1 0 3950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1039_
timestamp 0
transform -1 0 4550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1040_
timestamp 0
transform -1 0 4710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1041_
timestamp 0
transform 1 0 4030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1042_
timestamp 0
transform -1 0 4210 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1043_
timestamp 0
transform -1 0 4370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1044_
timestamp 0
transform 1 0 3730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1045_
timestamp 0
transform -1 0 4430 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1046_
timestamp 0
transform -1 0 2630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1047_
timestamp 0
transform 1 0 4230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1048_
timestamp 0
transform -1 0 4070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1049_
timestamp 0
transform -1 0 3810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1050_
timestamp 0
transform 1 0 3310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1051_
timestamp 0
transform -1 0 3510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1052_
timestamp 0
transform -1 0 4610 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1053_
timestamp 0
transform -1 0 4090 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1054_
timestamp 0
transform 1 0 3730 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1055_
timestamp 0
transform -1 0 3870 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1056_
timestamp 0
transform -1 0 3930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1057_
timestamp 0
transform 1 0 3730 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1058_
timestamp 0
transform -1 0 3570 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1059_
timestamp 0
transform -1 0 3090 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1060_
timestamp 0
transform 1 0 3410 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1061_
timestamp 0
transform -1 0 3590 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1062_
timestamp 0
transform -1 0 3450 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1063_
timestamp 0
transform 1 0 550 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1064_
timestamp 0
transform 1 0 710 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1065_
timestamp 0
transform 1 0 1110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1066_
timestamp 0
transform 1 0 810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1067_
timestamp 0
transform -1 0 970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1068_
timestamp 0
transform -1 0 1070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1069_
timestamp 0
transform -1 0 910 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1070_
timestamp 0
transform -1 0 1350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1071_
timestamp 0
transform 1 0 2430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1072_
timestamp 0
transform -1 0 3270 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1073_
timestamp 0
transform -1 0 3090 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1074_
timestamp 0
transform -1 0 2770 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1075_
timestamp 0
transform 1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1076_
timestamp 0
transform -1 0 1410 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1077_
timestamp 0
transform 1 0 1230 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1078_
timestamp 0
transform -1 0 3190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1079_
timestamp 0
transform -1 0 2850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1080_
timestamp 0
transform 1 0 1850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1081_
timestamp 0
transform -1 0 2710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1082_
timestamp 0
transform 1 0 1890 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1083_
timestamp 0
transform -1 0 2370 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1084_
timestamp 0
transform 1 0 1510 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1085_
timestamp 0
transform -1 0 1550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1086_
timestamp 0
transform 1 0 1070 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1087_
timestamp 0
transform -1 0 1550 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1088_
timestamp 0
transform -1 0 1230 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1089_
timestamp 0
transform 1 0 1350 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1090_
timestamp 0
transform -1 0 970 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1091_
timestamp 0
transform 1 0 430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1092_
timestamp 0
transform 1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1093_
timestamp 0
transform -1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1094_
timestamp 0
transform 1 0 70 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1095_
timestamp 0
transform 1 0 930 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1096_
timestamp 0
transform -1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1097_
timestamp 0
transform 1 0 750 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1098_
timestamp 0
transform -1 0 90 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1099_
timestamp 0
transform 1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1100_
timestamp 0
transform -1 0 1930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1101_
timestamp 0
transform -1 0 2470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1102_
timestamp 0
transform 1 0 2070 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1103_
timestamp 0
transform -1 0 2290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1104_
timestamp 0
transform -1 0 1190 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1105_
timestamp 0
transform -1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1106_
timestamp 0
transform -1 0 890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1107_
timestamp 0
transform -1 0 990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1108_
timestamp 0
transform 1 0 1030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1109_
timestamp 0
transform -1 0 630 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1110_
timestamp 0
transform -1 0 730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1111_
timestamp 0
transform -1 0 730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1112_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1113_
timestamp 0
transform 1 0 550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1114_
timestamp 0
transform -1 0 310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1115_
timestamp 0
transform -1 0 250 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1116_
timestamp 0
transform 1 0 390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1117_
timestamp 0
transform 1 0 210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1118_
timestamp 0
transform 1 0 250 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1119_
timestamp 0
transform 1 0 2170 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1120_
timestamp 0
transform -1 0 2330 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1121_
timestamp 0
transform 1 0 2010 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1122_
timestamp 0
transform -1 0 2410 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1123_
timestamp 0
transform 1 0 2230 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1124_
timestamp 0
transform 1 0 1670 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1125_
timestamp 0
transform 1 0 1850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1126_
timestamp 0
transform 1 0 1750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1127_
timestamp 0
transform 1 0 1590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1128_
timestamp 0
transform 1 0 1510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1129_
timestamp 0
transform 1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1130_
timestamp 0
transform -1 0 1730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1131_
timestamp 0
transform -1 0 2070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1132_
timestamp 0
transform -1 0 2110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1133_
timestamp 0
transform -1 0 1930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1134_
timestamp 0
transform -1 0 1730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1135_
timestamp 0
transform 1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1136_
timestamp 0
transform -1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1137_
timestamp 0
transform -1 0 1070 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1138_
timestamp 0
transform -1 0 610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1139_
timestamp 0
transform -1 0 450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1140_
timestamp 0
transform -1 0 3890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1141_
timestamp 0
transform 1 0 4090 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1142_
timestamp 0
transform -1 0 4630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1143_
timestamp 0
transform 1 0 5530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1144_
timestamp 0
transform 1 0 6550 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1145_
timestamp 0
transform -1 0 5530 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1146_
timestamp 0
transform 1 0 4810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1147_
timestamp 0
transform -1 0 5010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1148_
timestamp 0
transform -1 0 4650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1149_
timestamp 0
transform 1 0 5690 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1150_
timestamp 0
transform -1 0 5210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1151_
timestamp 0
transform -1 0 5190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1152_
timestamp 0
transform -1 0 4470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1153_
timestamp 0
transform -1 0 4310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1154_
timestamp 0
transform -1 0 6370 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1155_
timestamp 0
transform -1 0 6790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1156_
timestamp 0
transform 1 0 3230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1157_
timestamp 0
transform 1 0 3550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1158_
timestamp 0
transform -1 0 6150 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1159_
timestamp 0
transform 1 0 5350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1160_
timestamp 0
transform 1 0 5270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1161_
timestamp 0
transform 1 0 4210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1162_
timestamp 0
transform -1 0 5070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1163_
timestamp 0
transform 1 0 4850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1164_
timestamp 0
transform 1 0 5090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1165_
timestamp 0
transform 1 0 5110 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1166_
timestamp 0
transform -1 0 4870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1167_
timestamp 0
transform -1 0 5970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1168_
timestamp 0
transform 1 0 5830 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1169_
timestamp 0
transform 1 0 3870 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1170_
timestamp 0
transform 1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1171_
timestamp 0
transform 1 0 2910 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1172_
timestamp 0
transform -1 0 3090 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1173_
timestamp 0
transform 1 0 3050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1174_
timestamp 0
transform 1 0 3550 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1175_
timestamp 0
transform 1 0 3710 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1176_
timestamp 0
transform -1 0 4050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1177_
timestamp 0
transform 1 0 4370 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1178_
timestamp 0
transform -1 0 5050 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1179_
timestamp 0
transform 1 0 5350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1180_
timestamp 0
transform 1 0 4750 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1181_
timestamp 0
transform 1 0 5290 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1182_
timestamp 0
transform 1 0 5190 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1183_
timestamp 0
transform -1 0 5410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1184_
timestamp 0
transform 1 0 5190 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform -1 0 4570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1186_
timestamp 0
transform -1 0 5590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1187_
timestamp 0
transform -1 0 5170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1188_
timestamp 0
transform -1 0 4830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1189_
timestamp 0
transform -1 0 4530 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1190_
timestamp 0
transform 1 0 5710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1191_
timestamp 0
transform 1 0 6170 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1192_
timestamp 0
transform 1 0 4290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1193_
timestamp 0
transform -1 0 4350 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1194_
timestamp 0
transform -1 0 3670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1195_
timestamp 0
transform 1 0 3690 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1196_
timestamp 0
transform 1 0 3510 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1197_
timestamp 0
transform 1 0 3150 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1198_
timestamp 0
transform 1 0 3410 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1199_
timestamp 0
transform -1 0 3410 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1200_
timestamp 0
transform -1 0 2230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1201_
timestamp 0
transform 1 0 3570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1202_
timestamp 0
transform 1 0 3390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1203_
timestamp 0
transform -1 0 3250 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1204_
timestamp 0
transform 1 0 2550 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1205_
timestamp 0
transform 1 0 2450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1206_
timestamp 0
transform 1 0 2130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1207_
timestamp 0
transform 1 0 2750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1208_
timestamp 0
transform 1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1209_
timestamp 0
transform -1 0 3110 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1210_
timestamp 0
transform -1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1211_
timestamp 0
transform 1 0 2730 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1212_
timestamp 0
transform 1 0 4490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1213_
timestamp 0
transform 1 0 4650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1214_
timestamp 0
transform 1 0 4130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1215_
timestamp 0
transform -1 0 4030 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1216_
timestamp 0
transform 1 0 4710 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1217_
timestamp 0
transform 1 0 4170 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1218_
timestamp 0
transform -1 0 3870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1219_
timestamp 0
transform -1 0 3170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1220_
timestamp 0
transform 1 0 3790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1221_
timestamp 0
transform -1 0 3370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1222_
timestamp 0
transform 1 0 3350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1223_
timestamp 0
transform -1 0 3490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1224_
timestamp 0
transform 1 0 3610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1225_
timestamp 0
transform -1 0 3710 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1226_
timestamp 0
transform -1 0 3970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1227_
timestamp 0
transform 1 0 3310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1228_
timestamp 0
transform -1 0 3370 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1229_
timestamp 0
transform -1 0 3530 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1230_
timestamp 0
transform 1 0 2810 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1231_
timestamp 0
transform 1 0 2390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1232_
timestamp 0
transform 1 0 1970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1233_
timestamp 0
transform -1 0 1890 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1234_
timestamp 0
transform -1 0 2230 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1235_
timestamp 0
transform 1 0 2490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1236_
timestamp 0
transform -1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1237_
timestamp 0
transform 1 0 2850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1238_
timestamp 0
transform -1 0 1630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1239_
timestamp 0
transform -1 0 1830 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1240_
timestamp 0
transform 1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1241_
timestamp 0
transform -1 0 2410 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1242_
timestamp 0
transform -1 0 2010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1243_
timestamp 0
transform 1 0 2170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1244_
timestamp 0
transform 1 0 1310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1245_
timestamp 0
transform -1 0 1670 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1246_
timestamp 0
transform 1 0 1630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1247_
timestamp 0
transform -1 0 2750 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1248_
timestamp 0
transform 1 0 2550 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1249_
timestamp 0
transform -1 0 1530 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1250_
timestamp 0
transform -1 0 1470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1251_
timestamp 0
transform 1 0 1710 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1252_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1253_
timestamp 0
transform -1 0 2090 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1254_
timestamp 0
transform 1 0 1810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1255_
timestamp 0
transform 1 0 1890 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1256_
timestamp 0
transform -1 0 1710 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1257_
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1258_
timestamp 0
transform 1 0 2090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1259_
timestamp 0
transform 1 0 1850 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1260_
timestamp 0
transform -1 0 1470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1261_
timestamp 0
transform -1 0 1390 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1262_
timestamp 0
transform 1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1263_
timestamp 0
transform -1 0 2230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1264_
timestamp 0
transform -1 0 2070 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1265_
timestamp 0
transform -1 0 1910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1266_
timestamp 0
transform 1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1267_
timestamp 0
transform 1 0 2030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1268_
timestamp 0
transform -1 0 2250 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1269_
timestamp 0
transform 1 0 2210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1270_
timestamp 0
transform -1 0 2390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1271_
timestamp 0
transform 1 0 2410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1272_
timestamp 0
transform 1 0 2030 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1273_
timestamp 0
transform -1 0 2630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1274_
timestamp 0
transform -1 0 290 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1275_
timestamp 0
transform -1 0 450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1276_
timestamp 0
transform 1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1277_
timestamp 0
transform 1 0 410 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1278_
timestamp 0
transform -1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1279_
timestamp 0
transform 1 0 410 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1280_
timestamp 0
transform 1 0 230 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1281_
timestamp 0
transform -1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1282_
timestamp 0
transform -1 0 750 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1283_
timestamp 0
transform 1 0 590 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1284_
timestamp 0
transform 1 0 1550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1285_
timestamp 0
transform -1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1286_
timestamp 0
transform -1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1287_
timestamp 0
transform -1 0 1330 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1288_
timestamp 0
transform 1 0 1910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1289_
timestamp 0
transform -1 0 1130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1290_
timestamp 0
transform -1 0 1150 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1291_
timestamp 0
transform 1 0 550 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1292_
timestamp 0
transform -1 0 90 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1293_
timestamp 0
transform -1 0 90 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1294_
timestamp 0
transform -1 0 250 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1295_
timestamp 0
transform 1 0 570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1296_
timestamp 0
transform -1 0 810 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1297_
timestamp 0
transform 1 0 1750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1298_
timestamp 0
transform -1 0 1490 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1299_
timestamp 0
transform -1 0 990 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1300_
timestamp 0
transform -1 0 1670 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1301_
timestamp 0
transform 1 0 2150 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1302_
timestamp 0
transform 1 0 1970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1303_
timestamp 0
transform 1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1304_
timestamp 0
transform -1 0 2590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1305_
timestamp 0
transform -1 0 1550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1306_
timestamp 0
transform -1 0 1390 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1307_
timestamp 0
transform 1 0 1370 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1308_
timestamp 0
transform 1 0 1350 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1309_
timestamp 0
transform -1 0 5250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1310_
timestamp 0
transform 1 0 2950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1311_
timestamp 0
transform 1 0 2590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1312_
timestamp 0
transform 1 0 1670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1313_
timestamp 0
transform 1 0 1710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1314_
timestamp 0
transform 1 0 2770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1315_
timestamp 0
transform -1 0 4990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1316_
timestamp 0
transform 1 0 5650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1317_
timestamp 0
transform 1 0 5530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1318_
timestamp 0
transform 1 0 5810 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1319_
timestamp 0
transform -1 0 5710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1320_
timestamp 0
transform -1 0 6390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1321_
timestamp 0
transform -1 0 6690 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1322_
timestamp 0
transform -1 0 6750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1323_
timestamp 0
transform 1 0 6750 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1324_
timestamp 0
transform 1 0 5010 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1325_
timestamp 0
transform -1 0 5490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1326_
timestamp 0
transform 1 0 5330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1327_
timestamp 0
transform 1 0 5530 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1328_
timestamp 0
transform 1 0 5710 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1329_
timestamp 0
transform 1 0 5890 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1330_
timestamp 0
transform 1 0 5430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1331_
timestamp 0
transform 1 0 6430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1332_
timestamp 0
transform -1 0 5790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1333_
timestamp 0
transform 1 0 5930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1334_
timestamp 0
transform -1 0 6170 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1335_
timestamp 0
transform 1 0 6390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1336_
timestamp 0
transform 1 0 6550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1337_
timestamp 0
transform -1 0 6730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1338_
timestamp 0
transform -1 0 6730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1339_
timestamp 0
transform -1 0 6830 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1340_
timestamp 0
transform 1 0 6490 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1341_
timestamp 0
transform -1 0 6850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1342_
timestamp 0
transform 1 0 5610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1343_
timestamp 0
transform 1 0 6570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1344_
timestamp 0
transform -1 0 6750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1345_
timestamp 0
transform 1 0 6630 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1346_
timestamp 0
transform 1 0 6570 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1347_
timestamp 0
transform 1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1348_
timestamp 0
transform 1 0 6330 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1349_
timestamp 0
transform -1 0 6570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1350_
timestamp 0
transform 1 0 6510 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1351_
timestamp 0
transform 1 0 5510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1352_
timestamp 0
transform 1 0 5730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1353_
timestamp 0
transform -1 0 5910 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1354_
timestamp 0
transform 1 0 6070 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1355_
timestamp 0
transform 1 0 6370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1356_
timestamp 0
transform 1 0 6550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1357_
timestamp 0
transform -1 0 6210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1358_
timestamp 0
transform 1 0 6010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1359_
timestamp 0
transform 1 0 6470 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1360_
timestamp 0
transform 1 0 6090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1361_
timestamp 0
transform -1 0 6270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1362_
timestamp 0
transform -1 0 6710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1363_
timestamp 0
transform 1 0 6650 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1364_
timestamp 0
transform -1 0 6730 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1365_
timestamp 0
transform -1 0 6830 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1366_
timestamp 0
transform -1 0 6070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1367_
timestamp 0
transform -1 0 6230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1368_
timestamp 0
transform -1 0 5350 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1369_
timestamp 0
transform -1 0 4550 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1370_
timestamp 0
transform 1 0 3870 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1371_
timestamp 0
transform 1 0 4210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1372_
timestamp 0
transform -1 0 5110 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1373_
timestamp 0
transform -1 0 4690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1374_
timestamp 0
transform 1 0 5810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1375_
timestamp 0
transform -1 0 5370 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1376_
timestamp 0
transform 1 0 6530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1377_
timestamp 0
transform -1 0 6850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1378_
timestamp 0
transform -1 0 6610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1379_
timestamp 0
transform -1 0 6670 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1380_
timestamp 0
transform 1 0 6170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1381_
timestamp 0
transform -1 0 6370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1382_
timestamp 0
transform -1 0 5650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1383_
timestamp 0
transform 1 0 4790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1384_
timestamp 0
transform -1 0 4970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1385_
timestamp 0
transform -1 0 5210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1386_
timestamp 0
transform -1 0 5010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1387_
timestamp 0
transform -1 0 5010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1388_
timestamp 0
transform 1 0 4290 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1389_
timestamp 0
transform -1 0 4510 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1390_
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1391_
timestamp 0
transform -1 0 1370 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1392_
timestamp 0
transform -1 0 1390 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1393_
timestamp 0
transform -1 0 890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1394_
timestamp 0
transform 1 0 950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1395_
timestamp 0
transform -1 0 4130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1396_
timestamp 0
transform -1 0 3010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1397_
timestamp 0
transform 1 0 2810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1398_
timestamp 0
transform 1 0 4350 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1399_
timestamp 0
transform 1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1400_
timestamp 0
transform 1 0 5990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1401_
timestamp 0
transform -1 0 5910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1402_
timestamp 0
transform -1 0 4450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1403_
timestamp 0
transform 1 0 4750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1404_
timestamp 0
transform 1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1405_
timestamp 0
transform 1 0 4890 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1406_
timestamp 0
transform -1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1407_
timestamp 0
transform -1 0 5130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1408_
timestamp 0
transform 1 0 5050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1409_
timestamp 0
transform -1 0 5070 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1410_
timestamp 0
transform 1 0 4330 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1411_
timestamp 0
transform -1 0 6090 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1412_
timestamp 0
transform 1 0 5350 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1413_
timestamp 0
transform 1 0 6230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1414_
timestamp 0
transform -1 0 6570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1415_
timestamp 0
transform -1 0 6270 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1416_
timestamp 0
transform -1 0 6410 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1417_
timestamp 0
transform -1 0 5490 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1418_
timestamp 0
transform -1 0 5030 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1419_
timestamp 0
transform -1 0 4410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform -1 0 4790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1421_
timestamp 0
transform -1 0 4610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1422_
timestamp 0
transform 1 0 4390 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1423_
timestamp 0
transform -1 0 4610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1424_
timestamp 0
transform 1 0 4010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1425_
timestamp 0
transform -1 0 4230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1426_
timestamp 0
transform 1 0 770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1427_
timestamp 0
transform 1 0 590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1428_
timestamp 0
transform 1 0 2370 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1429_
timestamp 0
transform -1 0 4050 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1430_
timestamp 0
transform -1 0 4710 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1431_
timestamp 0
transform -1 0 4890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1432_
timestamp 0
transform -1 0 4710 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1433_
timestamp 0
transform -1 0 4890 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1434_
timestamp 0
transform 1 0 2390 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1435_
timestamp 0
transform 1 0 4690 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1436_
timestamp 0
transform -1 0 2270 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1437_
timestamp 0
transform 1 0 2350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1438_
timestamp 0
transform 1 0 2410 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1439_
timestamp 0
transform 1 0 2670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1440_
timestamp 0
transform 1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1441_
timestamp 0
transform -1 0 2850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1442_
timestamp 0
transform 1 0 2750 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1443_
timestamp 0
transform 1 0 2210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1444_
timestamp 0
transform 1 0 1690 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1445_
timestamp 0
transform 1 0 1730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1446_
timestamp 0
transform 1 0 2390 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1447_
timestamp 0
transform 1 0 2510 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1448_
timestamp 0
transform 1 0 2890 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1449_
timestamp 0
transform 1 0 4370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1450_
timestamp 0
transform -1 0 4210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1451_
timestamp 0
transform 1 0 4830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1452_
timestamp 0
transform 1 0 2830 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1453_
timestamp 0
transform 1 0 2650 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1454_
timestamp 0
transform -1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1455_
timestamp 0
transform -1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1456_
timestamp 0
transform 1 0 5270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1457_
timestamp 0
transform -1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1458_
timestamp 0
transform -1 0 5450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1459_
timestamp 0
transform 1 0 3670 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1460_
timestamp 0
transform 1 0 4430 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1461_
timestamp 0
transform 1 0 3490 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1462_
timestamp 0
transform -1 0 3130 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1463_
timestamp 0
transform 1 0 2790 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1464_
timestamp 0
transform 1 0 2230 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1465_
timestamp 0
transform 1 0 2530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1466_
timestamp 0
transform -1 0 2710 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1467_
timestamp 0
transform 1 0 3010 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1468_
timestamp 0
transform 1 0 3150 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1469_
timestamp 0
transform 1 0 2610 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1470_
timestamp 0
transform 1 0 3610 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1471_
timestamp 0
transform -1 0 3850 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1472_
timestamp 0
transform -1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1473_
timestamp 0
transform 1 0 4050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1474_
timestamp 0
transform 1 0 5150 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1475_
timestamp 0
transform -1 0 4250 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1476_
timestamp 0
transform -1 0 4830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1477_
timestamp 0
transform 1 0 4550 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1478_
timestamp 0
transform -1 0 4650 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1479_
timestamp 0
transform -1 0 4410 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1480_
timestamp 0
transform 1 0 5990 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1481_
timestamp 0
transform 1 0 5830 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1482_
timestamp 0
transform -1 0 5630 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1483_
timestamp 0
transform 1 0 3610 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1484_
timestamp 0
transform -1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1485_
timestamp 0
transform 1 0 3030 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1486_
timestamp 0
transform 1 0 3470 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1487_
timestamp 0
transform 1 0 3310 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1488_
timestamp 0
transform 1 0 2990 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1489_
timestamp 0
transform 1 0 2950 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1490_
timestamp 0
transform -1 0 3290 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1491_
timestamp 0
transform -1 0 4710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1492_
timestamp 0
transform -1 0 4610 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1493_
timestamp 0
transform -1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1494_
timestamp 0
transform 1 0 3530 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1495_
timestamp 0
transform 1 0 3710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1496_
timestamp 0
transform -1 0 4450 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1497_
timestamp 0
transform 1 0 4970 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1498_
timestamp 0
transform 1 0 4470 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1499_
timestamp 0
transform 1 0 4290 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1500_
timestamp 0
transform -1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1501_
timestamp 0
transform 1 0 4110 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1502_
timestamp 0
transform 1 0 4210 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1503_
timestamp 0
transform 1 0 4210 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1504_
timestamp 0
transform -1 0 4530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1505_
timestamp 0
transform -1 0 4170 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1506_
timestamp 0
transform 1 0 4370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1507_
timestamp 0
transform 1 0 4610 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1508_
timestamp 0
transform 1 0 4810 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1509_
timestamp 0
transform 1 0 2210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1510_
timestamp 0
transform -1 0 2610 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1511_
timestamp 0
transform 1 0 2390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1512_
timestamp 0
transform 1 0 2510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1513_
timestamp 0
transform -1 0 2590 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1514_
timestamp 0
transform -1 0 2590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1515_
timestamp 0
transform 1 0 2690 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1516_
timestamp 0
transform -1 0 2870 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1517_
timestamp 0
transform 1 0 3750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1518_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1519_
timestamp 0
transform -1 0 4210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1520_
timestamp 0
transform 1 0 3190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1521_
timestamp 0
transform -1 0 4010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1522_
timestamp 0
transform -1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1523_
timestamp 0
transform 1 0 3010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1524_
timestamp 0
transform -1 0 4070 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1525_
timestamp 0
transform 1 0 3190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1526_
timestamp 0
transform 1 0 3350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1527_
timestamp 0
transform 1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1528_
timestamp 0
transform -1 0 3030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1529_
timestamp 0
transform -1 0 1270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1530_
timestamp 0
transform 1 0 1410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1531_
timestamp 0
transform 1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1532_
timestamp 0
transform -1 0 1910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1533_
timestamp 0
transform -1 0 2070 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1534_
timestamp 0
transform -1 0 2370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1535_
timestamp 0
transform -1 0 2750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1536_
timestamp 0
transform -1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1537_
timestamp 0
transform 1 0 2490 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1538_
timestamp 0
transform 1 0 3890 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1539_
timestamp 0
transform -1 0 3270 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1540_
timestamp 0
transform 1 0 1830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1541_
timestamp 0
transform -1 0 3450 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1542_
timestamp 0
transform 1 0 2030 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1543_
timestamp 0
transform 1 0 3890 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1544_
timestamp 0
transform 1 0 3150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1545_
timestamp 0
transform 1 0 2450 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1546_
timestamp 0
transform 1 0 3590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1547_
timestamp 0
transform 1 0 4750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1548_
timestamp 0
transform 1 0 3890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1549_
timestamp 0
transform -1 0 4890 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1550_
timestamp 0
transform 1 0 5010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1551_
timestamp 0
transform -1 0 5210 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1552_
timestamp 0
transform 1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1553_
timestamp 0
transform -1 0 4530 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1554_
timestamp 0
transform 1 0 5230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1555_
timestamp 0
transform 1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1556_
timestamp 0
transform -1 0 5050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1557_
timestamp 0
transform -1 0 4850 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1558_
timestamp 0
transform -1 0 3830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1559_
timestamp 0
transform 1 0 4970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1560_
timestamp 0
transform -1 0 5010 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1561_
timestamp 0
transform -1 0 4650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1562_
timestamp 0
transform 1 0 3970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1563_
timestamp 0
transform -1 0 4170 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1564_
timestamp 0
transform -1 0 4870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1565_
timestamp 0
transform 1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1566_
timestamp 0
transform 1 0 3490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1567_
timestamp 0
transform -1 0 3010 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1568_
timestamp 0
transform 1 0 3650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1569_
timestamp 0
transform -1 0 3310 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1570_
timestamp 0
transform 1 0 3130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1571_
timestamp 0
transform 1 0 3190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1572_
timestamp 0
transform 1 0 3370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1573_
timestamp 0
transform 1 0 3930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1574_
timestamp 0
transform -1 0 4470 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1575_
timestamp 0
transform -1 0 3970 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1576_
timestamp 0
transform -1 0 4130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1577_
timestamp 0
transform -1 0 3450 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1578_
timestamp 0
transform -1 0 3810 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1579_
timestamp 0
transform 1 0 3610 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1580_
timestamp 0
transform 1 0 3690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1581_
timestamp 0
transform -1 0 3890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1582_
timestamp 0
transform 1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1583_
timestamp 0
transform -1 0 4070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1584_
timestamp 0
transform -1 0 4630 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1585_
timestamp 0
transform 1 0 4230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1586_
timestamp 0
transform -1 0 4710 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1587_
timestamp 0
transform -1 0 3290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1588_
timestamp 0
transform -1 0 3150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1589_
timestamp 0
transform -1 0 4450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1590_
timestamp 0
transform -1 0 4310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1591_
timestamp 0
transform 1 0 4270 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1592_
timestamp 0
transform 1 0 4110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1593_
timestamp 0
transform 1 0 2630 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1594_
timestamp 0
transform 1 0 2810 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1595_
timestamp 0
transform -1 0 3010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1596_
timestamp 0
transform -1 0 3210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1597_
timestamp 0
transform 1 0 3010 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1598_
timestamp 0
transform -1 0 3370 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1599_
timestamp 0
transform -1 0 3710 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1600_
timestamp 0
transform 1 0 3510 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1601_
timestamp 0
transform -1 0 3450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1602_
timestamp 0
transform -1 0 2910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1603_
timestamp 0
transform -1 0 3090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1604_
timestamp 0
transform -1 0 3270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1605_
timestamp 0
transform 1 0 4110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1606_
timestamp 0
transform 1 0 6330 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1607_
timestamp 0
transform 1 0 6270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1608_
timestamp 0
transform -1 0 6450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1609_
timestamp 0
transform 1 0 6210 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1610_
timestamp 0
transform 1 0 6610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1611_
timestamp 0
transform 1 0 5650 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1612_
timestamp 0
transform -1 0 6870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1613_
timestamp 0
transform -1 0 6490 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1614_
timestamp 0
transform -1 0 6310 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1615_
timestamp 0
transform -1 0 6130 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1616_
timestamp 0
transform 1 0 5930 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1617_
timestamp 0
transform 1 0 5670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1618_
timestamp 0
transform -1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1619_
timestamp 0
transform 1 0 5370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1620_
timestamp 0
transform -1 0 6150 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1621_
timestamp 0
transform 1 0 5370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1622_
timestamp 0
transform 1 0 6790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1623_
timestamp 0
transform 1 0 6450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1624_
timestamp 0
transform -1 0 6850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1625_
timestamp 0
transform -1 0 6590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1626_
timestamp 0
transform 1 0 6570 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1627_
timestamp 0
transform 1 0 6410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1628_
timestamp 0
transform -1 0 6210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1629_
timestamp 0
transform 1 0 5990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1630_
timestamp 0
transform 1 0 6710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1631_
timestamp 0
transform -1 0 6770 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1632_
timestamp 0
transform -1 0 6650 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1633_
timestamp 0
transform -1 0 6670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1634_
timestamp 0
transform -1 0 6490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1635_
timestamp 0
transform 1 0 6290 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1636_
timestamp 0
transform -1 0 6470 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1637_
timestamp 0
transform 1 0 6110 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1638_
timestamp 0
transform -1 0 6510 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1639_
timestamp 0
transform 1 0 6370 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1640_
timestamp 0
transform 1 0 5710 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1641_
timestamp 0
transform -1 0 6770 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1642_
timestamp 0
transform -1 0 6270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1643_
timestamp 0
transform -1 0 6570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1644_
timestamp 0
transform -1 0 6270 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1645_
timestamp 0
transform 1 0 6590 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1646_
timestamp 0
transform -1 0 6730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1647_
timestamp 0
transform -1 0 6050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1648_
timestamp 0
transform 1 0 5830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1649_
timestamp 0
transform -1 0 6730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1650_
timestamp 0
transform -1 0 6730 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1651_
timestamp 0
transform -1 0 6290 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1652_
timestamp 0
transform -1 0 6510 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1653_
timestamp 0
transform 1 0 5630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1654_
timestamp 0
transform 1 0 6410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1655_
timestamp 0
transform 1 0 6390 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1656_
timestamp 0
transform 1 0 6570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1657_
timestamp 0
transform -1 0 6830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1658_
timestamp 0
transform 1 0 6170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1659_
timestamp 0
transform -1 0 6870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1660_
timestamp 0
transform -1 0 6650 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1661_
timestamp 0
transform -1 0 6830 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1662_
timestamp 0
transform -1 0 6470 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1663_
timestamp 0
transform 1 0 6050 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1664_
timestamp 0
transform 1 0 6230 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1665_
timestamp 0
transform -1 0 6350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1666_
timestamp 0
transform -1 0 6670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1667_
timestamp 0
transform 1 0 6430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1668_
timestamp 0
transform 1 0 6730 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1669_
timestamp 0
transform -1 0 6010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1670_
timestamp 0
transform 1 0 5870 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1671_
timestamp 0
transform 1 0 5550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1672_
timestamp 0
transform -1 0 6110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1673_
timestamp 0
transform 1 0 5730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1674_
timestamp 0
transform -1 0 5930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1675_
timestamp 0
transform 1 0 4030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1676_
timestamp 0
transform 1 0 5210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1677_
timestamp 0
transform 1 0 5130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1711_
timestamp 0
transform -1 0 90 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1712_
timestamp 0
transform -1 0 90 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1713_
timestamp 0
transform -1 0 1090 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1714_
timestamp 0
transform 1 0 230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1715_
timestamp 0
transform -1 0 90 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1716_
timestamp 0
transform -1 0 90 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1717_
timestamp 0
transform 1 0 390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1718_
timestamp 0
transform -1 0 90 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1719_
timestamp 0
transform 1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1720_
timestamp 0
transform -1 0 90 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1721_
timestamp 0
transform -1 0 250 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1722_
timestamp 0
transform -1 0 90 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1723_
timestamp 0
transform 1 0 1530 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1724_
timestamp 0
transform 1 0 390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_3__1725_
timestamp 0
transform -1 0 450 0 1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert0
timestamp 0
transform -1 0 90 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert1
timestamp 0
transform 1 0 270 0 1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert2
timestamp 0
transform 1 0 230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform 1 0 390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform 1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform -1 0 5410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform 1 0 5650 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform -1 0 2510 0 1 790
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform 1 0 3370 0 1 1310
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert4
timestamp 0
transform 1 0 4990 0 1 790
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert5
timestamp 0
transform -1 0 1950 0 1 4950
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert6
timestamp 0
transform -1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert7
timestamp 0
transform 1 0 530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert8
timestamp 0
transform -1 0 430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert9
timestamp 0
transform 1 0 2610 0 1 1830
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert10
timestamp 0
transform -1 0 3590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__828_
timestamp 0
transform 1 0 870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__829_
timestamp 0
transform 1 0 1550 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__830_
timestamp 0
transform -1 0 2410 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__831_
timestamp 0
transform -1 0 1390 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__832_
timestamp 0
transform 1 0 2310 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__833_
timestamp 0
transform 1 0 2010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__834_
timestamp 0
transform -1 0 1630 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__835_
timestamp 0
transform -1 0 1710 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__836_
timestamp 0
transform -1 0 1030 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__838_
timestamp 0
transform -1 0 750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__839_
timestamp 0
transform -1 0 950 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__840_
timestamp 0
transform 1 0 90 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__841_
timestamp 0
transform -1 0 110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__842_
timestamp 0
transform 1 0 90 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__843_
timestamp 0
transform -1 0 270 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__844_
timestamp 0
transform 1 0 730 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__845_
timestamp 0
transform 1 0 270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__846_
timestamp 0
transform -1 0 790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__847_
timestamp 0
transform -1 0 950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__848_
timestamp 0
transform -1 0 610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__849_
timestamp 0
transform 1 0 250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__850_
timestamp 0
transform -1 0 270 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__851_
timestamp 0
transform -1 0 910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__852_
timestamp 0
transform -1 0 730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__853_
timestamp 0
transform 1 0 610 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__854_
timestamp 0
transform -1 0 110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__855_
timestamp 0
transform -1 0 590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__856_
timestamp 0
transform -1 0 790 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__857_
timestamp 0
transform 1 0 1050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__858_
timestamp 0
transform -1 0 530 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__859_
timestamp 0
transform 1 0 90 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__860_
timestamp 0
transform 1 0 1110 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__861_
timestamp 0
transform 1 0 870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__862_
timestamp 0
transform -1 0 750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__863_
timestamp 0
transform -1 0 570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__864_
timestamp 0
transform 1 0 870 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__865_
timestamp 0
transform 1 0 450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__866_
timestamp 0
transform -1 0 1410 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__867_
timestamp 0
transform 1 0 1030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__868_
timestamp 0
transform 1 0 1050 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__869_
timestamp 0
transform -1 0 1250 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__870_
timestamp 0
transform 1 0 1170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__871_
timestamp 0
transform -1 0 1470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__872_
timestamp 0
transform -1 0 910 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__873_
timestamp 0
transform 1 0 1070 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__874_
timestamp 0
transform 1 0 1050 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__875_
timestamp 0
transform 1 0 1290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__876_
timestamp 0
transform -1 0 1210 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__877_
timestamp 0
transform 1 0 1350 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__878_
timestamp 0
transform -1 0 890 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__879_
timestamp 0
transform -1 0 110 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__880_
timestamp 0
transform 1 0 1210 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__881_
timestamp 0
transform 1 0 250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__882_
timestamp 0
transform -1 0 250 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__883_
timestamp 0
transform 1 0 890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__884_
timestamp 0
transform -1 0 1050 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__886_
timestamp 0
transform -1 0 890 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__887_
timestamp 0
transform 1 0 890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__888_
timestamp 0
transform -1 0 710 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__889_
timestamp 0
transform 1 0 550 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__890_
timestamp 0
transform -1 0 730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__891_
timestamp 0
transform 1 0 370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__892_
timestamp 0
transform -1 0 550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__893_
timestamp 0
transform -1 0 250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__894_
timestamp 0
transform -1 0 570 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__895_
timestamp 0
transform -1 0 730 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__896_
timestamp 0
transform 1 0 1850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__897_
timestamp 0
transform -1 0 2570 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__898_
timestamp 0
transform -1 0 2230 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__899_
timestamp 0
transform 1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__900_
timestamp 0
transform -1 0 1790 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__901_
timestamp 0
transform 1 0 1670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__902_
timestamp 0
transform -1 0 1710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__903_
timestamp 0
transform -1 0 1850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__904_
timestamp 0
transform -1 0 1530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__905_
timestamp 0
transform -1 0 1450 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__906_
timestamp 0
transform 1 0 1250 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__907_
timestamp 0
transform 1 0 1830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__908_
timestamp 0
transform 1 0 2330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__909_
timestamp 0
transform 1 0 2050 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__910_
timestamp 0
transform -1 0 1890 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__911_
timestamp 0
transform 1 0 1650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__912_
timestamp 0
transform -1 0 1790 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__913_
timestamp 0
transform 1 0 2890 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__914_
timestamp 0
transform -1 0 3230 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__915_
timestamp 0
transform 1 0 2150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__916_
timestamp 0
transform -1 0 2150 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__917_
timestamp 0
transform 1 0 1590 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__918_
timestamp 0
transform 1 0 1990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__919_
timestamp 0
transform -1 0 3050 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__920_
timestamp 0
transform -1 0 3310 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__921_
timestamp 0
transform 1 0 2690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__922_
timestamp 0
transform -1 0 2530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__923_
timestamp 0
transform -1 0 2350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__924_
timestamp 0
transform 1 0 1950 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__925_
timestamp 0
transform 1 0 2630 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__926_
timestamp 0
transform -1 0 2790 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__927_
timestamp 0
transform -1 0 3450 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__928_
timestamp 0
transform -1 0 3130 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__929_
timestamp 0
transform -1 0 2610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__930_
timestamp 0
transform -1 0 2430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__931_
timestamp 0
transform -1 0 970 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__932_
timestamp 0
transform -1 0 2950 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__934_
timestamp 0
transform -1 0 2470 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__935_
timestamp 0
transform -1 0 790 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__936_
timestamp 0
transform -1 0 1230 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__937_
timestamp 0
transform -1 0 730 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__957_
timestamp 0
transform 1 0 1870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__958_
timestamp 0
transform -1 0 1270 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__959_
timestamp 0
transform -1 0 1730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__960_
timestamp 0
transform 1 0 1530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__961_
timestamp 0
transform 1 0 1030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__962_
timestamp 0
transform -1 0 430 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__963_
timestamp 0
transform -1 0 1210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__964_
timestamp 0
transform 1 0 2090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__965_
timestamp 0
transform 1 0 1570 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__966_
timestamp 0
transform 1 0 1750 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__967_
timestamp 0
transform 1 0 1590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__968_
timestamp 0
transform -1 0 3050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__969_
timestamp 0
transform -1 0 6110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__970_
timestamp 0
transform -1 0 6430 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__971_
timestamp 0
transform 1 0 5930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__972_
timestamp 0
transform -1 0 5770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__973_
timestamp 0
transform 1 0 5430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__974_
timestamp 0
transform 1 0 3270 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__975_
timestamp 0
transform 1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__976_
timestamp 0
transform -1 0 6550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__977_
timestamp 0
transform 1 0 5790 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__978_
timestamp 0
transform 1 0 5630 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__979_
timestamp 0
transform -1 0 5470 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__980_
timestamp 0
transform 1 0 5290 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__981_
timestamp 0
transform 1 0 3530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__982_
timestamp 0
transform -1 0 3550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__983_
timestamp 0
transform -1 0 5350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__984_
timestamp 0
transform 1 0 3930 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__985_
timestamp 0
transform -1 0 4150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__986_
timestamp 0
transform -1 0 3290 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__987_
timestamp 0
transform -1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__988_
timestamp 0
transform 1 0 3670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__989_
timestamp 0
transform -1 0 4510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__990_
timestamp 0
transform 1 0 2930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__991_
timestamp 0
transform -1 0 6390 0 1 790
box -6 -8 26 268
use FILL  FILL_4__992_
timestamp 0
transform -1 0 6270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__993_
timestamp 0
transform 1 0 6030 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__994_
timestamp 0
transform 1 0 6210 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__995_
timestamp 0
transform 1 0 4250 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__996_
timestamp 0
transform 1 0 4310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__997_
timestamp 0
transform -1 0 4290 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__998_
timestamp 0
transform 1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__999_
timestamp 0
transform 1 0 6090 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1000_
timestamp 0
transform -1 0 6850 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1001_
timestamp 0
transform -1 0 6030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1002_
timestamp 0
transform -1 0 5870 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1003_
timestamp 0
transform -1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1004_
timestamp 0
transform -1 0 4810 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1005_
timestamp 0
transform 1 0 6030 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1006_
timestamp 0
transform -1 0 5590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1007_
timestamp 0
transform -1 0 5510 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1008_
timestamp 0
transform -1 0 5810 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1009_
timestamp 0
transform -1 0 5650 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1010_
timestamp 0
transform -1 0 5170 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1011_
timestamp 0
transform 1 0 4970 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1012_
timestamp 0
transform 1 0 4730 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1013_
timestamp 0
transform 1 0 4890 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1014_
timestamp 0
transform -1 0 5370 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1015_
timestamp 0
transform -1 0 5550 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1016_
timestamp 0
transform 1 0 5410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1017_
timestamp 0
transform -1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1018_
timestamp 0
transform -1 0 4670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1019_
timestamp 0
transform -1 0 5310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1020_
timestamp 0
transform -1 0 5210 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1021_
timestamp 0
transform -1 0 3930 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1022_
timestamp 0
transform 1 0 3750 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1023_
timestamp 0
transform -1 0 3030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1024_
timestamp 0
transform -1 0 2710 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1025_
timestamp 0
transform -1 0 4110 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1026_
timestamp 0
transform 1 0 3690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1027_
timestamp 0
transform 1 0 2950 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1028_
timestamp 0
transform 1 0 6310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1029_
timestamp 0
transform 1 0 4890 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1030_
timestamp 0
transform 1 0 3810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1032_
timestamp 0
transform 1 0 4610 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1033_
timestamp 0
transform 1 0 4110 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1034_
timestamp 0
transform 1 0 3910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1035_
timestamp 0
transform -1 0 4470 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1036_
timestamp 0
transform -1 0 4290 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1037_
timestamp 0
transform 1 0 6430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1038_
timestamp 0
transform 1 0 3970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1039_
timestamp 0
transform -1 0 4570 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1040_
timestamp 0
transform -1 0 4730 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1041_
timestamp 0
transform 1 0 4050 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1042_
timestamp 0
transform -1 0 4230 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1043_
timestamp 0
transform -1 0 4390 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1044_
timestamp 0
transform 1 0 3750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1045_
timestamp 0
transform -1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1046_
timestamp 0
transform -1 0 2650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1047_
timestamp 0
transform 1 0 4250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1048_
timestamp 0
transform -1 0 4090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1049_
timestamp 0
transform -1 0 3830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1050_
timestamp 0
transform 1 0 3330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1051_
timestamp 0
transform -1 0 3530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1052_
timestamp 0
transform -1 0 4630 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1053_
timestamp 0
transform -1 0 4110 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1054_
timestamp 0
transform 1 0 3750 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1055_
timestamp 0
transform -1 0 3890 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1056_
timestamp 0
transform -1 0 3950 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1057_
timestamp 0
transform 1 0 3750 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1058_
timestamp 0
transform -1 0 3590 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1059_
timestamp 0
transform -1 0 3110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1060_
timestamp 0
transform 1 0 3430 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1061_
timestamp 0
transform -1 0 3610 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1062_
timestamp 0
transform -1 0 3470 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1063_
timestamp 0
transform 1 0 570 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1064_
timestamp 0
transform 1 0 730 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1065_
timestamp 0
transform 1 0 1130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1066_
timestamp 0
transform 1 0 830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1067_
timestamp 0
transform -1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1068_
timestamp 0
transform -1 0 1090 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1069_
timestamp 0
transform -1 0 930 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1070_
timestamp 0
transform -1 0 1370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1071_
timestamp 0
transform 1 0 2450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1072_
timestamp 0
transform -1 0 3290 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1073_
timestamp 0
transform -1 0 3110 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1074_
timestamp 0
transform -1 0 2790 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1075_
timestamp 0
transform 1 0 1530 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1076_
timestamp 0
transform -1 0 1430 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1077_
timestamp 0
transform 1 0 1250 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1078_
timestamp 0
transform -1 0 3210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1080_
timestamp 0
transform 1 0 1870 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1081_
timestamp 0
transform -1 0 2730 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1082_
timestamp 0
transform 1 0 1910 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1083_
timestamp 0
transform -1 0 2390 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1084_
timestamp 0
transform 1 0 1530 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1085_
timestamp 0
transform -1 0 1570 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1086_
timestamp 0
transform 1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1087_
timestamp 0
transform -1 0 1570 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1088_
timestamp 0
transform -1 0 1250 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1089_
timestamp 0
transform 1 0 1370 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1090_
timestamp 0
transform -1 0 990 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1091_
timestamp 0
transform 1 0 450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1092_
timestamp 0
transform 1 0 90 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1093_
timestamp 0
transform -1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1094_
timestamp 0
transform 1 0 90 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1095_
timestamp 0
transform 1 0 950 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1096_
timestamp 0
transform -1 0 1230 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1097_
timestamp 0
transform 1 0 770 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1098_
timestamp 0
transform -1 0 110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1099_
timestamp 0
transform 1 0 90 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1100_
timestamp 0
transform -1 0 1950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1101_
timestamp 0
transform -1 0 2490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1102_
timestamp 0
transform 1 0 2090 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1103_
timestamp 0
transform -1 0 2310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1104_
timestamp 0
transform -1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1105_
timestamp 0
transform -1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1106_
timestamp 0
transform -1 0 910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1107_
timestamp 0
transform -1 0 1010 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1108_
timestamp 0
transform 1 0 1050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1109_
timestamp 0
transform -1 0 650 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1110_
timestamp 0
transform -1 0 750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1111_
timestamp 0
transform -1 0 750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1112_
timestamp 0
transform -1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1113_
timestamp 0
transform 1 0 570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1114_
timestamp 0
transform -1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1115_
timestamp 0
transform -1 0 270 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1116_
timestamp 0
transform 1 0 410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1117_
timestamp 0
transform 1 0 230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1118_
timestamp 0
transform 1 0 270 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1119_
timestamp 0
transform 1 0 2190 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1120_
timestamp 0
transform -1 0 2350 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1121_
timestamp 0
transform 1 0 2030 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1122_
timestamp 0
transform -1 0 2430 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1123_
timestamp 0
transform 1 0 2250 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1124_
timestamp 0
transform 1 0 1690 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1125_
timestamp 0
transform 1 0 1870 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1126_
timestamp 0
transform 1 0 1770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1128_
timestamp 0
transform 1 0 1530 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1129_
timestamp 0
transform 1 0 1570 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1130_
timestamp 0
transform -1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1131_
timestamp 0
transform -1 0 2090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1132_
timestamp 0
transform -1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1133_
timestamp 0
transform -1 0 1950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1134_
timestamp 0
transform -1 0 1750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1135_
timestamp 0
transform 1 0 1230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1136_
timestamp 0
transform -1 0 1410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1137_
timestamp 0
transform -1 0 1090 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1138_
timestamp 0
transform -1 0 630 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1139_
timestamp 0
transform -1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1140_
timestamp 0
transform -1 0 3910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1141_
timestamp 0
transform 1 0 4110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1142_
timestamp 0
transform -1 0 4650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1143_
timestamp 0
transform 1 0 5550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1144_
timestamp 0
transform 1 0 6570 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1145_
timestamp 0
transform -1 0 5550 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1146_
timestamp 0
transform 1 0 4830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1147_
timestamp 0
transform -1 0 5030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1148_
timestamp 0
transform -1 0 4670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1149_
timestamp 0
transform 1 0 5710 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1150_
timestamp 0
transform -1 0 5230 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1151_
timestamp 0
transform -1 0 5210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1152_
timestamp 0
transform -1 0 4490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1153_
timestamp 0
transform -1 0 4330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1154_
timestamp 0
transform -1 0 6390 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1155_
timestamp 0
transform -1 0 6810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1156_
timestamp 0
transform 1 0 3250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1157_
timestamp 0
transform 1 0 3570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1158_
timestamp 0
transform -1 0 6170 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1159_
timestamp 0
transform 1 0 5370 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1160_
timestamp 0
transform 1 0 5290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1161_
timestamp 0
transform 1 0 4230 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1162_
timestamp 0
transform -1 0 5090 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1163_
timestamp 0
transform 1 0 4870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1164_
timestamp 0
transform 1 0 5110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1165_
timestamp 0
transform 1 0 5130 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1166_
timestamp 0
transform -1 0 4890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1167_
timestamp 0
transform -1 0 5990 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1168_
timestamp 0
transform 1 0 5850 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1169_
timestamp 0
transform 1 0 3890 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1170_
timestamp 0
transform 1 0 3170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1171_
timestamp 0
transform 1 0 2930 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1172_
timestamp 0
transform -1 0 3110 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1173_
timestamp 0
transform 1 0 3070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1174_
timestamp 0
transform 1 0 3570 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1176_
timestamp 0
transform -1 0 4070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1177_
timestamp 0
transform 1 0 4390 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1178_
timestamp 0
transform -1 0 5070 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1179_
timestamp 0
transform 1 0 5370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1180_
timestamp 0
transform 1 0 4770 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1181_
timestamp 0
transform 1 0 5310 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1182_
timestamp 0
transform 1 0 5210 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1183_
timestamp 0
transform -1 0 5430 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1184_
timestamp 0
transform 1 0 5210 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1185_
timestamp 0
transform -1 0 4590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1186_
timestamp 0
transform -1 0 5610 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1187_
timestamp 0
transform -1 0 5190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1188_
timestamp 0
transform -1 0 4850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1189_
timestamp 0
transform -1 0 4550 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1190_
timestamp 0
transform 1 0 5730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1191_
timestamp 0
transform 1 0 6190 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1192_
timestamp 0
transform 1 0 4310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1193_
timestamp 0
transform -1 0 4370 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1194_
timestamp 0
transform -1 0 3690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1195_
timestamp 0
transform 1 0 3710 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1196_
timestamp 0
transform 1 0 3530 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1197_
timestamp 0
transform 1 0 3170 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1198_
timestamp 0
transform 1 0 3430 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1199_
timestamp 0
transform -1 0 3430 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1200_
timestamp 0
transform -1 0 2250 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1201_
timestamp 0
transform 1 0 3590 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1202_
timestamp 0
transform 1 0 3410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1203_
timestamp 0
transform -1 0 3270 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1204_
timestamp 0
transform 1 0 2570 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1205_
timestamp 0
transform 1 0 2470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1206_
timestamp 0
transform 1 0 2150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1207_
timestamp 0
transform 1 0 2770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1208_
timestamp 0
transform 1 0 2290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1209_
timestamp 0
transform -1 0 3130 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1210_
timestamp 0
transform -1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1211_
timestamp 0
transform 1 0 2750 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1212_
timestamp 0
transform 1 0 4510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1213_
timestamp 0
transform 1 0 4670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1214_
timestamp 0
transform 1 0 4150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1215_
timestamp 0
transform -1 0 4050 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1216_
timestamp 0
transform 1 0 4730 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1217_
timestamp 0
transform 1 0 4190 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1218_
timestamp 0
transform -1 0 3890 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1219_
timestamp 0
transform -1 0 3190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1220_
timestamp 0
transform 1 0 3810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1221_
timestamp 0
transform -1 0 3390 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1222_
timestamp 0
transform 1 0 3370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1224_
timestamp 0
transform 1 0 3630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1225_
timestamp 0
transform -1 0 3730 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1226_
timestamp 0
transform -1 0 3990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1227_
timestamp 0
transform 1 0 3330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1228_
timestamp 0
transform -1 0 3390 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1229_
timestamp 0
transform -1 0 3550 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1230_
timestamp 0
transform 1 0 2830 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1231_
timestamp 0
transform 1 0 2410 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1232_
timestamp 0
transform 1 0 1990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1233_
timestamp 0
transform -1 0 1910 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1234_
timestamp 0
transform -1 0 2250 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1235_
timestamp 0
transform 1 0 2510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1236_
timestamp 0
transform -1 0 2710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1237_
timestamp 0
transform 1 0 2870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1238_
timestamp 0
transform -1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1239_
timestamp 0
transform -1 0 1850 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1240_
timestamp 0
transform 1 0 1910 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1241_
timestamp 0
transform -1 0 2430 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1242_
timestamp 0
transform -1 0 2030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1243_
timestamp 0
transform 1 0 2190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1244_
timestamp 0
transform 1 0 1330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1245_
timestamp 0
transform -1 0 1690 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1246_
timestamp 0
transform 1 0 1650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1247_
timestamp 0
transform -1 0 2770 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1248_
timestamp 0
transform 1 0 2570 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1249_
timestamp 0
transform -1 0 1550 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1250_
timestamp 0
transform -1 0 1490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1251_
timestamp 0
transform 1 0 1730 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1252_
timestamp 0
transform -1 0 2070 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1253_
timestamp 0
transform -1 0 2110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1254_
timestamp 0
transform 1 0 1830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1255_
timestamp 0
transform 1 0 1910 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1256_
timestamp 0
transform -1 0 1730 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1257_
timestamp 0
transform 1 0 2270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1258_
timestamp 0
transform 1 0 2110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1259_
timestamp 0
transform 1 0 1870 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1260_
timestamp 0
transform -1 0 1490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1261_
timestamp 0
transform -1 0 1410 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1262_
timestamp 0
transform 1 0 2010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1263_
timestamp 0
transform -1 0 2250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1264_
timestamp 0
transform -1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1265_
timestamp 0
transform -1 0 1930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1266_
timestamp 0
transform 1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1267_
timestamp 0
transform 1 0 2050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1268_
timestamp 0
transform -1 0 2270 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1269_
timestamp 0
transform 1 0 2230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1270_
timestamp 0
transform -1 0 2410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1272_
timestamp 0
transform 1 0 2050 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1273_
timestamp 0
transform -1 0 2650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1274_
timestamp 0
transform -1 0 310 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1275_
timestamp 0
transform -1 0 470 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1276_
timestamp 0
transform 1 0 90 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1277_
timestamp 0
transform 1 0 430 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1278_
timestamp 0
transform -1 0 810 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1279_
timestamp 0
transform 1 0 430 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1280_
timestamp 0
transform 1 0 250 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1281_
timestamp 0
transform -1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1282_
timestamp 0
transform -1 0 770 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1283_
timestamp 0
transform 1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1284_
timestamp 0
transform 1 0 1570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1285_
timestamp 0
transform -1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1286_
timestamp 0
transform -1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1287_
timestamp 0
transform -1 0 1350 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1288_
timestamp 0
transform 1 0 1930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1289_
timestamp 0
transform -1 0 1150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1290_
timestamp 0
transform -1 0 1170 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1291_
timestamp 0
transform 1 0 570 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1292_
timestamp 0
transform -1 0 110 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1293_
timestamp 0
transform -1 0 110 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1294_
timestamp 0
transform -1 0 270 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1295_
timestamp 0
transform 1 0 590 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1296_
timestamp 0
transform -1 0 830 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1297_
timestamp 0
transform 1 0 1770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1298_
timestamp 0
transform -1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1299_
timestamp 0
transform -1 0 1010 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1300_
timestamp 0
transform -1 0 1690 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1301_
timestamp 0
transform 1 0 2170 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1302_
timestamp 0
transform 1 0 1990 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1303_
timestamp 0
transform 1 0 2210 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1304_
timestamp 0
transform -1 0 2610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1305_
timestamp 0
transform -1 0 1570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1306_
timestamp 0
transform -1 0 1410 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1307_
timestamp 0
transform 1 0 1390 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1308_
timestamp 0
transform 1 0 1370 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1309_
timestamp 0
transform -1 0 5270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1310_
timestamp 0
transform 1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1311_
timestamp 0
transform 1 0 2610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1312_
timestamp 0
transform 1 0 1690 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1313_
timestamp 0
transform 1 0 1730 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1314_
timestamp 0
transform 1 0 2790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1315_
timestamp 0
transform -1 0 5010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1316_
timestamp 0
transform 1 0 5670 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1317_
timestamp 0
transform 1 0 5550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1318_
timestamp 0
transform 1 0 5830 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1320_
timestamp 0
transform -1 0 6410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1321_
timestamp 0
transform -1 0 6710 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1322_
timestamp 0
transform -1 0 6770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1323_
timestamp 0
transform 1 0 6770 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1324_
timestamp 0
transform 1 0 5030 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1325_
timestamp 0
transform -1 0 5510 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1326_
timestamp 0
transform 1 0 5350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1327_
timestamp 0
transform 1 0 5550 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1328_
timestamp 0
transform 1 0 5730 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1329_
timestamp 0
transform 1 0 5910 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1330_
timestamp 0
transform 1 0 5450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1331_
timestamp 0
transform 1 0 6450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1332_
timestamp 0
transform -1 0 5810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1333_
timestamp 0
transform 1 0 5950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1334_
timestamp 0
transform -1 0 6190 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1335_
timestamp 0
transform 1 0 6410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1336_
timestamp 0
transform 1 0 6570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1337_
timestamp 0
transform -1 0 6750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1338_
timestamp 0
transform -1 0 6750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1339_
timestamp 0
transform -1 0 6850 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1340_
timestamp 0
transform 1 0 6510 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1341_
timestamp 0
transform -1 0 6870 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1342_
timestamp 0
transform 1 0 5630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1343_
timestamp 0
transform 1 0 6590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1344_
timestamp 0
transform -1 0 6770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1345_
timestamp 0
transform 1 0 6650 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1346_
timestamp 0
transform 1 0 6590 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1347_
timestamp 0
transform 1 0 5850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1348_
timestamp 0
transform 1 0 6350 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1349_
timestamp 0
transform -1 0 6590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1350_
timestamp 0
transform 1 0 6530 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1351_
timestamp 0
transform 1 0 5530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1352_
timestamp 0
transform 1 0 5750 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1353_
timestamp 0
transform -1 0 5930 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1354_
timestamp 0
transform 1 0 6090 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1355_
timestamp 0
transform 1 0 6390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1356_
timestamp 0
transform 1 0 6570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1357_
timestamp 0
transform -1 0 6230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1358_
timestamp 0
transform 1 0 6030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4__1359_
timestamp 0
transform 1 0 6490 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1360_
timestamp 0
transform 1 0 6110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1361_
timestamp 0
transform -1 0 6290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1362_
timestamp 0
transform -1 0 6730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1363_
timestamp 0
transform 1 0 6670 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1364_
timestamp 0
transform -1 0 6750 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1365_
timestamp 0
transform -1 0 6850 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1366_
timestamp 0
transform -1 0 6090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1368_
timestamp 0
transform -1 0 5370 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1369_
timestamp 0
transform -1 0 4570 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1370_
timestamp 0
transform 1 0 3890 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1371_
timestamp 0
transform 1 0 4230 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1372_
timestamp 0
transform -1 0 5130 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1373_
timestamp 0
transform -1 0 4710 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1374_
timestamp 0
transform 1 0 5830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1375_
timestamp 0
transform -1 0 5390 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1376_
timestamp 0
transform 1 0 6550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1377_
timestamp 0
transform -1 0 6870 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1378_
timestamp 0
transform -1 0 6630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1379_
timestamp 0
transform -1 0 6690 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1380_
timestamp 0
transform 1 0 6190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1381_
timestamp 0
transform -1 0 6390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1382_
timestamp 0
transform -1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1383_
timestamp 0
transform 1 0 4810 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1384_
timestamp 0
transform -1 0 4990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1385_
timestamp 0
transform -1 0 5230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1386_
timestamp 0
transform -1 0 5030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1387_
timestamp 0
transform -1 0 5030 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1388_
timestamp 0
transform 1 0 4310 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1389_
timestamp 0
transform -1 0 4530 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1390_
timestamp 0
transform -1 0 1930 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1391_
timestamp 0
transform -1 0 1390 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1392_
timestamp 0
transform -1 0 1410 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1393_
timestamp 0
transform -1 0 910 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1394_
timestamp 0
transform 1 0 970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1395_
timestamp 0
transform -1 0 4150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1396_
timestamp 0
transform -1 0 3030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1397_
timestamp 0
transform 1 0 2830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1398_
timestamp 0
transform 1 0 4370 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1399_
timestamp 0
transform 1 0 4510 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1400_
timestamp 0
transform 1 0 6010 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1401_
timestamp 0
transform -1 0 5930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1402_
timestamp 0
transform -1 0 4470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1403_
timestamp 0
transform 1 0 4770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1404_
timestamp 0
transform 1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1405_
timestamp 0
transform 1 0 4910 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1406_
timestamp 0
transform -1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1407_
timestamp 0
transform -1 0 5150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1408_
timestamp 0
transform 1 0 5070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1409_
timestamp 0
transform -1 0 5090 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1410_
timestamp 0
transform 1 0 4350 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1411_
timestamp 0
transform -1 0 6110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1412_
timestamp 0
transform 1 0 5370 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1413_
timestamp 0
transform 1 0 6250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1414_
timestamp 0
transform -1 0 6590 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1416_
timestamp 0
transform -1 0 6430 0 1 5990
box -6 -8 26 268
use FILL  FILL_4__1417_
timestamp 0
transform -1 0 5510 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1418_
timestamp 0
transform -1 0 5050 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1419_
timestamp 0
transform -1 0 4430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1420_
timestamp 0
transform -1 0 4810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1421_
timestamp 0
transform -1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1422_
timestamp 0
transform 1 0 4410 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1423_
timestamp 0
transform -1 0 4630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1424_
timestamp 0
transform 1 0 4030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1425_
timestamp 0
transform -1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1426_
timestamp 0
transform 1 0 790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1427_
timestamp 0
transform 1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1428_
timestamp 0
transform 1 0 2390 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1429_
timestamp 0
transform -1 0 4070 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1430_
timestamp 0
transform -1 0 4730 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1431_
timestamp 0
transform -1 0 4910 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1432_
timestamp 0
transform -1 0 4730 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1433_
timestamp 0
transform -1 0 4910 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1434_
timestamp 0
transform 1 0 2410 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1435_
timestamp 0
transform 1 0 4710 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1436_
timestamp 0
transform -1 0 2290 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1437_
timestamp 0
transform 1 0 2370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1438_
timestamp 0
transform 1 0 2430 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1439_
timestamp 0
transform 1 0 2690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1440_
timestamp 0
transform 1 0 3010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1441_
timestamp 0
transform -1 0 2870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1442_
timestamp 0
transform 1 0 2770 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1443_
timestamp 0
transform 1 0 2230 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1444_
timestamp 0
transform 1 0 1710 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1445_
timestamp 0
transform 1 0 1750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1446_
timestamp 0
transform 1 0 2410 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1447_
timestamp 0
transform 1 0 2530 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1448_
timestamp 0
transform 1 0 2910 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1449_
timestamp 0
transform 1 0 4390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1450_
timestamp 0
transform -1 0 4230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1451_
timestamp 0
transform 1 0 4850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1452_
timestamp 0
transform 1 0 2850 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1453_
timestamp 0
transform 1 0 2670 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1454_
timestamp 0
transform -1 0 2850 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1455_
timestamp 0
transform -1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1456_
timestamp 0
transform 1 0 5290 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1457_
timestamp 0
transform -1 0 5450 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1458_
timestamp 0
transform -1 0 5470 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1459_
timestamp 0
transform 1 0 3690 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1460_
timestamp 0
transform 1 0 4450 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1461_
timestamp 0
transform 1 0 3510 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1463_
timestamp 0
transform 1 0 2810 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1464_
timestamp 0
transform 1 0 2250 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1465_
timestamp 0
transform 1 0 2550 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1466_
timestamp 0
transform -1 0 2730 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1467_
timestamp 0
transform 1 0 3030 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1468_
timestamp 0
transform 1 0 3170 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1469_
timestamp 0
transform 1 0 2630 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1470_
timestamp 0
transform 1 0 3630 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1471_
timestamp 0
transform -1 0 3870 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1472_
timestamp 0
transform -1 0 3830 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1473_
timestamp 0
transform 1 0 4070 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1474_
timestamp 0
transform 1 0 5170 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1475_
timestamp 0
transform -1 0 4270 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1476_
timestamp 0
transform -1 0 4850 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1477_
timestamp 0
transform 1 0 4570 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1478_
timestamp 0
transform -1 0 4670 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1479_
timestamp 0
transform -1 0 4430 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1480_
timestamp 0
transform 1 0 6010 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1481_
timestamp 0
transform 1 0 5850 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1482_
timestamp 0
transform -1 0 5650 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1483_
timestamp 0
transform 1 0 3630 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1484_
timestamp 0
transform -1 0 2890 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1485_
timestamp 0
transform 1 0 3050 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1486_
timestamp 0
transform 1 0 3490 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1487_
timestamp 0
transform 1 0 3330 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1488_
timestamp 0
transform 1 0 3010 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1489_
timestamp 0
transform 1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1490_
timestamp 0
transform -1 0 3310 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1491_
timestamp 0
transform -1 0 4730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1492_
timestamp 0
transform -1 0 4630 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1493_
timestamp 0
transform -1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1494_
timestamp 0
transform 1 0 3550 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1495_
timestamp 0
transform 1 0 3730 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1496_
timestamp 0
transform -1 0 4470 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1497_
timestamp 0
transform 1 0 4990 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1498_
timestamp 0
transform 1 0 4490 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1499_
timestamp 0
transform 1 0 4310 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1500_
timestamp 0
transform -1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1501_
timestamp 0
transform 1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1502_
timestamp 0
transform 1 0 4230 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1503_
timestamp 0
transform 1 0 4230 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1504_
timestamp 0
transform -1 0 4550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1505_
timestamp 0
transform -1 0 4190 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1506_
timestamp 0
transform 1 0 4390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1507_
timestamp 0
transform 1 0 4630 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1508_
timestamp 0
transform 1 0 4830 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1509_
timestamp 0
transform 1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1511_
timestamp 0
transform 1 0 2410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1512_
timestamp 0
transform 1 0 2530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4__1513_
timestamp 0
transform -1 0 2610 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1514_
timestamp 0
transform -1 0 2610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1515_
timestamp 0
transform 1 0 2710 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1516_
timestamp 0
transform -1 0 2890 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1517_
timestamp 0
transform 1 0 3770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1518_
timestamp 0
transform 1 0 4050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1519_
timestamp 0
transform -1 0 4230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1520_
timestamp 0
transform 1 0 3210 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1521_
timestamp 0
transform -1 0 4030 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1522_
timestamp 0
transform -1 0 3890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1523_
timestamp 0
transform 1 0 3030 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1524_
timestamp 0
transform -1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1525_
timestamp 0
transform 1 0 3210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1526_
timestamp 0
transform 1 0 3370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1527_
timestamp 0
transform 1 0 3010 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1528_
timestamp 0
transform -1 0 3050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_4__1529_
timestamp 0
transform -1 0 1290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1530_
timestamp 0
transform 1 0 1430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1531_
timestamp 0
transform 1 0 1570 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1532_
timestamp 0
transform -1 0 1930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1533_
timestamp 0
transform -1 0 2090 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1534_
timestamp 0
transform -1 0 2390 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1535_
timestamp 0
transform -1 0 2770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1536_
timestamp 0
transform -1 0 3390 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1537_
timestamp 0
transform 1 0 2510 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1538_
timestamp 0
transform 1 0 3910 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1539_
timestamp 0
transform -1 0 3290 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1540_
timestamp 0
transform 1 0 1850 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1541_
timestamp 0
transform -1 0 3470 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1542_
timestamp 0
transform 1 0 2050 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1543_
timestamp 0
transform 1 0 3910 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1544_
timestamp 0
transform 1 0 3170 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1545_
timestamp 0
transform 1 0 2470 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1546_
timestamp 0
transform 1 0 3610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1547_
timestamp 0
transform 1 0 4770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1548_
timestamp 0
transform 1 0 3910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1549_
timestamp 0
transform -1 0 4910 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1550_
timestamp 0
transform 1 0 5030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1551_
timestamp 0
transform -1 0 5230 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1552_
timestamp 0
transform 1 0 4470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1553_
timestamp 0
transform -1 0 4550 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1554_
timestamp 0
transform 1 0 5250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1555_
timestamp 0
transform 1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1556_
timestamp 0
transform -1 0 5070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1557_
timestamp 0
transform -1 0 4870 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1559_
timestamp 0
transform 1 0 4990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1560_
timestamp 0
transform -1 0 5030 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1561_
timestamp 0
transform -1 0 4670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1562_
timestamp 0
transform 1 0 3990 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1563_
timestamp 0
transform -1 0 4190 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1564_
timestamp 0
transform -1 0 4890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1565_
timestamp 0
transform 1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1566_
timestamp 0
transform 1 0 3510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1567_
timestamp 0
transform -1 0 3030 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1568_
timestamp 0
transform 1 0 3670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1569_
timestamp 0
transform -1 0 3330 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1570_
timestamp 0
transform 1 0 3150 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1571_
timestamp 0
transform 1 0 3210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1572_
timestamp 0
transform 1 0 3390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1573_
timestamp 0
transform 1 0 3950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1574_
timestamp 0
transform -1 0 4490 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1575_
timestamp 0
transform -1 0 3990 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1576_
timestamp 0
transform -1 0 4150 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1577_
timestamp 0
transform -1 0 3470 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1578_
timestamp 0
transform -1 0 3830 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1579_
timestamp 0
transform 1 0 3630 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1580_
timestamp 0
transform 1 0 3710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1581_
timestamp 0
transform -1 0 3910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1582_
timestamp 0
transform 1 0 4350 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1583_
timestamp 0
transform -1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1584_
timestamp 0
transform -1 0 4650 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1585_
timestamp 0
transform 1 0 4250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1586_
timestamp 0
transform -1 0 4730 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1587_
timestamp 0
transform -1 0 3310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1588_
timestamp 0
transform -1 0 3170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1589_
timestamp 0
transform -1 0 4470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1590_
timestamp 0
transform -1 0 4330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1591_
timestamp 0
transform 1 0 4290 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1592_
timestamp 0
transform 1 0 4130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1593_
timestamp 0
transform 1 0 2650 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1594_
timestamp 0
transform 1 0 2830 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1595_
timestamp 0
transform -1 0 3030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1596_
timestamp 0
transform -1 0 3230 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1597_
timestamp 0
transform 1 0 3030 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1598_
timestamp 0
transform -1 0 3390 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1599_
timestamp 0
transform -1 0 3730 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1600_
timestamp 0
transform 1 0 3530 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1601_
timestamp 0
transform -1 0 3470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1602_
timestamp 0
transform -1 0 2930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1603_
timestamp 0
transform -1 0 3110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1604_
timestamp 0
transform -1 0 3290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1605_
timestamp 0
transform 1 0 4130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1607_
timestamp 0
transform 1 0 6290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1608_
timestamp 0
transform -1 0 6470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1609_
timestamp 0
transform 1 0 6230 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1610_
timestamp 0
transform 1 0 6630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1611_
timestamp 0
transform 1 0 5670 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1612_
timestamp 0
transform -1 0 6890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_4__1613_
timestamp 0
transform -1 0 6510 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1614_
timestamp 0
transform -1 0 6330 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1615_
timestamp 0
transform -1 0 6150 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1616_
timestamp 0
transform 1 0 5950 0 1 3390
box -6 -8 26 268
use FILL  FILL_4__1617_
timestamp 0
transform 1 0 5690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4__1618_
timestamp 0
transform -1 0 5490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1619_
timestamp 0
transform 1 0 5390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1620_
timestamp 0
transform -1 0 6170 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1621_
timestamp 0
transform 1 0 5390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1622_
timestamp 0
transform 1 0 6810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1623_
timestamp 0
transform 1 0 6470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1624_
timestamp 0
transform -1 0 6870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1625_
timestamp 0
transform -1 0 6610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1626_
timestamp 0
transform 1 0 6590 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1627_
timestamp 0
transform 1 0 6430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1628_
timestamp 0
transform -1 0 6230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1629_
timestamp 0
transform 1 0 6010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1630_
timestamp 0
transform 1 0 6730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_4__1631_
timestamp 0
transform -1 0 6790 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1632_
timestamp 0
transform -1 0 6670 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1633_
timestamp 0
transform -1 0 6690 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1634_
timestamp 0
transform -1 0 6510 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1635_
timestamp 0
transform 1 0 6310 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1636_
timestamp 0
transform -1 0 6490 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1637_
timestamp 0
transform 1 0 6130 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1638_
timestamp 0
transform -1 0 6530 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1639_
timestamp 0
transform 1 0 6390 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1640_
timestamp 0
transform 1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1641_
timestamp 0
transform -1 0 6790 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1642_
timestamp 0
transform -1 0 6290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1643_
timestamp 0
transform -1 0 6590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1644_
timestamp 0
transform -1 0 6290 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1645_
timestamp 0
transform 1 0 6610 0 -1 790
box -6 -8 26 268
use FILL  FILL_4__1646_
timestamp 0
transform -1 0 6750 0 1 790
box -6 -8 26 268
use FILL  FILL_4__1647_
timestamp 0
transform -1 0 6070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1648_
timestamp 0
transform 1 0 5850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1649_
timestamp 0
transform -1 0 6750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1650_
timestamp 0
transform -1 0 6750 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1651_
timestamp 0
transform -1 0 6310 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1652_
timestamp 0
transform -1 0 6530 0 1 2870
box -6 -8 26 268
use FILL  FILL_4__1653_
timestamp 0
transform 1 0 5650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1655_
timestamp 0
transform 1 0 6410 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1656_
timestamp 0
transform 1 0 6590 0 1 2350
box -6 -8 26 268
use FILL  FILL_4__1657_
timestamp 0
transform -1 0 6850 0 1 270
box -6 -8 26 268
use FILL  FILL_4__1658_
timestamp 0
transform 1 0 6190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1659_
timestamp 0
transform -1 0 6890 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1660_
timestamp 0
transform -1 0 6670 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1661_
timestamp 0
transform -1 0 6850 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1662_
timestamp 0
transform -1 0 6490 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1663_
timestamp 0
transform 1 0 6070 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1664_
timestamp 0
transform 1 0 6250 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1665_
timestamp 0
transform -1 0 6370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1666_
timestamp 0
transform -1 0 6690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1667_
timestamp 0
transform 1 0 6450 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1668_
timestamp 0
transform 1 0 6750 0 1 1310
box -6 -8 26 268
use FILL  FILL_4__1669_
timestamp 0
transform -1 0 6030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1670_
timestamp 0
transform 1 0 5890 0 1 1830
box -6 -8 26 268
use FILL  FILL_4__1671_
timestamp 0
transform 1 0 5570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1672_
timestamp 0
transform -1 0 6130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1673_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1674_
timestamp 0
transform -1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1675_
timestamp 0
transform 1 0 4050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_4__1676_
timestamp 0
transform 1 0 5230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4__1677_
timestamp 0
transform 1 0 5150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_4__1711_
timestamp 0
transform -1 0 110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4__1712_
timestamp 0
transform -1 0 110 0 1 4950
box -6 -8 26 268
use FILL  FILL_4__1713_
timestamp 0
transform -1 0 1110 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1714_
timestamp 0
transform 1 0 250 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1715_
timestamp 0
transform -1 0 110 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1716_
timestamp 0
transform -1 0 110 0 1 4430
box -6 -8 26 268
use FILL  FILL_4__1717_
timestamp 0
transform 1 0 410 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1718_
timestamp 0
transform -1 0 110 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1719_
timestamp 0
transform 1 0 1250 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1720_
timestamp 0
transform -1 0 110 0 1 5470
box -6 -8 26 268
use FILL  FILL_4__1721_
timestamp 0
transform -1 0 270 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1722_
timestamp 0
transform -1 0 110 0 1 3910
box -6 -8 26 268
use FILL  FILL_4__1723_
timestamp 0
transform 1 0 1550 0 -1 270
box -6 -8 26 268
use FILL  FILL_4__1724_
timestamp 0
transform 1 0 410 0 -1 6510
box -6 -8 26 268
use FILL  FILL_4__1725_
timestamp 0
transform -1 0 470 0 1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert0
timestamp 0
transform -1 0 110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert1
timestamp 0
transform 1 0 290 0 1 5990
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert2
timestamp 0
transform 1 0 250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert3
timestamp 0
transform 1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert11
timestamp 0
transform 1 0 5850 0 -1 270
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert12
timestamp 0
transform -1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform 1 0 5670 0 1 2870
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform -1 0 2530 0 1 790
box -6 -8 26 268
use FILL  FILL_4_BUFX2_insert15
timestamp 0
transform 1 0 3390 0 1 1310
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert4
timestamp 0
transform 1 0 5010 0 1 790
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert5
timestamp 0
transform -1 0 1970 0 1 4950
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert6
timestamp 0
transform -1 0 4830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert7
timestamp 0
transform 1 0 550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert8
timestamp 0
transform -1 0 450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert9
timestamp 0
transform 1 0 2630 0 1 1830
box -6 -8 26 268
use FILL  FILL_4_CLKBUF1_insert10
timestamp 0
transform -1 0 3610 0 -1 1310
box -6 -8 26 268
<< labels >>
flabel metal1 s 6963 2 7023 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 4296 -16 4304 7 FreeSans 16 0 0 0 clk
port 2 nsew
flabel metal3 s 6996 3516 7004 3524 3 FreeSans 16 0 0 0 down
port 3 nsew
flabel metal3 s -24 4816 -16 4824 7 FreeSans 16 0 0 0 hsync
port 4 nsew
flabel metal3 s -24 5076 -16 5084 7 FreeSans 16 0 0 0 p_tick
port 5 nsew
flabel metal3 s -24 6116 -16 6124 7 FreeSans 16 0 0 0 reset
port 6 nsew
flabel metal3 s -24 4556 -16 4564 7 FreeSans 16 0 0 0 rgb[11]
port 7 nsew
flabel metal3 s -24 136 -16 144 7 FreeSans 16 0 0 0 rgb[10]
port 8 nsew
flabel metal2 s 477 6557 483 6563 3 FreeSans 16 90 0 0 rgb[9]
port 9 nsew
flabel metal2 s 1597 -23 1603 -17 7 FreeSans 16 270 0 0 rgb[8]
port 10 nsew
flabel metal3 s -24 4036 -16 4044 7 FreeSans 16 0 0 0 rgb[7]
port 11 nsew
flabel metal2 s 297 -23 303 -17 7 FreeSans 16 270 0 0 rgb[6]
port 12 nsew
flabel metal3 s -24 5596 -16 5604 7 FreeSans 16 0 0 0 rgb[5]
port 13 nsew
flabel metal2 s 1297 -23 1303 -17 7 FreeSans 16 270 0 0 rgb[4]
port 14 nsew
flabel metal3 s -24 6376 -16 6384 7 FreeSans 16 0 0 0 rgb[3]
port 15 nsew
flabel metal2 s 457 -23 463 -17 7 FreeSans 16 270 0 0 rgb[2]
port 16 nsew
flabel metal2 s 297 6557 303 6563 3 FreeSans 16 90 0 0 rgb[1]
port 17 nsew
flabel metal2 s 1137 -23 1143 -17 7 FreeSans 16 270 0 0 rgb[0]
port 18 nsew
flabel metal3 s 6996 2216 7004 2224 3 FreeSans 16 0 0 0 up
port 19 nsew
flabel metal2 s 437 6557 443 6563 3 FreeSans 16 90 0 0 vsync
port 20 nsew
<< properties >>
string FIXED_BBOX -40 -40 7000 6560
<< end >>
