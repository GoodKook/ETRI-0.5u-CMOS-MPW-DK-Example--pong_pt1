VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pong_pt1
  CLASS BLOCK ;
  FOREIGN pong_pt1 ;
  ORIGIN 6.000 6.000 ;
  SIZE 1056.000 BY 990.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 975.300 1053.450 977.700 ;
        RECT 1044.450 899.700 1053.450 975.300 ;
        RECT 0.600 897.300 1053.450 899.700 ;
        RECT 1044.450 821.700 1053.450 897.300 ;
        RECT 0.600 819.300 1053.450 821.700 ;
        RECT 1044.450 743.700 1053.450 819.300 ;
        RECT 0.600 741.300 1053.450 743.700 ;
        RECT 1044.450 665.700 1053.450 741.300 ;
        RECT 0.600 663.300 1053.450 665.700 ;
        RECT 1044.450 587.700 1053.450 663.300 ;
        RECT 0.600 585.300 1053.450 587.700 ;
        RECT 1044.450 509.700 1053.450 585.300 ;
        RECT 0.600 507.300 1053.450 509.700 ;
        RECT 1044.450 431.700 1053.450 507.300 ;
        RECT 0.600 429.300 1053.450 431.700 ;
        RECT 1044.450 353.700 1053.450 429.300 ;
        RECT 0.600 351.300 1053.450 353.700 ;
        RECT 1044.450 275.700 1053.450 351.300 ;
        RECT 0.600 273.300 1053.450 275.700 ;
        RECT 1044.450 197.700 1053.450 273.300 ;
        RECT 0.600 195.300 1053.450 197.700 ;
        RECT 1044.450 119.700 1053.450 195.300 ;
        RECT 0.600 117.300 1053.450 119.700 ;
        RECT 1044.450 41.700 1053.450 117.300 ;
        RECT 0.600 39.300 1053.450 41.700 ;
        RECT 1044.450 0.300 1053.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 938.700 -0.450 977.700 ;
        RECT -9.450 936.300 1043.400 938.700 ;
        RECT -9.450 860.700 -0.450 936.300 ;
        RECT 34.950 933.450 37.050 934.050 ;
        RECT 41.550 933.450 42.450 936.300 ;
        RECT 79.950 934.950 82.050 936.300 ;
        RECT 142.950 934.950 145.050 936.300 ;
        RECT 226.950 934.950 229.050 936.300 ;
        RECT 292.950 934.950 295.050 936.300 ;
        RECT 34.950 932.550 42.450 933.450 ;
        RECT 34.950 931.950 37.050 932.550 ;
        RECT -9.450 858.300 1043.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT 172.950 856.950 175.050 858.300 ;
        RECT 178.950 856.950 181.050 858.300 ;
        RECT 150.000 840.450 154.050 841.050 ;
        RECT 149.550 838.950 154.050 840.450 ;
        RECT 149.550 835.050 150.450 838.950 ;
        RECT 149.550 833.550 154.050 835.050 ;
        RECT 150.000 832.950 154.050 833.550 ;
        RECT -9.450 780.300 1043.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 13.950 778.950 16.050 780.300 ;
        RECT 37.950 778.950 40.050 780.300 ;
        RECT 178.950 778.950 181.050 780.300 ;
        RECT -9.450 702.300 1043.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT -9.450 624.300 1043.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 121.950 622.950 124.050 624.300 ;
        RECT -9.450 546.300 1043.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 97.950 544.950 100.050 546.300 ;
        RECT 178.950 544.950 181.050 546.300 ;
        RECT 607.950 544.950 610.050 546.300 ;
        RECT 643.950 544.950 646.050 546.300 ;
        RECT 721.950 544.950 724.050 546.300 ;
        RECT 883.950 544.950 886.050 546.300 ;
        RECT -9.450 468.300 1043.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 595.950 466.950 598.050 468.300 ;
        RECT 790.950 466.950 793.050 468.300 ;
        RECT 871.950 426.450 874.050 427.050 ;
        RECT 877.950 426.450 880.050 427.050 ;
        RECT 871.950 425.550 880.050 426.450 ;
        RECT 871.950 424.950 874.050 425.550 ;
        RECT 877.950 424.950 880.050 425.550 ;
        RECT -9.450 390.300 1043.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 52.950 388.950 55.050 390.300 ;
        RECT 100.950 388.950 103.050 390.300 ;
        RECT 901.950 387.450 904.050 388.050 ;
        RECT 911.550 387.450 912.450 390.300 ;
        RECT 901.950 386.550 912.450 387.450 ;
        RECT 901.950 385.950 904.050 386.550 ;
        RECT -9.450 312.300 1043.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 13.950 310.950 16.050 312.300 ;
        RECT 385.950 310.950 388.050 312.300 ;
        RECT 424.950 310.950 427.050 312.300 ;
        RECT 433.950 310.950 436.050 312.300 ;
        RECT 586.950 310.950 589.050 312.300 ;
        RECT 872.550 306.450 873.450 312.300 ;
        RECT 880.950 306.450 883.050 307.050 ;
        RECT 872.550 305.550 883.050 306.450 ;
        RECT 880.950 304.950 883.050 305.550 ;
        RECT -9.450 234.300 1043.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 442.950 232.950 445.050 234.300 ;
        RECT 445.950 232.950 448.050 234.300 ;
        RECT 472.950 232.950 475.050 234.300 ;
        RECT 502.950 232.950 505.050 234.300 ;
        RECT 733.950 232.950 736.050 234.300 ;
        RECT 838.950 232.950 841.050 234.300 ;
        RECT 847.950 232.950 850.050 234.300 ;
        RECT -9.450 156.300 1043.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 352.950 154.950 355.050 156.300 ;
        RECT 466.950 154.950 469.050 156.300 ;
        RECT 835.950 154.950 838.050 156.300 ;
        RECT 874.950 154.950 877.050 156.300 ;
        RECT 913.950 154.950 916.050 156.300 ;
        RECT -9.450 78.300 1043.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT 301.950 76.950 304.050 78.300 ;
        RECT 328.950 76.950 331.050 78.300 ;
        RECT 760.950 76.950 763.050 78.300 ;
        RECT 967.950 76.950 970.050 78.300 ;
        RECT 322.950 51.450 325.050 51.750 ;
        RECT 328.950 51.450 331.050 52.050 ;
        RECT 322.950 50.550 331.050 51.450 ;
        RECT 322.950 49.650 325.050 50.550 ;
        RECT 328.950 49.950 331.050 50.550 ;
        RECT -9.450 0.300 1043.400 2.700 ;
      LAYER metal2 ;
        RECT 139.950 958.950 142.050 961.050 ;
        RECT 151.950 959.100 154.050 961.200 ;
        RECT 221.400 960.450 222.600 960.600 ;
        RECT 290.400 960.450 291.600 960.600 ;
        RECT 221.400 959.400 225.450 960.450 ;
        RECT 77.400 953.400 78.600 955.650 ;
        RECT 77.400 937.050 78.450 953.400 ;
        RECT 140.400 937.050 141.450 958.950 ;
        RECT 152.400 958.350 153.600 959.100 ;
        RECT 221.400 958.350 222.600 959.400 ;
        RECT 224.400 937.050 225.450 959.400 ;
        RECT 290.400 959.400 294.450 960.450 ;
        RECT 290.400 958.350 291.600 959.400 ;
        RECT 293.400 937.050 294.450 959.400 ;
        RECT 77.400 935.400 82.050 937.050 ;
        RECT 140.400 935.400 145.050 937.050 ;
        RECT 224.400 935.400 229.050 937.050 ;
        RECT 78.000 934.950 82.050 935.400 ;
        RECT 141.000 934.950 145.050 935.400 ;
        RECT 225.000 934.950 229.050 935.400 ;
        RECT 292.950 934.950 295.050 937.050 ;
        RECT 34.950 931.950 37.050 934.050 ;
        RECT 35.400 882.600 36.450 931.950 ;
        RECT 167.400 914.400 168.600 916.650 ;
        RECT 167.400 895.050 168.450 914.400 ;
        RECT 166.950 892.950 169.050 895.050 ;
        RECT 178.950 894.450 181.050 895.050 ;
        RECT 176.400 893.400 181.050 894.450 ;
        RECT 176.400 882.600 177.450 893.400 ;
        RECT 178.950 892.950 181.050 893.400 ;
        RECT 35.400 880.350 36.600 882.600 ;
        RECT 176.400 880.350 177.600 882.600 ;
        RECT 179.400 859.050 180.450 892.950 ;
        RECT 172.950 856.950 175.050 859.050 ;
        RECT 178.950 856.950 181.050 859.050 ;
        RECT 173.400 847.050 174.450 856.950 ;
        RECT 151.950 844.950 154.050 847.050 ;
        RECT 172.950 844.950 175.050 847.050 ;
        RECT 152.400 841.050 153.450 844.950 ;
        RECT 151.950 838.950 154.050 841.050 ;
        RECT 35.400 836.400 36.600 838.650 ;
        RECT 35.400 820.050 36.450 836.400 ;
        RECT 151.950 832.950 154.050 835.050 ;
        RECT 34.950 817.950 37.050 820.050 ;
        RECT 49.950 817.950 52.050 820.050 ;
        RECT 11.400 804.450 12.600 804.600 ;
        RECT 11.400 803.400 15.450 804.450 ;
        RECT 11.400 802.350 12.600 803.400 ;
        RECT 14.400 781.050 15.450 803.400 ;
        RECT 50.400 781.050 51.450 817.950 ;
        RECT 152.400 804.450 153.450 832.950 ;
        RECT 155.400 804.450 156.600 804.600 ;
        RECT 152.400 803.400 156.600 804.450 ;
        RECT 155.400 802.350 156.600 803.400 ;
        RECT 13.950 778.950 16.050 781.050 ;
        RECT 37.950 778.950 40.050 781.050 ;
        RECT 49.950 778.950 52.050 781.050 ;
        RECT 178.950 778.950 181.050 781.050 ;
        RECT 35.400 681.450 36.600 682.650 ;
        RECT 38.400 681.450 39.450 778.950 ;
        RECT 179.400 726.600 180.450 778.950 ;
        RECT 179.400 724.350 180.600 726.600 ;
        RECT 35.400 680.400 39.450 681.450 ;
        RECT 38.400 667.050 39.450 680.400 ;
        RECT 37.950 664.950 40.050 667.050 ;
        RECT 55.950 664.950 58.050 667.050 ;
        RECT 56.400 609.600 57.450 664.950 ;
        RECT 104.400 648.450 105.600 648.600 ;
        RECT 104.400 647.400 108.450 648.450 ;
        RECT 104.400 646.350 105.600 647.400 ;
        RECT 107.400 625.050 108.450 647.400 ;
        RECT 106.950 622.950 109.050 625.050 ;
        RECT 121.950 622.950 124.050 625.050 ;
        RECT 56.400 607.350 57.600 609.600 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 175.800 568.950 177.900 571.050 ;
        RECT 161.400 568.350 162.600 568.950 ;
        RECT 176.400 561.450 177.450 568.950 ;
        RECT 176.400 560.400 180.450 561.450 ;
        RECT 179.400 547.050 180.450 560.400 ;
        RECT 67.950 541.950 70.050 544.050 ;
        RECT 97.950 541.950 100.050 547.050 ;
        RECT 178.950 544.950 181.050 547.050 ;
        RECT 607.950 544.950 610.050 547.050 ;
        RECT 643.950 544.950 646.050 547.050 ;
        RECT 721.950 544.950 724.050 547.050 ;
        RECT 883.950 544.950 886.050 547.050 ;
        RECT 11.400 525.000 12.600 526.650 ;
        RECT 10.950 520.950 13.050 525.000 ;
        RECT 68.400 523.050 69.450 541.950 ;
        RECT 590.400 525.900 591.600 526.650 ;
        RECT 608.400 526.050 609.450 544.950 ;
        RECT 589.950 523.800 592.050 525.900 ;
        RECT 607.950 523.950 610.050 526.050 ;
        RECT 67.950 520.950 70.050 523.050 ;
        RECT 644.400 522.450 645.450 544.950 ;
        RECT 722.400 529.050 723.450 544.950 ;
        RECT 721.950 526.950 724.050 529.050 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 644.400 521.400 648.450 522.450 ;
        RECT 647.400 504.450 648.450 521.400 ;
        RECT 647.400 503.400 651.450 504.450 ;
        RECT 650.400 492.600 651.450 503.400 ;
        RECT 761.400 492.600 762.450 523.950 ;
        RECT 884.400 514.050 885.450 544.950 ;
        RECT 874.950 511.950 877.050 514.050 ;
        RECT 883.950 511.950 886.050 514.050 ;
        RECT 875.400 492.600 876.450 511.950 ;
        RECT 596.400 492.450 597.600 492.600 ;
        RECT 593.400 491.400 597.600 492.450 ;
        RECT 593.400 469.050 594.450 491.400 ;
        RECT 596.400 490.350 597.600 491.400 ;
        RECT 650.400 490.350 651.600 492.600 ;
        RECT 761.400 490.350 762.600 492.600 ;
        RECT 875.400 490.350 876.600 492.600 ;
        RECT 593.400 467.400 598.050 469.050 ;
        RECT 594.000 466.950 598.050 467.400 ;
        RECT 790.950 466.950 793.050 469.050 ;
        RECT 11.400 447.450 12.600 448.650 ;
        RECT 779.400 447.900 780.600 448.650 ;
        RECT 791.400 448.050 792.450 466.950 ;
        RECT 8.400 446.400 12.600 447.450 ;
        RECT 8.400 427.050 9.450 446.400 ;
        RECT 778.950 445.800 781.050 447.900 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 872.400 446.400 873.600 448.650 ;
        RECT 872.400 427.050 873.450 446.400 ;
        RECT 7.950 424.950 10.050 427.050 ;
        RECT 34.950 424.950 37.050 427.050 ;
        RECT 871.950 424.950 874.050 427.050 ;
        RECT 877.950 424.950 880.050 427.050 ;
        RECT 35.400 400.050 36.450 424.950 ;
        RECT 61.950 418.950 64.050 421.050 ;
        RECT 100.950 418.950 103.050 421.050 ;
        RECT 62.400 414.600 63.450 418.950 ;
        RECT 62.400 412.350 63.600 414.600 ;
        RECT 34.950 397.950 37.050 400.050 ;
        RECT 52.950 397.950 55.050 400.050 ;
        RECT 53.400 391.050 54.450 397.950 ;
        RECT 101.400 391.050 102.450 418.950 ;
        RECT 878.400 406.050 879.450 424.950 ;
        RECT 877.950 403.950 880.050 406.050 ;
        RECT 901.950 403.950 904.050 406.050 ;
        RECT 52.950 388.950 55.050 391.050 ;
        RECT 100.950 388.950 103.050 391.050 ;
        RECT 902.400 388.050 903.450 403.950 ;
        RECT 901.950 385.950 904.050 388.050 ;
        RECT 821.400 369.450 822.600 370.650 ;
        RECT 821.400 368.400 825.450 369.450 ;
        RECT 824.400 355.050 825.450 368.400 ;
        RECT 842.400 368.400 843.600 370.650 ;
        RECT 842.400 366.450 843.450 368.400 ;
        RECT 839.400 365.400 843.450 366.450 ;
        RECT 823.950 352.950 826.050 355.050 ;
        RECT 829.950 352.950 832.050 355.050 ;
        RECT 830.400 349.050 831.450 352.950 ;
        RECT 839.400 349.050 840.450 365.400 ;
        RECT 829.950 346.950 832.050 349.050 ;
        RECT 838.950 346.950 841.050 349.050 ;
        RECT 11.400 336.450 12.600 336.600 ;
        RECT 428.400 336.450 429.600 336.600 ;
        RECT 11.400 335.400 15.450 336.450 ;
        RECT 11.400 334.350 12.600 335.400 ;
        RECT 14.400 313.050 15.450 335.400 ;
        RECT 425.400 335.400 429.600 336.450 ;
        RECT 425.400 313.050 426.450 335.400 ;
        RECT 428.400 334.350 429.600 335.400 ;
        RECT 830.400 316.050 831.450 346.950 ;
        RECT 829.950 313.950 832.050 316.050 ;
        RECT 859.950 313.950 862.050 316.050 ;
        RECT 13.950 310.950 16.050 313.050 ;
        RECT 385.950 310.950 388.050 313.050 ;
        RECT 424.950 310.950 427.050 313.050 ;
        RECT 433.950 310.950 436.050 313.050 ;
        RECT 529.950 310.950 532.050 313.050 ;
        RECT 586.950 310.950 589.050 313.050 ;
        RECT 386.400 286.050 387.450 310.950 ;
        RECT 434.400 292.050 435.450 310.950 ;
        RECT 433.950 289.950 436.050 292.050 ;
        RECT 458.400 291.900 459.600 292.650 ;
        RECT 457.950 289.800 460.050 291.900 ;
        RECT 527.400 291.450 528.600 292.650 ;
        RECT 530.400 291.450 531.450 310.950 ;
        RECT 860.400 304.050 861.450 313.950 ;
        RECT 880.950 306.450 883.050 307.050 ;
        RECT 880.950 305.400 885.450 306.450 ;
        RECT 859.950 301.950 862.050 304.050 ;
        RECT 880.950 301.950 883.050 305.400 ;
        RECT 884.400 295.050 885.450 305.400 ;
        RECT 883.950 292.950 886.050 295.050 ;
        RECT 860.400 291.900 861.600 292.650 ;
        RECT 527.400 290.400 531.450 291.450 ;
        RECT 859.950 289.800 862.050 291.900 ;
        RECT 379.950 283.950 382.050 286.050 ;
        RECT 385.950 283.950 388.050 286.050 ;
        RECT 380.400 258.600 381.450 283.950 ;
        RECT 380.400 256.350 381.600 258.600 ;
        RECT 449.400 258.450 450.600 258.600 ;
        RECT 446.400 257.400 450.600 258.450 ;
        RECT 446.400 235.050 447.450 257.400 ;
        RECT 449.400 256.350 450.600 257.400 ;
        RECT 470.400 258.450 471.600 258.600 ;
        RECT 470.400 257.400 474.450 258.450 ;
        RECT 470.400 256.350 471.600 257.400 ;
        RECT 473.400 235.050 474.450 257.400 ;
        RECT 730.950 257.100 733.050 259.200 ;
        RECT 731.400 256.350 732.600 257.100 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 830.400 258.450 831.600 258.600 ;
        RECT 830.400 257.400 834.450 258.450 ;
        RECT 743.400 235.050 744.450 256.950 ;
        RECT 830.400 256.350 831.600 257.400 ;
        RECT 442.950 232.950 445.050 235.050 ;
        RECT 445.950 232.950 448.050 235.050 ;
        RECT 472.950 232.950 475.050 235.050 ;
        RECT 502.950 232.950 505.050 235.050 ;
        RECT 733.950 232.950 736.050 235.050 ;
        RECT 742.950 232.950 745.050 235.050 ;
        RECT 431.400 213.900 432.600 214.650 ;
        RECT 443.400 214.050 444.450 232.950 ;
        RECT 503.400 214.050 504.450 232.950 ;
        RECT 833.400 232.050 834.450 257.400 ;
        RECT 832.950 229.950 835.050 232.050 ;
        RECT 838.950 229.950 841.050 235.050 ;
        RECT 847.950 232.950 850.050 235.050 ;
        RECT 833.400 219.600 834.450 229.950 ;
        RECT 833.400 217.350 834.600 219.600 ;
        RECT 430.950 211.800 433.050 213.900 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 530.400 213.900 531.600 214.650 ;
        RECT 529.950 211.800 532.050 213.900 ;
        RECT 848.400 208.050 849.450 232.950 ;
        RECT 869.400 212.400 870.600 214.650 ;
        RECT 869.400 208.050 870.450 212.400 ;
        RECT 847.950 205.950 850.050 208.050 ;
        RECT 868.950 205.950 871.050 208.050 ;
        RECT 467.400 180.450 468.600 180.600 ;
        RECT 878.400 180.450 879.600 180.600 ;
        RECT 467.400 179.400 471.450 180.450 ;
        RECT 467.400 178.350 468.600 179.400 ;
        RECT 470.400 157.050 471.450 179.400 ;
        RECT 875.400 179.400 879.600 180.450 ;
        RECT 875.400 157.050 876.450 179.400 ;
        RECT 878.400 178.350 879.600 179.400 ;
        RECT 352.950 154.950 355.050 157.050 ;
        RECT 466.950 155.400 471.450 157.050 ;
        RECT 466.950 154.950 471.000 155.400 ;
        RECT 835.950 154.950 838.050 157.050 ;
        RECT 874.950 154.950 877.050 157.050 ;
        RECT 913.950 154.950 916.050 157.050 ;
        RECT 353.400 102.600 354.450 154.950 ;
        RECT 836.400 123.450 837.450 154.950 ;
        RECT 833.400 122.400 837.450 123.450 ;
        RECT 353.400 100.350 354.600 102.600 ;
        RECT 767.400 102.450 768.600 102.600 ;
        RECT 764.400 101.400 768.600 102.450 ;
        RECT 764.400 79.050 765.450 101.400 ;
        RECT 767.400 100.350 768.600 101.400 ;
        RECT 301.950 76.950 304.050 79.050 ;
        RECT 328.950 76.950 331.050 79.050 ;
        RECT 760.950 77.400 765.450 79.050 ;
        RECT 760.950 76.950 765.000 77.400 ;
        RECT 302.400 24.600 303.450 76.950 ;
        RECT 329.400 52.050 330.450 76.950 ;
        RECT 833.400 67.050 834.450 122.400 ;
        RECT 914.400 121.050 915.450 154.950 ;
        RECT 886.950 118.950 889.050 121.050 ;
        RECT 913.950 118.950 916.050 121.050 ;
        RECT 887.400 102.600 888.450 118.950 ;
        RECT 887.400 100.350 888.600 102.600 ;
        RECT 967.950 76.950 970.050 79.050 ;
        RECT 823.950 64.950 826.050 67.050 ;
        RECT 832.950 64.950 835.050 67.050 ;
        RECT 322.950 49.650 325.050 51.750 ;
        RECT 328.950 49.950 331.050 52.050 ;
        RECT 323.400 24.600 324.450 49.650 ;
        RECT 824.400 49.050 825.450 64.950 ;
        RECT 833.400 63.600 834.450 64.950 ;
        RECT 833.400 61.350 834.600 63.600 ;
        RECT 848.400 56.400 849.600 58.650 ;
        RECT 848.400 49.050 849.450 56.400 ;
        RECT 823.950 46.950 826.050 49.050 ;
        RECT 847.950 46.950 850.050 49.050 ;
        RECT 302.400 22.350 303.600 24.600 ;
        RECT 323.400 22.350 324.600 24.600 ;
        RECT 853.950 23.100 856.050 25.200 ;
        RECT 854.400 22.350 855.600 23.100 ;
        RECT 874.950 22.950 877.050 25.050 ;
        RECT 899.400 24.450 900.600 24.600 ;
        RECT 899.400 23.400 903.450 24.450 ;
        RECT 875.400 13.050 876.450 22.950 ;
        RECT 899.400 22.350 900.600 23.400 ;
        RECT 902.400 13.050 903.450 23.400 ;
        RECT 968.400 13.050 969.450 76.950 ;
        RECT 874.950 10.950 877.050 13.050 ;
        RECT 901.950 10.950 904.050 13.050 ;
        RECT 967.950 10.950 970.050 13.050 ;
      LAYER metal3 ;
        RECT 139.950 960.600 142.050 961.050 ;
        RECT 151.950 960.600 154.050 961.200 ;
        RECT 139.950 959.400 154.050 960.600 ;
        RECT 139.950 958.950 142.050 959.400 ;
        RECT 151.950 959.100 154.050 959.400 ;
        RECT 166.950 894.600 169.050 895.050 ;
        RECT 178.950 894.600 181.050 895.050 ;
        RECT 166.950 893.400 181.050 894.600 ;
        RECT 166.950 892.950 169.050 893.400 ;
        RECT 178.950 892.950 181.050 893.400 ;
        RECT 151.950 846.600 154.050 847.050 ;
        RECT 172.950 846.600 175.050 847.050 ;
        RECT 151.950 845.400 175.050 846.600 ;
        RECT 151.950 844.950 154.050 845.400 ;
        RECT 172.950 844.950 175.050 845.400 ;
        RECT 34.950 819.600 37.050 820.050 ;
        RECT 49.950 819.600 52.050 820.050 ;
        RECT 34.950 818.400 52.050 819.600 ;
        RECT 34.950 817.950 37.050 818.400 ;
        RECT 49.950 817.950 52.050 818.400 ;
        RECT 37.950 780.600 40.050 781.050 ;
        RECT 49.950 780.600 52.050 781.050 ;
        RECT 37.950 779.400 52.050 780.600 ;
        RECT 37.950 778.950 40.050 779.400 ;
        RECT 49.950 778.950 52.050 779.400 ;
        RECT 37.950 666.600 40.050 667.050 ;
        RECT 55.950 666.600 58.050 667.050 ;
        RECT 37.950 665.400 58.050 666.600 ;
        RECT 37.950 664.950 40.050 665.400 ;
        RECT 55.950 664.950 58.050 665.400 ;
        RECT 106.950 624.600 109.050 625.050 ;
        RECT 121.950 624.600 124.050 625.050 ;
        RECT 106.950 623.400 124.050 624.600 ;
        RECT 106.950 622.950 109.050 623.400 ;
        RECT 121.950 622.950 124.050 623.400 ;
        RECT 160.950 570.600 163.050 571.050 ;
        RECT 175.800 570.600 177.900 571.050 ;
        RECT 160.950 569.400 177.900 570.600 ;
        RECT 160.950 568.950 163.050 569.400 ;
        RECT 175.800 568.950 177.900 569.400 ;
        RECT 67.950 543.600 70.050 544.050 ;
        RECT 97.950 543.600 100.050 544.050 ;
        RECT 67.950 542.400 100.050 543.600 ;
        RECT 67.950 541.950 70.050 542.400 ;
        RECT 97.950 541.950 100.050 542.400 ;
        RECT 589.950 525.600 592.050 525.900 ;
        RECT 607.950 525.600 610.050 526.050 ;
        RECT 589.950 524.400 610.050 525.600 ;
        RECT 721.950 525.600 724.050 529.050 ;
        RECT 760.950 525.600 763.050 526.050 ;
        RECT 721.950 525.000 763.050 525.600 ;
        RECT 722.400 524.400 763.050 525.000 ;
        RECT 589.950 523.800 592.050 524.400 ;
        RECT 607.950 523.950 610.050 524.400 ;
        RECT 760.950 523.950 763.050 524.400 ;
        RECT 10.950 522.600 13.050 523.050 ;
        RECT 67.950 522.600 70.050 523.050 ;
        RECT 10.950 521.400 70.050 522.600 ;
        RECT 10.950 520.950 13.050 521.400 ;
        RECT 67.950 520.950 70.050 521.400 ;
        RECT 874.950 513.600 877.050 514.050 ;
        RECT 883.950 513.600 886.050 514.050 ;
        RECT 874.950 512.400 886.050 513.600 ;
        RECT 874.950 511.950 877.050 512.400 ;
        RECT 883.950 511.950 886.050 512.400 ;
        RECT 778.950 447.600 781.050 447.900 ;
        RECT 790.950 447.600 793.050 448.050 ;
        RECT 778.950 446.400 793.050 447.600 ;
        RECT 778.950 445.800 781.050 446.400 ;
        RECT 790.950 445.950 793.050 446.400 ;
        RECT 7.950 426.600 10.050 427.050 ;
        RECT 34.950 426.600 37.050 427.050 ;
        RECT 7.950 425.400 37.050 426.600 ;
        RECT 7.950 424.950 10.050 425.400 ;
        RECT 34.950 424.950 37.050 425.400 ;
        RECT 61.950 420.600 64.050 421.050 ;
        RECT 100.950 420.600 103.050 421.050 ;
        RECT 61.950 419.400 103.050 420.600 ;
        RECT 61.950 418.950 64.050 419.400 ;
        RECT 100.950 418.950 103.050 419.400 ;
        RECT 877.950 405.600 880.050 406.050 ;
        RECT 901.950 405.600 904.050 406.050 ;
        RECT 877.950 404.400 904.050 405.600 ;
        RECT 877.950 403.950 880.050 404.400 ;
        RECT 901.950 403.950 904.050 404.400 ;
        RECT 34.950 399.600 37.050 400.050 ;
        RECT 52.950 399.600 55.050 400.050 ;
        RECT 34.950 398.400 55.050 399.600 ;
        RECT 34.950 397.950 37.050 398.400 ;
        RECT 52.950 397.950 55.050 398.400 ;
        RECT 823.950 354.600 826.050 355.050 ;
        RECT 829.950 354.600 832.050 355.050 ;
        RECT 823.950 353.400 832.050 354.600 ;
        RECT 823.950 352.950 826.050 353.400 ;
        RECT 829.950 352.950 832.050 353.400 ;
        RECT 829.950 348.600 832.050 349.050 ;
        RECT 838.950 348.600 841.050 349.050 ;
        RECT 829.950 347.400 841.050 348.600 ;
        RECT 829.950 346.950 832.050 347.400 ;
        RECT 838.950 346.950 841.050 347.400 ;
        RECT 829.950 315.600 832.050 316.050 ;
        RECT 859.950 315.600 862.050 316.050 ;
        RECT 829.950 314.400 862.050 315.600 ;
        RECT 829.950 313.950 832.050 314.400 ;
        RECT 859.950 313.950 862.050 314.400 ;
        RECT 529.950 312.600 532.050 313.050 ;
        RECT 586.950 312.600 589.050 313.050 ;
        RECT 529.950 311.400 589.050 312.600 ;
        RECT 529.950 310.950 532.050 311.400 ;
        RECT 586.950 310.950 589.050 311.400 ;
        RECT 859.950 303.600 862.050 304.050 ;
        RECT 880.950 303.600 883.050 304.050 ;
        RECT 859.950 302.400 883.050 303.600 ;
        RECT 859.950 301.950 862.050 302.400 ;
        RECT 880.950 301.950 883.050 302.400 ;
        RECT 433.950 291.600 436.050 292.050 ;
        RECT 457.950 291.600 460.050 291.900 ;
        RECT 433.950 290.400 460.050 291.600 ;
        RECT 433.950 289.950 436.050 290.400 ;
        RECT 457.950 289.800 460.050 290.400 ;
        RECT 859.950 291.600 862.050 291.900 ;
        RECT 883.950 291.600 886.050 295.050 ;
        RECT 859.950 291.000 886.050 291.600 ;
        RECT 859.950 290.400 885.600 291.000 ;
        RECT 859.950 289.800 862.050 290.400 ;
        RECT 379.950 285.600 382.050 286.050 ;
        RECT 385.950 285.600 388.050 286.050 ;
        RECT 379.950 284.400 388.050 285.600 ;
        RECT 379.950 283.950 382.050 284.400 ;
        RECT 385.950 283.950 388.050 284.400 ;
        RECT 730.950 258.600 733.050 259.200 ;
        RECT 742.950 258.600 745.050 259.050 ;
        RECT 730.950 257.400 745.050 258.600 ;
        RECT 730.950 257.100 733.050 257.400 ;
        RECT 742.950 256.950 745.050 257.400 ;
        RECT 733.950 234.600 736.050 235.050 ;
        RECT 742.950 234.600 745.050 235.050 ;
        RECT 733.950 233.400 745.050 234.600 ;
        RECT 733.950 232.950 736.050 233.400 ;
        RECT 742.950 232.950 745.050 233.400 ;
        RECT 832.950 231.600 835.050 232.050 ;
        RECT 838.950 231.600 841.050 232.050 ;
        RECT 832.950 230.400 841.050 231.600 ;
        RECT 832.950 229.950 835.050 230.400 ;
        RECT 838.950 229.950 841.050 230.400 ;
        RECT 430.950 213.600 433.050 213.900 ;
        RECT 442.950 213.600 445.050 214.050 ;
        RECT 430.950 212.400 445.050 213.600 ;
        RECT 430.950 211.800 433.050 212.400 ;
        RECT 442.950 211.950 445.050 212.400 ;
        RECT 502.950 213.600 505.050 214.050 ;
        RECT 529.950 213.600 532.050 213.900 ;
        RECT 502.950 212.400 532.050 213.600 ;
        RECT 502.950 211.950 505.050 212.400 ;
        RECT 529.950 211.800 532.050 212.400 ;
        RECT 847.950 207.600 850.050 208.050 ;
        RECT 868.950 207.600 871.050 208.050 ;
        RECT 847.950 206.400 871.050 207.600 ;
        RECT 847.950 205.950 850.050 206.400 ;
        RECT 868.950 205.950 871.050 206.400 ;
        RECT 886.950 120.600 889.050 121.050 ;
        RECT 913.950 120.600 916.050 121.050 ;
        RECT 886.950 119.400 916.050 120.600 ;
        RECT 886.950 118.950 889.050 119.400 ;
        RECT 913.950 118.950 916.050 119.400 ;
        RECT 823.950 66.600 826.050 67.050 ;
        RECT 832.950 66.600 835.050 67.050 ;
        RECT 823.950 65.400 835.050 66.600 ;
        RECT 823.950 64.950 826.050 65.400 ;
        RECT 832.950 64.950 835.050 65.400 ;
        RECT 823.950 48.600 826.050 49.050 ;
        RECT 847.950 48.600 850.050 49.050 ;
        RECT 823.950 47.400 850.050 48.600 ;
        RECT 823.950 46.950 826.050 47.400 ;
        RECT 847.950 46.950 850.050 47.400 ;
        RECT 853.950 24.600 856.050 25.200 ;
        RECT 874.950 24.600 877.050 25.050 ;
        RECT 853.950 23.400 877.050 24.600 ;
        RECT 853.950 23.100 856.050 23.400 ;
        RECT 874.950 22.950 877.050 23.400 ;
        RECT 874.950 12.600 877.050 13.050 ;
        RECT 901.950 12.600 904.050 13.050 ;
        RECT 967.950 12.600 970.050 13.050 ;
        RECT 874.950 11.400 970.050 12.600 ;
        RECT 874.950 10.950 877.050 11.400 ;
        RECT 901.950 10.950 904.050 11.400 ;
        RECT 967.950 10.950 970.050 11.400 ;
    END
  END vdd
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 317.400 762.450 318.600 762.600 ;
        RECT 314.400 761.400 318.600 762.450 ;
        RECT 314.400 706.050 315.450 761.400 ;
        RECT 317.400 760.350 318.600 761.400 ;
        RECT 283.950 703.950 286.050 706.050 ;
        RECT 313.950 703.950 316.050 706.050 ;
        RECT 82.950 697.950 85.050 700.050 ;
        RECT 1.950 643.950 4.050 646.050 ;
        RECT 2.400 589.050 3.450 643.950 ;
        RECT 83.400 643.050 84.450 697.950 ;
        RECT 284.400 697.050 285.450 703.950 ;
        RECT 283.950 694.950 286.050 697.050 ;
        RECT 89.400 645.000 90.600 646.650 ;
        RECT 82.950 640.950 85.050 643.050 ;
        RECT 88.950 640.950 91.050 645.000 ;
        RECT 1.950 586.950 4.050 589.050 ;
        RECT 61.950 586.950 64.050 589.050 ;
        RECT 62.400 553.050 63.450 586.950 ;
        RECT 61.950 550.950 64.050 553.050 ;
        RECT 127.950 547.950 130.050 550.050 ;
        RECT 128.400 486.450 129.450 547.950 ;
        RECT 746.400 489.900 747.600 490.650 ;
        RECT 730.950 487.800 733.050 489.900 ;
        RECT 745.950 487.800 748.050 489.900 ;
        RECT 125.400 485.400 129.450 486.450 ;
        RECT 125.400 379.050 126.450 485.400 ;
        RECT 731.400 433.050 732.450 487.800 ;
        RECT 730.950 430.950 733.050 433.050 ;
        RECT 742.950 430.950 745.050 433.050 ;
        RECT 373.950 394.950 376.050 397.050 ;
        RECT 205.950 388.950 208.050 391.050 ;
        RECT 232.950 388.950 235.050 391.050 ;
        RECT 206.400 379.050 207.450 388.950 ;
        RECT 233.400 385.050 234.450 388.950 ;
        RECT 374.400 388.050 375.450 394.950 ;
        RECT 388.950 394.800 391.050 396.900 ;
        RECT 373.950 385.950 376.050 388.050 ;
        RECT 232.950 382.950 235.050 385.050 ;
        RECT 100.950 376.950 103.050 379.050 ;
        RECT 124.950 376.950 127.050 379.050 ;
        RECT 205.950 376.950 208.050 379.050 ;
        RECT 89.400 333.900 90.600 334.650 ;
        RECT 101.400 333.900 102.450 376.950 ;
        RECT 88.950 331.800 91.050 333.900 ;
        RECT 100.950 331.800 103.050 333.900 ;
        RECT 389.400 316.050 390.450 394.800 ;
        RECT 743.400 351.450 744.450 430.950 ;
        RECT 743.400 350.400 747.450 351.450 ;
        RECT 746.400 339.450 747.450 350.400 ;
        RECT 746.400 338.400 750.450 339.450 ;
        RECT 388.950 313.950 391.050 316.050 ;
        RECT 400.950 313.950 403.050 316.050 ;
        RECT 401.400 294.600 402.450 313.950 ;
        RECT 401.400 294.450 402.600 294.600 ;
        RECT 401.400 293.400 405.450 294.450 ;
        RECT 401.400 292.350 402.600 293.400 ;
        RECT 404.400 274.050 405.450 293.400 ;
        RECT 403.950 271.950 406.050 274.050 ;
        RECT 445.950 271.950 448.050 274.050 ;
        RECT 446.400 265.050 447.450 271.950 ;
        RECT 445.950 262.950 448.050 265.050 ;
        RECT 532.950 262.950 535.050 265.050 ;
        RECT 533.400 193.050 534.450 262.950 ;
        RECT 749.400 193.050 750.450 338.400 ;
        RECT 532.950 190.950 535.050 193.050 ;
        RECT 559.950 190.950 562.050 193.050 ;
        RECT 748.950 190.950 751.050 193.050 ;
        RECT 757.950 190.950 760.050 193.050 ;
        RECT 560.400 177.450 561.450 190.950 ;
        RECT 563.400 177.450 564.600 178.650 ;
        RECT 560.400 176.400 564.600 177.450 ;
        RECT 758.400 138.600 759.450 190.950 ;
        RECT 758.400 136.350 759.600 138.600 ;
      LAYER metal3 ;
        RECT 283.950 705.600 286.050 706.050 ;
        RECT 313.950 705.600 316.050 706.050 ;
        RECT 283.950 704.400 316.050 705.600 ;
        RECT 283.950 703.950 286.050 704.400 ;
        RECT 313.950 703.950 316.050 704.400 ;
        RECT 82.950 699.600 85.050 700.050 ;
        RECT 82.950 698.400 165.600 699.600 ;
        RECT 82.950 697.950 85.050 698.400 ;
        RECT 164.400 696.600 165.600 698.400 ;
        RECT 283.950 696.600 286.050 697.050 ;
        RECT 164.400 695.400 286.050 696.600 ;
        RECT 283.950 694.950 286.050 695.400 ;
        RECT 1.950 645.600 4.050 646.050 ;
        RECT -3.600 644.400 4.050 645.600 ;
        RECT 1.950 643.950 4.050 644.400 ;
        RECT 2.400 642.600 3.600 643.950 ;
        RECT 82.950 642.600 85.050 643.050 ;
        RECT 88.950 642.600 91.050 643.050 ;
        RECT 2.400 641.400 91.050 642.600 ;
        RECT 82.950 640.950 85.050 641.400 ;
        RECT 88.950 640.950 91.050 641.400 ;
        RECT 1.950 588.600 4.050 589.050 ;
        RECT 61.950 588.600 64.050 589.050 ;
        RECT 1.950 587.400 64.050 588.600 ;
        RECT 1.950 586.950 4.050 587.400 ;
        RECT 61.950 586.950 64.050 587.400 ;
        RECT 61.950 552.600 64.050 553.050 ;
        RECT 61.950 551.400 81.600 552.600 ;
        RECT 61.950 550.950 64.050 551.400 ;
        RECT 80.400 549.600 81.600 551.400 ;
        RECT 127.950 549.600 130.050 550.050 ;
        RECT 80.400 548.400 130.050 549.600 ;
        RECT 127.950 547.950 130.050 548.400 ;
        RECT 730.950 489.450 733.050 489.900 ;
        RECT 745.950 489.450 748.050 489.900 ;
        RECT 730.950 488.250 748.050 489.450 ;
        RECT 730.950 487.800 733.050 488.250 ;
        RECT 745.950 487.800 748.050 488.250 ;
        RECT 730.950 432.600 733.050 433.050 ;
        RECT 742.950 432.600 745.050 433.050 ;
        RECT 730.950 431.400 745.050 432.600 ;
        RECT 730.950 430.950 733.050 431.400 ;
        RECT 742.950 430.950 745.050 431.400 ;
        RECT 373.950 396.600 376.050 397.050 ;
        RECT 388.950 396.600 391.050 396.900 ;
        RECT 373.950 395.400 391.050 396.600 ;
        RECT 373.950 394.950 376.050 395.400 ;
        RECT 388.950 394.800 391.050 395.400 ;
        RECT 205.950 390.600 208.050 391.050 ;
        RECT 232.950 390.600 235.050 391.050 ;
        RECT 205.950 389.400 235.050 390.600 ;
        RECT 205.950 388.950 208.050 389.400 ;
        RECT 232.950 388.950 235.050 389.400 ;
        RECT 373.950 387.600 376.050 388.050 ;
        RECT 251.400 386.400 376.050 387.600 ;
        RECT 232.950 384.600 235.050 385.050 ;
        RECT 251.400 384.600 252.600 386.400 ;
        RECT 373.950 385.950 376.050 386.400 ;
        RECT 232.950 383.400 252.600 384.600 ;
        RECT 232.950 382.950 235.050 383.400 ;
        RECT 100.950 378.600 103.050 379.050 ;
        RECT 124.950 378.600 127.050 379.050 ;
        RECT 205.950 378.600 208.050 379.050 ;
        RECT 100.950 377.400 208.050 378.600 ;
        RECT 100.950 376.950 103.050 377.400 ;
        RECT 124.950 376.950 127.050 377.400 ;
        RECT 205.950 376.950 208.050 377.400 ;
        RECT 88.950 333.450 91.050 333.900 ;
        RECT 100.950 333.450 103.050 333.900 ;
        RECT 88.950 332.250 103.050 333.450 ;
        RECT 88.950 331.800 91.050 332.250 ;
        RECT 100.950 331.800 103.050 332.250 ;
        RECT 388.950 315.600 391.050 316.050 ;
        RECT 400.950 315.600 403.050 316.050 ;
        RECT 388.950 314.400 403.050 315.600 ;
        RECT 388.950 313.950 391.050 314.400 ;
        RECT 400.950 313.950 403.050 314.400 ;
        RECT 403.950 273.600 406.050 274.050 ;
        RECT 445.950 273.600 448.050 274.050 ;
        RECT 403.950 272.400 448.050 273.600 ;
        RECT 403.950 271.950 406.050 272.400 ;
        RECT 445.950 271.950 448.050 272.400 ;
        RECT 445.950 264.600 448.050 265.050 ;
        RECT 532.950 264.600 535.050 265.050 ;
        RECT 445.950 263.400 535.050 264.600 ;
        RECT 445.950 262.950 448.050 263.400 ;
        RECT 532.950 262.950 535.050 263.400 ;
        RECT 532.950 192.600 535.050 193.050 ;
        RECT 559.950 192.600 562.050 193.050 ;
        RECT 748.950 192.600 751.050 193.050 ;
        RECT 757.950 192.600 760.050 193.050 ;
        RECT 532.950 191.400 760.050 192.600 ;
        RECT 532.950 190.950 535.050 191.400 ;
        RECT 559.950 190.950 562.050 191.400 ;
        RECT 748.950 190.950 751.050 191.400 ;
        RECT 757.950 190.950 760.050 191.400 ;
    END
  END clk
  PIN down
    PORT
      LAYER metal2 ;
        RECT 931.950 541.950 934.050 544.050 ;
        RECT 1042.950 541.950 1045.050 544.050 ;
        RECT 892.950 538.950 895.050 541.050 ;
        RECT 893.400 528.450 894.450 538.950 ;
        RECT 932.400 538.050 933.450 541.950 ;
        RECT 931.950 535.950 934.050 538.050 ;
        RECT 1043.400 529.050 1044.450 541.950 ;
        RECT 896.400 528.450 897.600 528.600 ;
        RECT 893.400 527.400 897.600 528.450 ;
        RECT 896.400 526.350 897.600 527.400 ;
        RECT 1042.950 526.950 1045.050 529.050 ;
      LAYER metal3 ;
        RECT 931.950 543.600 934.050 544.050 ;
        RECT 1042.950 543.600 1045.050 544.050 ;
        RECT 931.950 542.400 1045.050 543.600 ;
        RECT 931.950 541.950 934.050 542.400 ;
        RECT 1042.950 541.950 1045.050 542.400 ;
        RECT 892.950 540.600 895.050 541.050 ;
        RECT 892.950 539.400 915.600 540.600 ;
        RECT 892.950 538.950 895.050 539.400 ;
        RECT 914.400 537.600 915.600 539.400 ;
        RECT 931.950 537.600 934.050 538.050 ;
        RECT 914.400 536.400 934.050 537.600 ;
        RECT 931.950 535.950 934.050 536.400 ;
        RECT 1042.950 528.600 1045.050 529.050 ;
        RECT 1042.950 527.400 1050.600 528.600 ;
        RECT 1042.950 526.950 1045.050 527.400 ;
    END
  END down
  PIN hsync
    PORT
      LAYER metal2 ;
        RECT 17.400 723.900 18.600 724.650 ;
        RECT 16.950 721.800 19.050 723.900 ;
      LAYER metal3 ;
        RECT 16.950 723.600 19.050 723.900 ;
        RECT -3.600 722.400 19.050 723.600 ;
        RECT 16.950 721.800 19.050 722.400 ;
    END
  END hsync
  PIN p_tick
    PORT
      LAYER metal2 ;
        RECT 16.950 761.100 19.050 763.200 ;
        RECT 17.400 760.350 18.600 761.100 ;
      LAYER metal3 ;
        RECT 16.950 762.600 19.050 763.200 ;
        RECT -3.600 761.400 19.050 762.600 ;
        RECT 16.950 761.100 19.050 761.400 ;
    END
  END p_tick
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 1.950 916.950 4.050 919.050 ;
        RECT 2.400 912.900 3.450 916.950 ;
        RECT 20.400 912.900 21.600 913.650 ;
        RECT 1.950 910.800 4.050 912.900 ;
        RECT 19.950 910.800 22.050 912.900 ;
        RECT 2.400 805.050 3.450 910.800 ;
        RECT 1.950 802.950 4.050 805.050 ;
        RECT 1.800 796.950 3.900 799.050 ;
        RECT 2.400 793.050 3.450 796.950 ;
        RECT 1.950 790.950 4.050 793.050 ;
        RECT 7.950 790.950 10.050 793.050 ;
        RECT 8.400 559.050 9.450 790.950 ;
        RECT 7.950 556.950 10.050 559.050 ;
        RECT 52.950 556.950 55.050 559.050 ;
        RECT 53.400 535.050 54.450 556.950 ;
        RECT 52.950 532.950 55.050 535.050 ;
        RECT 73.950 532.950 76.050 535.050 ;
        RECT 74.400 478.050 75.450 532.950 ;
        RECT 73.950 475.950 76.050 478.050 ;
        RECT 208.950 475.950 211.050 478.050 ;
        RECT 209.400 444.450 210.450 475.950 ;
        RECT 212.400 444.450 213.600 445.650 ;
        RECT 209.400 443.400 213.600 444.450 ;
      LAYER metal3 ;
        RECT 1.950 918.600 4.050 919.050 ;
        RECT -3.600 917.400 4.050 918.600 ;
        RECT 1.950 916.950 4.050 917.400 ;
        RECT 1.950 912.450 4.050 912.900 ;
        RECT 19.950 912.450 22.050 912.900 ;
        RECT 1.950 911.250 22.050 912.450 ;
        RECT 1.950 910.800 4.050 911.250 ;
        RECT 19.950 910.800 22.050 911.250 ;
        RECT 1.950 802.950 4.050 805.050 ;
        RECT 2.400 799.050 3.600 802.950 ;
        RECT 1.800 796.950 3.900 799.050 ;
        RECT 1.950 792.600 4.050 793.050 ;
        RECT 7.950 792.600 10.050 793.050 ;
        RECT 1.950 791.400 10.050 792.600 ;
        RECT 1.950 790.950 4.050 791.400 ;
        RECT 7.950 790.950 10.050 791.400 ;
        RECT 7.950 558.600 10.050 559.050 ;
        RECT 52.950 558.600 55.050 559.050 ;
        RECT 7.950 557.400 55.050 558.600 ;
        RECT 7.950 556.950 10.050 557.400 ;
        RECT 52.950 556.950 55.050 557.400 ;
        RECT 52.950 534.600 55.050 535.050 ;
        RECT 73.950 534.600 76.050 535.050 ;
        RECT 52.950 533.400 76.050 534.600 ;
        RECT 52.950 532.950 55.050 533.400 ;
        RECT 73.950 532.950 76.050 533.400 ;
        RECT 73.950 477.600 76.050 478.050 ;
        RECT 208.950 477.600 211.050 478.050 ;
        RECT 73.950 476.400 211.050 477.600 ;
        RECT 73.950 475.950 76.050 476.400 ;
        RECT 208.950 475.950 211.050 476.400 ;
    END
  END reset
  PIN rgb[11]
    PORT
      LAYER metal2 ;
        RECT 16.950 683.100 19.050 685.200 ;
        RECT 17.400 682.350 18.600 683.100 ;
      LAYER metal3 ;
        RECT 16.950 684.600 19.050 685.200 ;
        RECT -3.600 683.400 19.050 684.600 ;
        RECT 16.950 683.100 19.050 683.400 ;
    END
  END rgb[11]
  PIN rgb[10]
    PORT
      LAYER metal2 ;
        RECT 17.400 21.900 18.600 22.650 ;
        RECT 16.950 19.800 19.050 21.900 ;
      LAYER metal3 ;
        RECT 16.950 21.600 19.050 21.900 ;
        RECT -3.600 20.400 19.050 21.600 ;
        RECT 16.950 19.800 19.050 20.400 ;
    END
  END rgb[10]
  PIN rgb[9]
    PORT
      LAYER metal2 ;
        RECT 71.400 983.400 75.450 984.450 ;
        RECT 74.400 961.050 75.450 983.400 ;
        RECT 73.950 958.950 76.050 961.050 ;
        RECT 71.400 957.900 72.600 958.650 ;
        RECT 70.950 955.800 73.050 957.900 ;
      LAYER metal3 ;
        RECT 70.950 957.600 73.050 957.900 ;
        RECT 73.950 957.600 76.050 961.050 ;
        RECT 70.950 957.000 76.050 957.600 ;
        RECT 70.950 956.400 75.600 957.000 ;
        RECT 70.950 955.800 73.050 956.400 ;
    END
  END rgb[9]
  PIN rgb[8]
    PORT
      LAYER metal2 ;
        RECT 242.400 20.400 243.600 22.650 ;
        RECT 242.400 -2.550 243.450 20.400 ;
        RECT 239.400 -3.600 243.450 -2.550 ;
    END
  END rgb[8]
  PIN rgb[7]
    PORT
      LAYER metal2 ;
        RECT 16.950 605.100 19.050 607.200 ;
        RECT 17.400 604.350 18.600 605.100 ;
      LAYER metal3 ;
        RECT 16.950 606.600 19.050 607.200 ;
        RECT -3.600 605.400 19.050 606.600 ;
        RECT 16.950 605.100 19.050 605.400 ;
    END
  END rgb[7]
  PIN rgb[6]
    PORT
      LAYER metal2 ;
        RECT 41.400 20.400 42.600 22.650 ;
        RECT 41.400 -2.550 42.450 20.400 ;
        RECT 41.400 -3.600 45.450 -2.550 ;
    END
  END rgb[6]
  PIN rgb[5]
    PORT
      LAYER metal2 ;
        RECT 16.950 839.100 19.050 841.200 ;
        RECT 17.400 838.350 18.600 839.100 ;
      LAYER metal3 ;
        RECT 16.950 840.600 19.050 841.200 ;
        RECT -3.600 839.400 19.050 840.600 ;
        RECT 16.950 839.100 19.050 839.400 ;
    END
  END rgb[5]
  PIN rgb[4]
    PORT
      LAYER metal2 ;
        RECT 197.400 20.400 198.600 22.650 ;
        RECT 197.400 -2.550 198.450 20.400 ;
        RECT 194.400 -3.600 198.450 -2.550 ;
    END
  END rgb[4]
  PIN rgb[3]
    PORT
      LAYER metal2 ;
        RECT 17.400 957.900 18.600 958.650 ;
        RECT 16.950 955.800 19.050 957.900 ;
      LAYER metal3 ;
        RECT 16.950 957.600 19.050 957.900 ;
        RECT -3.600 956.400 19.050 957.600 ;
        RECT 16.950 955.800 19.050 956.400 ;
    END
  END rgb[3]
  PIN rgb[2]
    PORT
      LAYER metal2 ;
        RECT 71.400 20.400 72.600 22.650 ;
        RECT 71.400 -2.550 72.450 20.400 ;
        RECT 68.400 -3.600 72.450 -2.550 ;
    END
  END rgb[2]
  PIN rgb[1]
    PORT
      LAYER metal2 ;
        RECT 44.400 979.050 45.450 984.450 ;
        RECT 43.950 976.950 46.050 979.050 ;
        RECT 49.950 976.950 52.050 979.050 ;
        RECT 47.400 957.450 48.600 958.650 ;
        RECT 50.400 957.450 51.450 976.950 ;
        RECT 47.400 956.400 51.450 957.450 ;
      LAYER metal3 ;
        RECT 43.950 978.600 46.050 979.050 ;
        RECT 49.950 978.600 52.050 979.050 ;
        RECT 43.950 977.400 52.050 978.600 ;
        RECT 43.950 976.950 46.050 977.400 ;
        RECT 49.950 976.950 52.050 977.400 ;
    END
  END rgb[1]
  PIN rgb[0]
    PORT
      LAYER metal2 ;
        RECT 167.400 20.400 168.600 22.650 ;
        RECT 167.400 -2.550 168.450 20.400 ;
        RECT 167.400 -3.600 171.450 -2.550 ;
    END
  END rgb[0]
  PIN up
    PORT
      LAYER metal2 ;
        RECT 1024.950 338.100 1027.050 340.200 ;
        RECT 1025.400 337.350 1026.600 338.100 ;
        RECT 1007.400 333.900 1008.600 334.650 ;
        RECT 1006.950 331.800 1009.050 333.900 ;
      LAYER metal3 ;
        RECT 1024.950 339.600 1027.050 340.200 ;
        RECT 1024.950 338.400 1050.600 339.600 ;
        RECT 1024.950 338.100 1027.050 338.400 ;
        RECT 1006.950 333.600 1009.050 333.900 ;
        RECT 1025.400 333.600 1026.600 338.100 ;
        RECT 1006.950 332.400 1026.600 333.600 ;
        RECT 1049.400 332.400 1050.600 338.400 ;
        RECT 1006.950 331.800 1009.050 332.400 ;
    END
  END up
  PIN vsync
    PORT
      LAYER metal2 ;
        RECT 65.400 967.050 66.450 984.450 ;
        RECT 64.950 964.950 67.050 967.050 ;
        RECT 70.950 949.950 73.050 952.050 ;
        RECT 71.400 918.600 72.450 949.950 ;
        RECT 71.400 916.350 72.600 918.600 ;
      LAYER metal3 ;
        RECT 64.950 964.950 67.050 967.050 ;
        RECT 65.400 951.600 66.600 964.950 ;
        RECT 70.950 951.600 73.050 952.050 ;
        RECT 65.400 950.400 73.050 951.600 ;
        RECT 70.950 949.950 73.050 950.400 ;
    END
  END vsync
  OBS
      LAYER metal1 ;
        RECT 17.100 968.400 18.900 974.400 ;
        RECT 20.100 968.400 21.900 975.000 ;
        RECT 23.100 971.400 24.900 974.400 ;
        RECT 17.100 961.050 18.300 968.400 ;
        RECT 23.700 967.500 24.900 971.400 ;
        RECT 19.200 966.600 24.900 967.500 ;
        RECT 41.100 971.400 42.900 974.400 ;
        RECT 41.100 967.500 42.300 971.400 ;
        RECT 44.100 968.400 45.900 975.000 ;
        RECT 47.100 968.400 48.900 974.400 ;
        RECT 41.100 966.600 46.800 967.500 ;
        RECT 19.200 965.700 21.000 966.600 ;
        RECT 17.100 958.950 19.200 961.050 ;
        RECT 17.100 951.600 18.300 958.950 ;
        RECT 20.100 954.300 21.000 965.700 ;
        RECT 45.000 965.700 46.800 966.600 ;
        RECT 22.500 958.950 24.600 961.050 ;
        RECT 22.800 957.150 24.600 958.950 ;
        RECT 41.400 958.950 43.500 961.050 ;
        RECT 41.400 957.150 43.200 958.950 ;
        RECT 19.200 953.400 21.000 954.300 ;
        RECT 45.000 954.300 45.900 965.700 ;
        RECT 47.700 961.050 48.900 968.400 ;
        RECT 65.100 971.400 66.900 974.400 ;
        RECT 65.100 967.500 66.300 971.400 ;
        RECT 68.100 968.400 69.900 975.000 ;
        RECT 71.100 968.400 72.900 974.400 ;
        RECT 65.100 966.600 70.800 967.500 ;
        RECT 69.000 965.700 70.800 966.600 ;
        RECT 46.800 958.950 48.900 961.050 ;
        RECT 45.000 953.400 46.800 954.300 ;
        RECT 19.200 952.500 24.900 953.400 ;
        RECT 17.100 939.600 18.900 951.600 ;
        RECT 20.100 939.000 21.900 949.800 ;
        RECT 23.700 945.600 24.900 952.500 ;
        RECT 23.100 939.600 24.900 945.600 ;
        RECT 41.100 952.500 46.800 953.400 ;
        RECT 41.100 945.600 42.300 952.500 ;
        RECT 47.700 951.600 48.900 958.950 ;
        RECT 65.400 958.950 67.500 961.050 ;
        RECT 65.400 957.150 67.200 958.950 ;
        RECT 69.000 954.300 69.900 965.700 ;
        RECT 71.700 961.050 72.900 968.400 ;
        RECT 70.800 958.950 72.900 961.050 ;
        RECT 69.000 953.400 70.800 954.300 ;
        RECT 41.100 939.600 42.900 945.600 ;
        RECT 44.100 939.000 45.900 949.800 ;
        RECT 47.100 939.600 48.900 951.600 ;
        RECT 65.100 952.500 70.800 953.400 ;
        RECT 65.100 945.600 66.300 952.500 ;
        RECT 71.700 951.600 72.900 958.950 ;
        RECT 65.100 939.600 66.900 945.600 ;
        RECT 68.100 939.000 69.900 949.800 ;
        RECT 71.100 939.600 72.900 951.600 ;
        RECT 74.700 968.400 76.500 974.400 ;
        RECT 80.100 968.400 81.900 975.000 ;
        RECT 85.500 968.400 87.300 974.400 ;
        RECT 89.700 971.400 91.500 974.400 ;
        RECT 92.700 971.400 94.500 974.400 ;
        RECT 95.700 971.400 97.500 974.400 ;
        RECT 98.700 971.400 100.500 975.000 ;
        RECT 89.700 969.300 91.800 971.400 ;
        RECT 92.700 969.300 94.800 971.400 ;
        RECT 95.700 969.300 97.800 971.400 ;
        RECT 103.200 970.500 105.000 974.400 ;
        RECT 106.200 971.400 108.000 975.000 ;
        RECT 109.200 971.400 111.000 974.400 ;
        RECT 112.200 971.400 114.000 974.400 ;
        RECT 115.200 971.400 117.000 974.400 ;
        RECT 118.200 971.400 120.000 974.400 ;
        RECT 99.600 969.600 101.400 970.500 ;
        RECT 98.700 968.400 101.400 969.600 ;
        RECT 103.200 968.400 105.900 970.500 ;
        RECT 109.200 969.300 111.300 971.400 ;
        RECT 112.200 969.300 114.300 971.400 ;
        RECT 115.200 969.300 117.300 971.400 ;
        RECT 118.200 969.300 120.300 971.400 ;
        RECT 122.400 969.600 124.200 974.400 ;
        RECT 122.400 968.400 126.600 969.600 ;
        RECT 127.500 968.400 129.300 975.000 ;
        RECT 132.900 968.400 134.700 974.400 ;
        RECT 74.700 964.800 75.900 968.400 ;
        RECT 85.800 967.500 87.300 968.400 ;
        RECT 94.800 967.800 96.600 968.400 ;
        RECT 98.700 967.800 99.600 968.400 ;
        RECT 78.900 966.300 87.300 967.500 ;
        RECT 92.400 966.600 99.600 967.800 ;
        RECT 114.300 966.600 120.900 968.400 ;
        RECT 78.900 965.700 80.700 966.300 ;
        RECT 89.400 964.800 91.500 965.700 ;
        RECT 74.700 963.600 91.500 964.800 ;
        RECT 92.400 963.600 93.300 966.600 ;
        RECT 97.800 963.900 99.600 964.800 ;
        RECT 107.100 964.500 108.900 966.300 ;
        RECT 125.100 965.100 126.600 968.400 ;
        RECT 100.800 963.900 102.900 964.050 ;
        RECT 74.700 947.400 75.900 963.600 ;
        RECT 92.400 961.800 94.200 963.600 ;
        RECT 97.800 963.000 102.900 963.900 ;
        RECT 100.800 961.950 102.900 963.000 ;
        RECT 107.100 963.900 109.200 964.500 ;
        RECT 107.100 962.400 124.200 963.900 ;
        RECT 125.100 963.300 132.900 965.100 ;
        RECT 122.700 960.900 129.300 962.400 ;
        RECT 77.100 959.700 121.500 960.900 ;
        RECT 77.100 958.050 78.900 959.700 ;
        RECT 76.800 955.950 78.900 958.050 ;
        RECT 82.800 957.750 84.900 958.050 ;
        RECT 95.400 957.900 97.200 958.500 ;
        RECT 104.400 957.900 117.900 958.800 ;
        RECT 82.800 955.950 86.700 957.750 ;
        RECT 95.400 956.700 106.500 957.900 ;
        RECT 84.900 955.200 86.700 955.950 ;
        RECT 104.400 955.800 106.500 956.700 ;
        RECT 108.000 955.200 111.900 957.000 ;
        RECT 117.000 956.700 117.900 957.900 ;
        RECT 84.900 954.300 98.400 955.200 ;
        RECT 109.800 954.900 111.900 955.200 ;
        RECT 116.100 954.900 117.900 956.700 ;
        RECT 120.600 958.200 121.500 959.700 ;
        RECT 120.600 956.400 125.700 958.200 ;
        RECT 127.800 958.050 129.300 960.900 ;
        RECT 127.800 955.950 129.900 958.050 ;
        RECT 97.200 953.700 98.400 954.300 ;
        RECT 131.100 953.700 132.900 954.300 ;
        RECT 92.400 952.500 94.500 952.800 ;
        RECT 97.200 952.500 132.900 953.700 ;
        RECT 82.500 951.300 94.500 952.500 ;
        RECT 133.800 951.600 134.700 968.400 ;
        RECT 82.500 950.700 84.300 951.300 ;
        RECT 92.400 950.700 94.500 951.300 ;
        RECT 97.200 950.400 114.900 951.600 ;
        RECT 79.200 949.800 81.000 950.100 ;
        RECT 97.200 949.800 98.400 950.400 ;
        RECT 79.200 948.600 98.400 949.800 ;
        RECT 112.800 949.500 114.900 950.400 ;
        RECT 118.200 950.700 134.700 951.600 ;
        RECT 118.200 949.500 120.300 950.700 ;
        RECT 79.200 948.300 81.000 948.600 ;
        RECT 74.700 946.500 78.300 947.400 ;
        RECT 77.400 945.600 78.300 946.500 ;
        RECT 74.700 939.000 76.500 945.600 ;
        RECT 77.400 944.700 79.500 945.600 ;
        RECT 77.700 939.600 79.500 944.700 ;
        RECT 80.700 939.000 82.500 945.600 ;
        RECT 83.700 939.600 85.500 948.600 ;
        RECT 95.700 945.600 97.800 947.700 ;
        RECT 103.200 947.100 106.500 949.200 ;
        RECT 86.700 939.000 88.500 945.600 ;
        RECT 90.300 942.600 92.400 944.700 ;
        RECT 93.300 942.600 95.400 944.700 ;
        RECT 90.300 939.600 92.100 942.600 ;
        RECT 93.300 939.600 95.100 942.600 ;
        RECT 96.300 939.600 98.100 945.600 ;
        RECT 99.300 939.000 101.100 945.600 ;
        RECT 103.200 939.600 105.000 947.100 ;
        RECT 109.200 945.600 111.900 949.500 ;
        RECT 124.200 948.600 129.900 949.800 ;
        RECT 121.500 947.700 123.300 948.300 ;
        RECT 115.200 946.500 123.300 947.700 ;
        RECT 115.200 945.600 117.300 946.500 ;
        RECT 124.200 945.600 125.400 948.600 ;
        RECT 128.100 948.000 129.900 948.600 ;
        RECT 133.800 947.400 134.700 950.700 ;
        RECT 130.800 946.500 134.700 947.400 ;
        RECT 136.500 971.400 138.300 974.400 ;
        RECT 139.500 971.400 141.300 975.000 ;
        RECT 136.500 958.050 138.000 971.400 ;
        RECT 143.700 968.400 145.500 974.400 ;
        RECT 149.100 968.400 150.900 975.000 ;
        RECT 154.500 968.400 156.300 974.400 ;
        RECT 158.700 971.400 160.500 974.400 ;
        RECT 161.700 971.400 163.500 974.400 ;
        RECT 164.700 971.400 166.500 974.400 ;
        RECT 167.700 971.400 169.500 975.000 ;
        RECT 158.700 969.300 160.800 971.400 ;
        RECT 161.700 969.300 163.800 971.400 ;
        RECT 164.700 969.300 166.800 971.400 ;
        RECT 172.200 970.500 174.000 974.400 ;
        RECT 175.200 971.400 177.000 975.000 ;
        RECT 178.200 971.400 180.000 974.400 ;
        RECT 181.200 971.400 183.000 974.400 ;
        RECT 184.200 971.400 186.000 974.400 ;
        RECT 187.200 971.400 189.000 974.400 ;
        RECT 168.600 969.600 170.400 970.500 ;
        RECT 167.700 968.400 170.400 969.600 ;
        RECT 172.200 968.400 174.900 970.500 ;
        RECT 178.200 969.300 180.300 971.400 ;
        RECT 181.200 969.300 183.300 971.400 ;
        RECT 184.200 969.300 186.300 971.400 ;
        RECT 187.200 969.300 189.300 971.400 ;
        RECT 191.400 969.600 193.200 974.400 ;
        RECT 191.400 968.400 195.600 969.600 ;
        RECT 196.500 968.400 198.300 975.000 ;
        RECT 201.900 968.400 203.700 974.400 ;
        RECT 143.700 964.800 144.900 968.400 ;
        RECT 154.800 967.500 156.300 968.400 ;
        RECT 163.800 967.800 165.600 968.400 ;
        RECT 167.700 967.800 168.600 968.400 ;
        RECT 147.900 966.300 156.300 967.500 ;
        RECT 161.400 966.600 168.600 967.800 ;
        RECT 183.300 966.600 189.900 968.400 ;
        RECT 147.900 965.700 149.700 966.300 ;
        RECT 158.400 964.800 160.500 965.700 ;
        RECT 143.700 963.600 160.500 964.800 ;
        RECT 161.400 963.600 162.300 966.600 ;
        RECT 166.800 963.900 168.600 964.800 ;
        RECT 176.100 964.500 177.900 966.300 ;
        RECT 194.100 965.100 195.600 968.400 ;
        RECT 169.800 963.900 171.900 964.050 ;
        RECT 136.500 955.950 138.900 958.050 ;
        RECT 130.800 945.600 132.000 946.500 ;
        RECT 136.500 945.600 138.000 955.950 ;
        RECT 143.700 947.400 144.900 963.600 ;
        RECT 161.400 961.800 163.200 963.600 ;
        RECT 166.800 963.000 171.900 963.900 ;
        RECT 169.800 961.950 171.900 963.000 ;
        RECT 176.100 963.900 178.200 964.500 ;
        RECT 176.100 962.400 193.200 963.900 ;
        RECT 194.100 963.300 201.900 965.100 ;
        RECT 191.700 960.900 198.300 962.400 ;
        RECT 146.100 959.700 190.500 960.900 ;
        RECT 146.100 958.050 147.900 959.700 ;
        RECT 145.800 955.950 147.900 958.050 ;
        RECT 151.800 957.750 153.900 958.050 ;
        RECT 164.400 957.900 166.200 958.500 ;
        RECT 173.400 957.900 186.900 958.800 ;
        RECT 151.800 955.950 155.700 957.750 ;
        RECT 164.400 956.700 175.500 957.900 ;
        RECT 153.900 955.200 155.700 955.950 ;
        RECT 173.400 955.800 175.500 956.700 ;
        RECT 177.000 955.200 180.900 957.000 ;
        RECT 186.000 956.700 186.900 957.900 ;
        RECT 153.900 954.300 167.400 955.200 ;
        RECT 178.800 954.900 180.900 955.200 ;
        RECT 185.100 954.900 186.900 956.700 ;
        RECT 189.600 958.200 190.500 959.700 ;
        RECT 189.600 956.400 194.700 958.200 ;
        RECT 196.800 958.050 198.300 960.900 ;
        RECT 196.800 955.950 198.900 958.050 ;
        RECT 166.200 953.700 167.400 954.300 ;
        RECT 200.100 953.700 201.900 954.300 ;
        RECT 161.400 952.500 163.500 952.800 ;
        RECT 166.200 952.500 201.900 953.700 ;
        RECT 151.500 951.300 163.500 952.500 ;
        RECT 202.800 951.600 203.700 968.400 ;
        RECT 151.500 950.700 153.300 951.300 ;
        RECT 161.400 950.700 163.500 951.300 ;
        RECT 166.200 950.400 183.900 951.600 ;
        RECT 148.200 949.800 150.000 950.100 ;
        RECT 166.200 949.800 167.400 950.400 ;
        RECT 148.200 948.600 167.400 949.800 ;
        RECT 181.800 949.500 183.900 950.400 ;
        RECT 187.200 950.700 203.700 951.600 ;
        RECT 187.200 949.500 189.300 950.700 ;
        RECT 148.200 948.300 150.000 948.600 ;
        RECT 143.700 946.500 147.300 947.400 ;
        RECT 146.400 945.600 147.300 946.500 ;
        RECT 106.200 939.000 108.000 945.600 ;
        RECT 109.200 939.600 111.000 945.600 ;
        RECT 112.200 942.600 114.300 944.700 ;
        RECT 115.200 942.600 117.300 944.700 ;
        RECT 118.200 942.600 120.300 944.700 ;
        RECT 112.200 939.600 114.000 942.600 ;
        RECT 115.200 939.600 117.000 942.600 ;
        RECT 118.200 939.600 120.000 942.600 ;
        RECT 121.200 939.000 123.000 945.600 ;
        RECT 124.200 939.600 126.000 945.600 ;
        RECT 127.200 939.000 129.000 945.600 ;
        RECT 130.200 939.600 132.000 945.600 ;
        RECT 133.200 939.000 135.000 945.600 ;
        RECT 136.500 939.600 138.300 945.600 ;
        RECT 139.500 939.000 141.300 945.600 ;
        RECT 143.700 939.000 145.500 945.600 ;
        RECT 146.400 944.700 148.500 945.600 ;
        RECT 146.700 939.600 148.500 944.700 ;
        RECT 149.700 939.000 151.500 945.600 ;
        RECT 152.700 939.600 154.500 948.600 ;
        RECT 164.700 945.600 166.800 947.700 ;
        RECT 172.200 947.100 175.500 949.200 ;
        RECT 155.700 939.000 157.500 945.600 ;
        RECT 159.300 942.600 161.400 944.700 ;
        RECT 162.300 942.600 164.400 944.700 ;
        RECT 159.300 939.600 161.100 942.600 ;
        RECT 162.300 939.600 164.100 942.600 ;
        RECT 165.300 939.600 167.100 945.600 ;
        RECT 168.300 939.000 170.100 945.600 ;
        RECT 172.200 939.600 174.000 947.100 ;
        RECT 178.200 945.600 180.900 949.500 ;
        RECT 193.200 948.600 198.900 949.800 ;
        RECT 190.500 947.700 192.300 948.300 ;
        RECT 184.200 946.500 192.300 947.700 ;
        RECT 184.200 945.600 186.300 946.500 ;
        RECT 193.200 945.600 194.400 948.600 ;
        RECT 197.100 948.000 198.900 948.600 ;
        RECT 202.800 947.400 203.700 950.700 ;
        RECT 199.800 946.500 203.700 947.400 ;
        RECT 205.500 971.400 207.300 974.400 ;
        RECT 208.500 971.400 210.300 975.000 ;
        RECT 205.500 958.050 207.000 971.400 ;
        RECT 212.700 968.400 214.500 974.400 ;
        RECT 218.100 968.400 219.900 975.000 ;
        RECT 223.500 968.400 225.300 974.400 ;
        RECT 227.700 971.400 229.500 974.400 ;
        RECT 230.700 971.400 232.500 974.400 ;
        RECT 233.700 971.400 235.500 974.400 ;
        RECT 236.700 971.400 238.500 975.000 ;
        RECT 227.700 969.300 229.800 971.400 ;
        RECT 230.700 969.300 232.800 971.400 ;
        RECT 233.700 969.300 235.800 971.400 ;
        RECT 241.200 970.500 243.000 974.400 ;
        RECT 244.200 971.400 246.000 975.000 ;
        RECT 247.200 971.400 249.000 974.400 ;
        RECT 250.200 971.400 252.000 974.400 ;
        RECT 253.200 971.400 255.000 974.400 ;
        RECT 256.200 971.400 258.000 974.400 ;
        RECT 237.600 969.600 239.400 970.500 ;
        RECT 236.700 968.400 239.400 969.600 ;
        RECT 241.200 968.400 243.900 970.500 ;
        RECT 247.200 969.300 249.300 971.400 ;
        RECT 250.200 969.300 252.300 971.400 ;
        RECT 253.200 969.300 255.300 971.400 ;
        RECT 256.200 969.300 258.300 971.400 ;
        RECT 260.400 969.600 262.200 974.400 ;
        RECT 260.400 968.400 264.600 969.600 ;
        RECT 265.500 968.400 267.300 975.000 ;
        RECT 270.900 968.400 272.700 974.400 ;
        RECT 212.700 964.800 213.900 968.400 ;
        RECT 223.800 967.500 225.300 968.400 ;
        RECT 232.800 967.800 234.600 968.400 ;
        RECT 236.700 967.800 237.600 968.400 ;
        RECT 216.900 966.300 225.300 967.500 ;
        RECT 230.400 966.600 237.600 967.800 ;
        RECT 252.300 966.600 258.900 968.400 ;
        RECT 216.900 965.700 218.700 966.300 ;
        RECT 227.400 964.800 229.500 965.700 ;
        RECT 212.700 963.600 229.500 964.800 ;
        RECT 230.400 963.600 231.300 966.600 ;
        RECT 235.800 963.900 237.600 964.800 ;
        RECT 245.100 964.500 246.900 966.300 ;
        RECT 263.100 965.100 264.600 968.400 ;
        RECT 238.800 963.900 240.900 964.050 ;
        RECT 205.500 955.950 207.900 958.050 ;
        RECT 199.800 945.600 201.000 946.500 ;
        RECT 205.500 945.600 207.000 955.950 ;
        RECT 212.700 947.400 213.900 963.600 ;
        RECT 230.400 961.800 232.200 963.600 ;
        RECT 235.800 963.000 240.900 963.900 ;
        RECT 238.800 961.950 240.900 963.000 ;
        RECT 245.100 963.900 247.200 964.500 ;
        RECT 245.100 962.400 262.200 963.900 ;
        RECT 263.100 963.300 270.900 965.100 ;
        RECT 260.700 960.900 267.300 962.400 ;
        RECT 215.100 959.700 259.500 960.900 ;
        RECT 215.100 958.050 216.900 959.700 ;
        RECT 214.800 955.950 216.900 958.050 ;
        RECT 220.800 957.750 222.900 958.050 ;
        RECT 233.400 957.900 235.200 958.500 ;
        RECT 242.400 957.900 255.900 958.800 ;
        RECT 220.800 955.950 224.700 957.750 ;
        RECT 233.400 956.700 244.500 957.900 ;
        RECT 222.900 955.200 224.700 955.950 ;
        RECT 242.400 955.800 244.500 956.700 ;
        RECT 246.000 955.200 249.900 957.000 ;
        RECT 255.000 956.700 255.900 957.900 ;
        RECT 222.900 954.300 236.400 955.200 ;
        RECT 247.800 954.900 249.900 955.200 ;
        RECT 254.100 954.900 255.900 956.700 ;
        RECT 258.600 958.200 259.500 959.700 ;
        RECT 258.600 956.400 263.700 958.200 ;
        RECT 265.800 958.050 267.300 960.900 ;
        RECT 265.800 955.950 267.900 958.050 ;
        RECT 235.200 953.700 236.400 954.300 ;
        RECT 269.100 953.700 270.900 954.300 ;
        RECT 230.400 952.500 232.500 952.800 ;
        RECT 235.200 952.500 270.900 953.700 ;
        RECT 220.500 951.300 232.500 952.500 ;
        RECT 271.800 951.600 272.700 968.400 ;
        RECT 220.500 950.700 222.300 951.300 ;
        RECT 230.400 950.700 232.500 951.300 ;
        RECT 235.200 950.400 252.900 951.600 ;
        RECT 217.200 949.800 219.000 950.100 ;
        RECT 235.200 949.800 236.400 950.400 ;
        RECT 217.200 948.600 236.400 949.800 ;
        RECT 250.800 949.500 252.900 950.400 ;
        RECT 256.200 950.700 272.700 951.600 ;
        RECT 256.200 949.500 258.300 950.700 ;
        RECT 217.200 948.300 219.000 948.600 ;
        RECT 212.700 946.500 216.300 947.400 ;
        RECT 215.400 945.600 216.300 946.500 ;
        RECT 175.200 939.000 177.000 945.600 ;
        RECT 178.200 939.600 180.000 945.600 ;
        RECT 181.200 942.600 183.300 944.700 ;
        RECT 184.200 942.600 186.300 944.700 ;
        RECT 187.200 942.600 189.300 944.700 ;
        RECT 181.200 939.600 183.000 942.600 ;
        RECT 184.200 939.600 186.000 942.600 ;
        RECT 187.200 939.600 189.000 942.600 ;
        RECT 190.200 939.000 192.000 945.600 ;
        RECT 193.200 939.600 195.000 945.600 ;
        RECT 196.200 939.000 198.000 945.600 ;
        RECT 199.200 939.600 201.000 945.600 ;
        RECT 202.200 939.000 204.000 945.600 ;
        RECT 205.500 939.600 207.300 945.600 ;
        RECT 208.500 939.000 210.300 945.600 ;
        RECT 212.700 939.000 214.500 945.600 ;
        RECT 215.400 944.700 217.500 945.600 ;
        RECT 215.700 939.600 217.500 944.700 ;
        RECT 218.700 939.000 220.500 945.600 ;
        RECT 221.700 939.600 223.500 948.600 ;
        RECT 233.700 945.600 235.800 947.700 ;
        RECT 241.200 947.100 244.500 949.200 ;
        RECT 224.700 939.000 226.500 945.600 ;
        RECT 228.300 942.600 230.400 944.700 ;
        RECT 231.300 942.600 233.400 944.700 ;
        RECT 228.300 939.600 230.100 942.600 ;
        RECT 231.300 939.600 233.100 942.600 ;
        RECT 234.300 939.600 236.100 945.600 ;
        RECT 237.300 939.000 239.100 945.600 ;
        RECT 241.200 939.600 243.000 947.100 ;
        RECT 247.200 945.600 249.900 949.500 ;
        RECT 262.200 948.600 267.900 949.800 ;
        RECT 259.500 947.700 261.300 948.300 ;
        RECT 253.200 946.500 261.300 947.700 ;
        RECT 253.200 945.600 255.300 946.500 ;
        RECT 262.200 945.600 263.400 948.600 ;
        RECT 266.100 948.000 267.900 948.600 ;
        RECT 271.800 947.400 272.700 950.700 ;
        RECT 268.800 946.500 272.700 947.400 ;
        RECT 274.500 971.400 276.300 974.400 ;
        RECT 277.500 971.400 279.300 975.000 ;
        RECT 274.500 958.050 276.000 971.400 ;
        RECT 281.700 968.400 283.500 974.400 ;
        RECT 287.100 968.400 288.900 975.000 ;
        RECT 292.500 968.400 294.300 974.400 ;
        RECT 296.700 971.400 298.500 974.400 ;
        RECT 299.700 971.400 301.500 974.400 ;
        RECT 302.700 971.400 304.500 974.400 ;
        RECT 305.700 971.400 307.500 975.000 ;
        RECT 296.700 969.300 298.800 971.400 ;
        RECT 299.700 969.300 301.800 971.400 ;
        RECT 302.700 969.300 304.800 971.400 ;
        RECT 310.200 970.500 312.000 974.400 ;
        RECT 313.200 971.400 315.000 975.000 ;
        RECT 316.200 971.400 318.000 974.400 ;
        RECT 319.200 971.400 321.000 974.400 ;
        RECT 322.200 971.400 324.000 974.400 ;
        RECT 325.200 971.400 327.000 974.400 ;
        RECT 306.600 969.600 308.400 970.500 ;
        RECT 305.700 968.400 308.400 969.600 ;
        RECT 310.200 968.400 312.900 970.500 ;
        RECT 316.200 969.300 318.300 971.400 ;
        RECT 319.200 969.300 321.300 971.400 ;
        RECT 322.200 969.300 324.300 971.400 ;
        RECT 325.200 969.300 327.300 971.400 ;
        RECT 329.400 969.600 331.200 974.400 ;
        RECT 329.400 968.400 333.600 969.600 ;
        RECT 334.500 968.400 336.300 975.000 ;
        RECT 339.900 968.400 341.700 974.400 ;
        RECT 281.700 964.800 282.900 968.400 ;
        RECT 292.800 967.500 294.300 968.400 ;
        RECT 301.800 967.800 303.600 968.400 ;
        RECT 305.700 967.800 306.600 968.400 ;
        RECT 285.900 966.300 294.300 967.500 ;
        RECT 299.400 966.600 306.600 967.800 ;
        RECT 321.300 966.600 327.900 968.400 ;
        RECT 285.900 965.700 287.700 966.300 ;
        RECT 296.400 964.800 298.500 965.700 ;
        RECT 281.700 963.600 298.500 964.800 ;
        RECT 299.400 963.600 300.300 966.600 ;
        RECT 304.800 963.900 306.600 964.800 ;
        RECT 314.100 964.500 315.900 966.300 ;
        RECT 332.100 965.100 333.600 968.400 ;
        RECT 307.800 963.900 309.900 964.050 ;
        RECT 274.500 955.950 276.900 958.050 ;
        RECT 268.800 945.600 270.000 946.500 ;
        RECT 274.500 945.600 276.000 955.950 ;
        RECT 281.700 947.400 282.900 963.600 ;
        RECT 299.400 961.800 301.200 963.600 ;
        RECT 304.800 963.000 309.900 963.900 ;
        RECT 307.800 961.950 309.900 963.000 ;
        RECT 314.100 963.900 316.200 964.500 ;
        RECT 314.100 962.400 331.200 963.900 ;
        RECT 332.100 963.300 339.900 965.100 ;
        RECT 329.700 960.900 336.300 962.400 ;
        RECT 284.100 959.700 328.500 960.900 ;
        RECT 284.100 958.050 285.900 959.700 ;
        RECT 283.800 955.950 285.900 958.050 ;
        RECT 289.800 957.750 291.900 958.050 ;
        RECT 302.400 957.900 304.200 958.500 ;
        RECT 311.400 957.900 324.900 958.800 ;
        RECT 289.800 955.950 293.700 957.750 ;
        RECT 302.400 956.700 313.500 957.900 ;
        RECT 291.900 955.200 293.700 955.950 ;
        RECT 311.400 955.800 313.500 956.700 ;
        RECT 315.000 955.200 318.900 957.000 ;
        RECT 324.000 956.700 324.900 957.900 ;
        RECT 291.900 954.300 305.400 955.200 ;
        RECT 316.800 954.900 318.900 955.200 ;
        RECT 323.100 954.900 324.900 956.700 ;
        RECT 327.600 958.200 328.500 959.700 ;
        RECT 327.600 956.400 332.700 958.200 ;
        RECT 334.800 958.050 336.300 960.900 ;
        RECT 334.800 955.950 336.900 958.050 ;
        RECT 304.200 953.700 305.400 954.300 ;
        RECT 338.100 953.700 339.900 954.300 ;
        RECT 299.400 952.500 301.500 952.800 ;
        RECT 304.200 952.500 339.900 953.700 ;
        RECT 289.500 951.300 301.500 952.500 ;
        RECT 340.800 951.600 341.700 968.400 ;
        RECT 289.500 950.700 291.300 951.300 ;
        RECT 299.400 950.700 301.500 951.300 ;
        RECT 304.200 950.400 321.900 951.600 ;
        RECT 286.200 949.800 288.000 950.100 ;
        RECT 304.200 949.800 305.400 950.400 ;
        RECT 286.200 948.600 305.400 949.800 ;
        RECT 319.800 949.500 321.900 950.400 ;
        RECT 325.200 950.700 341.700 951.600 ;
        RECT 325.200 949.500 327.300 950.700 ;
        RECT 286.200 948.300 288.000 948.600 ;
        RECT 281.700 946.500 285.300 947.400 ;
        RECT 284.400 945.600 285.300 946.500 ;
        RECT 244.200 939.000 246.000 945.600 ;
        RECT 247.200 939.600 249.000 945.600 ;
        RECT 250.200 942.600 252.300 944.700 ;
        RECT 253.200 942.600 255.300 944.700 ;
        RECT 256.200 942.600 258.300 944.700 ;
        RECT 250.200 939.600 252.000 942.600 ;
        RECT 253.200 939.600 255.000 942.600 ;
        RECT 256.200 939.600 258.000 942.600 ;
        RECT 259.200 939.000 261.000 945.600 ;
        RECT 262.200 939.600 264.000 945.600 ;
        RECT 265.200 939.000 267.000 945.600 ;
        RECT 268.200 939.600 270.000 945.600 ;
        RECT 271.200 939.000 273.000 945.600 ;
        RECT 274.500 939.600 276.300 945.600 ;
        RECT 277.500 939.000 279.300 945.600 ;
        RECT 281.700 939.000 283.500 945.600 ;
        RECT 284.400 944.700 286.500 945.600 ;
        RECT 284.700 939.600 286.500 944.700 ;
        RECT 287.700 939.000 289.500 945.600 ;
        RECT 290.700 939.600 292.500 948.600 ;
        RECT 302.700 945.600 304.800 947.700 ;
        RECT 310.200 947.100 313.500 949.200 ;
        RECT 293.700 939.000 295.500 945.600 ;
        RECT 297.300 942.600 299.400 944.700 ;
        RECT 300.300 942.600 302.400 944.700 ;
        RECT 297.300 939.600 299.100 942.600 ;
        RECT 300.300 939.600 302.100 942.600 ;
        RECT 303.300 939.600 305.100 945.600 ;
        RECT 306.300 939.000 308.100 945.600 ;
        RECT 310.200 939.600 312.000 947.100 ;
        RECT 316.200 945.600 318.900 949.500 ;
        RECT 331.200 948.600 336.900 949.800 ;
        RECT 328.500 947.700 330.300 948.300 ;
        RECT 322.200 946.500 330.300 947.700 ;
        RECT 322.200 945.600 324.300 946.500 ;
        RECT 331.200 945.600 332.400 948.600 ;
        RECT 335.100 948.000 336.900 948.600 ;
        RECT 340.800 947.400 341.700 950.700 ;
        RECT 337.800 946.500 341.700 947.400 ;
        RECT 343.500 971.400 345.300 974.400 ;
        RECT 346.500 971.400 348.300 975.000 ;
        RECT 343.500 958.050 345.000 971.400 ;
        RECT 365.100 968.400 366.900 974.400 ;
        RECT 365.700 966.300 366.900 968.400 ;
        RECT 368.100 969.300 369.900 974.400 ;
        RECT 371.100 970.200 372.900 975.000 ;
        RECT 374.100 969.300 375.900 974.400 ;
        RECT 368.100 967.950 375.900 969.300 ;
        RECT 365.700 965.400 369.300 966.300 ;
        RECT 394.500 966.000 396.300 974.400 ;
        RECT 365.100 961.050 366.900 962.850 ;
        RECT 368.100 961.050 369.300 965.400 ;
        RECT 393.000 964.800 396.300 966.000 ;
        RECT 401.100 965.400 402.900 975.000 ;
        RECT 419.700 967.200 421.500 974.400 ;
        RECT 424.800 968.400 426.600 975.000 ;
        RECT 419.700 966.300 423.900 967.200 ;
        RECT 371.100 961.050 372.900 962.850 ;
        RECT 393.000 961.050 393.900 964.800 ;
        RECT 395.100 961.050 396.900 962.850 ;
        RECT 401.100 961.050 402.900 962.850 ;
        RECT 419.100 961.050 420.900 962.850 ;
        RECT 422.700 961.050 423.900 966.300 ;
        RECT 445.500 966.000 447.300 974.400 ;
        RECT 444.000 964.800 447.300 966.000 ;
        RECT 452.100 965.400 453.900 975.000 ;
        RECT 470.100 968.400 471.900 974.400 ;
        RECT 470.700 966.300 471.900 968.400 ;
        RECT 473.100 969.300 474.900 974.400 ;
        RECT 476.100 970.200 477.900 975.000 ;
        RECT 479.100 969.300 480.900 974.400 ;
        RECT 497.100 971.400 498.900 974.400 ;
        RECT 500.100 971.400 501.900 975.000 ;
        RECT 518.100 971.400 519.900 974.400 ;
        RECT 521.100 971.400 522.900 975.000 ;
        RECT 473.100 967.950 480.900 969.300 ;
        RECT 470.700 965.400 474.300 966.300 ;
        RECT 424.950 961.050 426.750 962.850 ;
        RECT 444.000 961.050 444.900 964.800 ;
        RECT 446.100 961.050 447.900 962.850 ;
        RECT 452.100 961.050 453.900 962.850 ;
        RECT 470.100 961.050 471.900 962.850 ;
        RECT 473.100 961.050 474.300 965.400 ;
        RECT 476.100 961.050 477.900 962.850 ;
        RECT 497.700 961.050 498.900 971.400 ;
        RECT 518.700 961.050 519.900 971.400 ;
        RECT 539.400 968.400 541.200 975.000 ;
        RECT 544.500 967.200 546.300 974.400 ;
        RECT 561.000 968.400 562.800 975.000 ;
        RECT 565.500 969.600 567.300 974.400 ;
        RECT 568.500 971.400 570.300 975.000 ;
        RECT 587.100 971.400 588.900 975.000 ;
        RECT 590.100 971.400 591.900 974.400 ;
        RECT 593.100 971.400 594.900 975.000 ;
        RECT 565.500 968.400 570.600 969.600 ;
        RECT 542.100 966.300 546.300 967.200 ;
        RECT 539.250 961.050 541.050 962.850 ;
        RECT 542.100 961.050 543.300 966.300 ;
        RECT 545.100 961.050 546.900 962.850 ;
        RECT 560.100 961.050 561.900 962.850 ;
        RECT 566.250 961.050 568.050 962.850 ;
        RECT 569.700 961.050 570.600 968.400 ;
        RECT 590.400 961.050 591.300 971.400 ;
        RECT 611.100 968.400 612.900 974.400 ;
        RECT 611.700 966.300 612.900 968.400 ;
        RECT 614.100 969.300 615.900 974.400 ;
        RECT 617.100 970.200 618.900 975.000 ;
        RECT 620.100 969.300 621.900 974.400 ;
        RECT 614.100 967.950 621.900 969.300 ;
        RECT 638.400 968.400 640.200 975.000 ;
        RECT 643.500 967.200 645.300 974.400 ;
        RECT 641.100 966.300 645.300 967.200 ;
        RECT 611.700 965.400 615.300 966.300 ;
        RECT 611.100 961.050 612.900 962.850 ;
        RECT 614.100 961.050 615.300 965.400 ;
        RECT 617.100 961.050 618.900 962.850 ;
        RECT 638.250 961.050 640.050 962.850 ;
        RECT 641.100 961.050 642.300 966.300 ;
        RECT 662.100 965.400 663.900 975.000 ;
        RECT 668.700 966.000 670.500 974.400 ;
        RECT 689.700 967.200 691.500 974.400 ;
        RECT 694.800 968.400 696.600 975.000 ;
        RECT 713.100 971.400 714.900 975.000 ;
        RECT 716.100 971.400 717.900 974.400 ;
        RECT 689.700 966.300 693.900 967.200 ;
        RECT 668.700 964.800 672.000 966.000 ;
        RECT 644.100 961.050 645.900 962.850 ;
        RECT 662.100 961.050 663.900 962.850 ;
        RECT 668.100 961.050 669.900 962.850 ;
        RECT 671.100 961.050 672.000 964.800 ;
        RECT 689.100 961.050 690.900 962.850 ;
        RECT 692.700 961.050 693.900 966.300 ;
        RECT 694.950 961.050 696.750 962.850 ;
        RECT 716.100 961.050 717.300 971.400 ;
        RECT 734.100 968.400 735.900 974.400 ;
        RECT 734.700 966.300 735.900 968.400 ;
        RECT 737.100 969.300 738.900 974.400 ;
        RECT 740.100 970.200 741.900 975.000 ;
        RECT 743.100 969.300 744.900 974.400 ;
        RECT 761.100 971.400 762.900 975.000 ;
        RECT 764.100 971.400 765.900 974.400 ;
        RECT 767.100 971.400 768.900 975.000 ;
        RECT 737.100 967.950 744.900 969.300 ;
        RECT 734.700 965.400 738.300 966.300 ;
        RECT 734.100 961.050 735.900 962.850 ;
        RECT 737.100 961.050 738.300 965.400 ;
        RECT 740.100 961.050 741.900 962.850 ;
        RECT 764.700 961.050 765.600 971.400 ;
        RECT 785.700 968.400 787.500 975.000 ;
        RECT 790.200 968.400 792.000 974.400 ;
        RECT 794.700 968.400 796.500 975.000 ;
        RECT 816.600 970.200 818.400 974.400 ;
        RECT 815.700 968.400 818.400 970.200 ;
        RECT 819.600 968.400 821.400 975.000 ;
        RECT 785.250 961.050 787.050 962.850 ;
        RECT 791.100 961.050 792.300 968.400 ;
        RECT 797.100 961.050 798.900 962.850 ;
        RECT 815.700 961.050 816.600 968.400 ;
        RECT 817.500 966.600 819.300 967.500 ;
        RECT 824.100 966.600 825.900 974.400 ;
        RECT 817.500 965.700 825.900 966.600 ;
        RECT 842.700 967.200 844.500 974.400 ;
        RECT 847.800 968.400 849.600 975.000 ;
        RECT 866.400 968.400 868.200 975.000 ;
        RECT 871.500 967.200 873.300 974.400 ;
        RECT 890.100 968.400 891.900 974.400 ;
        RECT 842.700 966.300 846.900 967.200 ;
        RECT 364.950 958.950 367.050 961.050 ;
        RECT 367.950 958.950 370.050 961.050 ;
        RECT 370.950 958.950 373.050 961.050 ;
        RECT 373.950 958.950 376.050 961.050 ;
        RECT 391.950 958.950 394.050 961.050 ;
        RECT 394.950 958.950 397.050 961.050 ;
        RECT 397.950 958.950 400.050 961.050 ;
        RECT 400.950 958.950 403.050 961.050 ;
        RECT 418.950 958.950 421.050 961.050 ;
        RECT 421.950 958.950 424.050 961.050 ;
        RECT 424.950 958.950 427.050 961.050 ;
        RECT 442.950 958.950 445.050 961.050 ;
        RECT 445.950 958.950 448.050 961.050 ;
        RECT 448.950 958.950 451.050 961.050 ;
        RECT 451.950 958.950 454.050 961.050 ;
        RECT 469.950 958.950 472.050 961.050 ;
        RECT 472.950 958.950 475.050 961.050 ;
        RECT 475.950 958.950 478.050 961.050 ;
        RECT 478.950 958.950 481.050 961.050 ;
        RECT 496.950 958.950 499.050 961.050 ;
        RECT 499.950 958.950 502.050 961.050 ;
        RECT 517.950 958.950 520.050 961.050 ;
        RECT 520.950 958.950 523.050 961.050 ;
        RECT 538.950 958.950 541.050 961.050 ;
        RECT 541.950 958.950 544.050 961.050 ;
        RECT 544.950 958.950 547.050 961.050 ;
        RECT 559.950 958.950 562.050 961.050 ;
        RECT 562.950 958.950 565.050 961.050 ;
        RECT 565.950 958.950 568.050 961.050 ;
        RECT 568.950 958.950 571.050 961.050 ;
        RECT 586.950 958.950 589.050 961.050 ;
        RECT 589.950 958.950 592.050 961.050 ;
        RECT 592.950 958.950 595.050 961.050 ;
        RECT 610.950 958.950 613.050 961.050 ;
        RECT 613.950 958.950 616.050 961.050 ;
        RECT 616.950 958.950 619.050 961.050 ;
        RECT 619.950 958.950 622.050 961.050 ;
        RECT 637.950 958.950 640.050 961.050 ;
        RECT 640.950 958.950 643.050 961.050 ;
        RECT 643.950 958.950 646.050 961.050 ;
        RECT 661.950 958.950 664.050 961.050 ;
        RECT 664.950 958.950 667.050 961.050 ;
        RECT 667.950 958.950 670.050 961.050 ;
        RECT 670.950 958.950 673.050 961.050 ;
        RECT 688.950 958.950 691.050 961.050 ;
        RECT 691.950 958.950 694.050 961.050 ;
        RECT 694.950 958.950 697.050 961.050 ;
        RECT 712.950 958.950 715.050 961.050 ;
        RECT 715.950 958.950 718.050 961.050 ;
        RECT 733.950 958.950 736.050 961.050 ;
        RECT 736.950 958.950 739.050 961.050 ;
        RECT 739.950 958.950 742.050 961.050 ;
        RECT 742.950 958.950 745.050 961.050 ;
        RECT 760.950 958.950 763.050 961.050 ;
        RECT 763.950 958.950 766.050 961.050 ;
        RECT 766.950 958.950 769.050 961.050 ;
        RECT 784.950 958.950 787.050 961.050 ;
        RECT 787.950 958.950 790.050 961.050 ;
        RECT 790.950 958.950 793.050 961.050 ;
        RECT 793.950 958.950 796.050 961.050 ;
        RECT 796.950 958.950 799.050 961.050 ;
        RECT 815.100 958.950 817.200 961.050 ;
        RECT 818.400 958.950 820.500 961.050 ;
        RECT 343.500 955.950 345.900 958.050 ;
        RECT 337.800 945.600 339.000 946.500 ;
        RECT 343.500 945.600 345.000 955.950 ;
        RECT 368.100 951.600 369.300 958.950 ;
        RECT 374.100 957.150 375.900 958.950 ;
        RECT 368.100 950.100 370.500 951.600 ;
        RECT 366.000 947.100 367.800 948.900 ;
        RECT 313.200 939.000 315.000 945.600 ;
        RECT 316.200 939.600 318.000 945.600 ;
        RECT 319.200 942.600 321.300 944.700 ;
        RECT 322.200 942.600 324.300 944.700 ;
        RECT 325.200 942.600 327.300 944.700 ;
        RECT 319.200 939.600 321.000 942.600 ;
        RECT 322.200 939.600 324.000 942.600 ;
        RECT 325.200 939.600 327.000 942.600 ;
        RECT 328.200 939.000 330.000 945.600 ;
        RECT 331.200 939.600 333.000 945.600 ;
        RECT 334.200 939.000 336.000 945.600 ;
        RECT 337.200 939.600 339.000 945.600 ;
        RECT 340.200 939.000 342.000 945.600 ;
        RECT 343.500 939.600 345.300 945.600 ;
        RECT 346.500 939.000 348.300 945.600 ;
        RECT 365.700 939.000 367.500 945.600 ;
        RECT 368.700 939.600 370.500 950.100 ;
        RECT 373.800 939.000 375.600 951.600 ;
        RECT 393.000 946.800 393.900 958.950 ;
        RECT 398.100 957.150 399.900 958.950 ;
        RECT 393.000 945.900 399.600 946.800 ;
        RECT 393.000 945.600 393.900 945.900 ;
        RECT 392.100 939.600 393.900 945.600 ;
        RECT 398.100 945.600 399.600 945.900 ;
        RECT 422.700 945.600 423.900 958.950 ;
        RECT 444.000 946.800 444.900 958.950 ;
        RECT 449.100 957.150 450.900 958.950 ;
        RECT 473.100 951.600 474.300 958.950 ;
        RECT 479.100 957.150 480.900 958.950 ;
        RECT 473.100 950.100 475.500 951.600 ;
        RECT 471.000 947.100 472.800 948.900 ;
        RECT 444.000 945.900 450.600 946.800 ;
        RECT 444.000 945.600 444.900 945.900 ;
        RECT 395.100 939.000 396.900 945.000 ;
        RECT 398.100 939.600 399.900 945.600 ;
        RECT 401.100 939.000 402.900 945.600 ;
        RECT 419.100 939.000 420.900 945.600 ;
        RECT 422.100 939.600 423.900 945.600 ;
        RECT 425.100 939.000 426.900 945.600 ;
        RECT 443.100 939.600 444.900 945.600 ;
        RECT 449.100 945.600 450.600 945.900 ;
        RECT 446.100 939.000 447.900 945.000 ;
        RECT 449.100 939.600 450.900 945.600 ;
        RECT 452.100 939.000 453.900 945.600 ;
        RECT 470.700 939.000 472.500 945.600 ;
        RECT 473.700 939.600 475.500 950.100 ;
        RECT 478.800 939.000 480.600 951.600 ;
        RECT 497.700 945.600 498.900 958.950 ;
        RECT 500.100 957.150 501.900 958.950 ;
        RECT 518.700 945.600 519.900 958.950 ;
        RECT 521.100 957.150 522.900 958.950 ;
        RECT 542.100 945.600 543.300 958.950 ;
        RECT 563.250 957.150 565.050 958.950 ;
        RECT 569.700 951.600 570.600 958.950 ;
        RECT 587.250 957.150 589.050 958.950 ;
        RECT 590.400 951.600 591.300 958.950 ;
        RECT 593.100 957.150 594.900 958.950 ;
        RECT 595.950 954.450 598.050 955.050 ;
        RECT 610.950 954.450 613.050 955.050 ;
        RECT 595.950 953.550 613.050 954.450 ;
        RECT 595.950 952.950 598.050 953.550 ;
        RECT 610.950 952.950 613.050 953.550 ;
        RECT 614.100 951.600 615.300 958.950 ;
        RECT 620.100 957.150 621.900 958.950 ;
        RECT 560.100 950.700 567.900 951.600 ;
        RECT 497.100 939.600 498.900 945.600 ;
        RECT 500.100 939.000 501.900 945.600 ;
        RECT 518.100 939.600 519.900 945.600 ;
        RECT 521.100 939.000 522.900 945.600 ;
        RECT 539.100 939.000 540.900 945.600 ;
        RECT 542.100 939.600 543.900 945.600 ;
        RECT 545.100 939.000 546.900 945.600 ;
        RECT 560.100 939.600 561.900 950.700 ;
        RECT 563.100 939.000 564.900 949.800 ;
        RECT 566.100 939.600 567.900 950.700 ;
        RECT 569.100 939.600 570.900 951.600 ;
        RECT 587.100 939.000 588.900 951.600 ;
        RECT 590.400 950.400 594.000 951.600 ;
        RECT 592.200 939.600 594.000 950.400 ;
        RECT 614.100 950.100 616.500 951.600 ;
        RECT 612.000 947.100 613.800 948.900 ;
        RECT 611.700 939.000 613.500 945.600 ;
        RECT 614.700 939.600 616.500 950.100 ;
        RECT 619.800 939.000 621.600 951.600 ;
        RECT 641.100 945.600 642.300 958.950 ;
        RECT 665.100 957.150 666.900 958.950 ;
        RECT 671.100 946.800 672.000 958.950 ;
        RECT 665.400 945.900 672.000 946.800 ;
        RECT 665.400 945.600 666.900 945.900 ;
        RECT 638.100 939.000 639.900 945.600 ;
        RECT 641.100 939.600 642.900 945.600 ;
        RECT 644.100 939.000 645.900 945.600 ;
        RECT 662.100 939.000 663.900 945.600 ;
        RECT 665.100 939.600 666.900 945.600 ;
        RECT 671.100 945.600 672.000 945.900 ;
        RECT 692.700 945.600 693.900 958.950 ;
        RECT 713.100 957.150 714.900 958.950 ;
        RECT 716.100 945.600 717.300 958.950 ;
        RECT 737.100 951.600 738.300 958.950 ;
        RECT 743.100 957.150 744.900 958.950 ;
        RECT 761.100 957.150 762.900 958.950 ;
        RECT 739.950 954.450 742.050 955.050 ;
        RECT 748.950 954.450 751.050 955.050 ;
        RECT 739.950 953.550 751.050 954.450 ;
        RECT 739.950 952.950 742.050 953.550 ;
        RECT 748.950 952.950 751.050 953.550 ;
        RECT 764.700 951.600 765.600 958.950 ;
        RECT 766.950 957.150 768.750 958.950 ;
        RECT 788.250 957.150 790.050 958.950 ;
        RECT 791.100 953.400 792.000 958.950 ;
        RECT 794.100 957.150 795.900 958.950 ;
        RECT 791.100 952.500 795.900 953.400 ;
        RECT 737.100 950.100 739.500 951.600 ;
        RECT 735.000 947.100 736.800 948.900 ;
        RECT 668.100 939.000 669.900 945.000 ;
        RECT 671.100 939.600 672.900 945.600 ;
        RECT 689.100 939.000 690.900 945.600 ;
        RECT 692.100 939.600 693.900 945.600 ;
        RECT 695.100 939.000 696.900 945.600 ;
        RECT 713.100 939.000 714.900 945.600 ;
        RECT 716.100 939.600 717.900 945.600 ;
        RECT 734.700 939.000 736.500 945.600 ;
        RECT 737.700 939.600 739.500 950.100 ;
        RECT 742.800 939.000 744.600 951.600 ;
        RECT 762.000 950.400 765.600 951.600 ;
        RECT 762.000 939.600 763.800 950.400 ;
        RECT 767.100 939.000 768.900 951.600 ;
        RECT 785.100 950.400 792.900 951.300 ;
        RECT 785.100 939.600 786.900 950.400 ;
        RECT 788.100 939.000 789.900 949.500 ;
        RECT 791.100 940.500 792.900 950.400 ;
        RECT 794.100 941.400 795.900 952.500 ;
        RECT 815.700 951.600 816.600 958.950 ;
        RECT 819.000 957.150 820.800 958.950 ;
        RECT 797.100 940.500 798.900 951.600 ;
        RECT 791.100 939.600 798.900 940.500 ;
        RECT 815.100 939.600 816.900 951.600 ;
        RECT 818.100 939.000 819.900 951.000 ;
        RECT 822.000 945.600 822.900 965.700 ;
        RECT 823.950 961.050 825.750 962.850 ;
        RECT 842.100 961.050 843.900 962.850 ;
        RECT 845.700 961.050 846.900 966.300 ;
        RECT 869.100 966.300 873.300 967.200 ;
        RECT 890.700 966.300 891.900 968.400 ;
        RECT 893.100 969.300 894.900 974.400 ;
        RECT 896.100 970.200 897.900 975.000 ;
        RECT 899.100 969.300 900.900 974.400 ;
        RECT 893.100 967.950 900.900 969.300 ;
        RECT 917.700 967.200 919.500 974.400 ;
        RECT 922.800 968.400 924.600 975.000 ;
        RECT 917.700 966.300 921.900 967.200 ;
        RECT 847.950 961.050 849.750 962.850 ;
        RECT 866.250 961.050 868.050 962.850 ;
        RECT 869.100 961.050 870.300 966.300 ;
        RECT 890.700 965.400 894.300 966.300 ;
        RECT 872.100 961.050 873.900 962.850 ;
        RECT 890.100 961.050 891.900 962.850 ;
        RECT 893.100 961.050 894.300 965.400 ;
        RECT 896.100 961.050 897.900 962.850 ;
        RECT 917.100 961.050 918.900 962.850 ;
        RECT 920.700 961.050 921.900 966.300 ;
        RECT 941.100 965.400 942.900 975.000 ;
        RECT 947.700 966.000 949.500 974.400 ;
        RECT 968.100 968.400 969.900 975.000 ;
        RECT 971.100 968.400 972.900 974.400 ;
        RECT 997.200 971.400 999.900 974.400 ;
        RECT 1001.100 971.400 1002.900 975.000 ;
        RECT 1004.100 971.400 1005.900 974.400 ;
        RECT 1007.100 971.400 1009.200 975.000 ;
        RECT 997.200 970.500 998.100 971.400 ;
        RECT 1004.400 970.500 1005.300 971.400 ;
        RECT 992.700 969.600 1005.300 970.500 ;
        RECT 947.700 964.800 951.000 966.000 ;
        RECT 922.950 961.050 924.750 962.850 ;
        RECT 941.100 961.050 942.900 962.850 ;
        RECT 947.100 961.050 948.900 962.850 ;
        RECT 950.100 961.050 951.000 964.800 ;
        RECT 968.100 961.050 969.900 962.850 ;
        RECT 971.100 961.050 972.300 968.400 ;
        RECT 973.950 963.450 976.050 964.050 ;
        RECT 988.950 963.450 991.050 964.050 ;
        RECT 973.950 962.550 991.050 963.450 ;
        RECT 973.950 961.950 976.050 962.550 ;
        RECT 988.950 961.950 991.050 962.550 ;
        RECT 992.700 961.050 993.900 969.600 ;
        RECT 1028.700 967.200 1030.500 974.400 ;
        RECT 1033.800 968.400 1035.600 975.000 ;
        RECT 1028.700 966.300 1032.900 967.200 ;
        RECT 1001.250 961.050 1003.050 962.850 ;
        RECT 1028.100 961.050 1029.900 962.850 ;
        RECT 1031.700 961.050 1032.900 966.300 ;
        RECT 1033.950 961.050 1035.750 962.850 ;
        RECT 823.800 958.950 825.900 961.050 ;
        RECT 841.950 958.950 844.050 961.050 ;
        RECT 844.950 958.950 847.050 961.050 ;
        RECT 847.950 958.950 850.050 961.050 ;
        RECT 865.950 958.950 868.050 961.050 ;
        RECT 868.950 958.950 871.050 961.050 ;
        RECT 871.950 958.950 874.050 961.050 ;
        RECT 889.950 958.950 892.050 961.050 ;
        RECT 892.950 958.950 895.050 961.050 ;
        RECT 895.950 958.950 898.050 961.050 ;
        RECT 898.950 958.950 901.050 961.050 ;
        RECT 916.950 958.950 919.050 961.050 ;
        RECT 919.950 958.950 922.050 961.050 ;
        RECT 922.950 958.950 925.050 961.050 ;
        RECT 940.950 958.950 943.050 961.050 ;
        RECT 943.950 958.950 946.050 961.050 ;
        RECT 946.950 958.950 949.050 961.050 ;
        RECT 949.950 958.950 952.050 961.050 ;
        RECT 967.950 958.950 970.050 961.050 ;
        RECT 970.950 958.950 973.050 961.050 ;
        RECT 992.400 958.950 994.500 961.050 ;
        RECT 997.950 958.950 1000.050 961.050 ;
        RECT 1000.950 958.950 1003.050 961.050 ;
        RECT 1007.100 958.950 1009.200 961.050 ;
        RECT 1027.950 958.950 1030.050 961.050 ;
        RECT 1030.950 958.950 1033.050 961.050 ;
        RECT 1033.950 958.950 1036.050 961.050 ;
        RECT 845.700 945.600 846.900 958.950 ;
        RECT 869.100 945.600 870.300 958.950 ;
        RECT 893.100 951.600 894.300 958.950 ;
        RECT 899.100 957.150 900.900 958.950 ;
        RECT 893.100 950.100 895.500 951.600 ;
        RECT 891.000 947.100 892.800 948.900 ;
        RECT 821.100 939.600 822.900 945.600 ;
        RECT 824.100 939.000 825.900 945.600 ;
        RECT 842.100 939.000 843.900 945.600 ;
        RECT 845.100 939.600 846.900 945.600 ;
        RECT 848.100 939.000 849.900 945.600 ;
        RECT 866.100 939.000 867.900 945.600 ;
        RECT 869.100 939.600 870.900 945.600 ;
        RECT 872.100 939.000 873.900 945.600 ;
        RECT 890.700 939.000 892.500 945.600 ;
        RECT 893.700 939.600 895.500 950.100 ;
        RECT 898.800 939.000 900.600 951.600 ;
        RECT 920.700 945.600 921.900 958.950 ;
        RECT 944.100 957.150 945.900 958.950 ;
        RECT 950.100 946.800 951.000 958.950 ;
        RECT 955.950 954.450 958.050 955.050 ;
        RECT 967.950 954.450 970.050 955.050 ;
        RECT 955.950 953.550 970.050 954.450 ;
        RECT 955.950 952.950 958.050 953.550 ;
        RECT 967.950 952.950 970.050 953.550 ;
        RECT 971.100 951.600 972.300 958.950 ;
        RECT 944.400 945.900 951.000 946.800 ;
        RECT 944.400 945.600 945.900 945.900 ;
        RECT 917.100 939.000 918.900 945.600 ;
        RECT 920.100 939.600 921.900 945.600 ;
        RECT 923.100 939.000 924.900 945.600 ;
        RECT 941.100 939.000 942.900 945.600 ;
        RECT 944.100 939.600 945.900 945.600 ;
        RECT 950.100 945.600 951.000 945.900 ;
        RECT 947.100 939.000 948.900 945.000 ;
        RECT 950.100 939.600 951.900 945.600 ;
        RECT 968.100 939.000 969.900 951.600 ;
        RECT 971.100 939.600 972.900 951.600 ;
        RECT 989.100 940.500 990.900 949.800 ;
        RECT 992.700 949.200 993.900 958.950 ;
        RECT 997.950 957.150 999.750 958.950 ;
        RECT 1007.100 957.150 1008.900 958.950 ;
        RECT 992.100 941.400 993.900 949.200 ;
        RECT 995.100 949.200 1002.900 950.100 ;
        RECT 995.100 940.500 996.900 949.200 ;
        RECT 989.100 939.600 996.900 940.500 ;
        RECT 998.100 940.500 999.900 948.300 ;
        RECT 1001.100 941.400 1002.900 949.200 ;
        RECT 1004.100 949.500 1011.900 950.400 ;
        RECT 1004.100 940.500 1005.900 949.500 ;
        RECT 998.100 939.600 1005.900 940.500 ;
        RECT 1007.100 939.000 1008.900 948.600 ;
        RECT 1010.100 939.600 1011.900 949.500 ;
        RECT 1031.700 945.600 1032.900 958.950 ;
        RECT 1028.100 939.000 1029.900 945.600 ;
        RECT 1031.100 939.600 1032.900 945.600 ;
        RECT 1034.100 939.000 1035.900 945.600 ;
        RECT 17.100 923.400 18.900 936.000 ;
        RECT 20.100 922.500 21.900 935.400 ;
        RECT 23.100 923.400 24.900 936.000 ;
        RECT 26.100 923.400 27.900 935.400 ;
        RECT 29.100 923.400 30.900 936.000 ;
        RECT 47.100 929.400 48.900 935.400 ;
        RECT 26.100 922.500 27.300 923.400 ;
        RECT 20.100 921.600 27.300 922.500 ;
        RECT 47.100 922.500 48.300 929.400 ;
        RECT 50.100 925.200 51.900 936.000 ;
        RECT 53.100 923.400 54.900 935.400 ;
        RECT 47.100 921.600 52.800 922.500 ;
        RECT 20.100 916.050 21.900 917.850 ;
        RECT 26.100 916.050 27.300 921.600 ;
        RECT 51.000 920.700 52.800 921.600 ;
        RECT 47.400 916.050 49.200 917.850 ;
        RECT 20.100 913.950 22.200 916.050 ;
        RECT 26.100 913.950 28.200 916.050 ;
        RECT 47.400 913.950 49.500 916.050 ;
        RECT 26.100 908.700 27.300 913.950 ;
        RECT 20.100 907.500 27.300 908.700 ;
        RECT 51.000 909.300 51.900 920.700 ;
        RECT 53.700 916.050 54.900 923.400 ;
        RECT 52.800 913.950 54.900 916.050 ;
        RECT 51.000 908.400 52.800 909.300 ;
        RECT 20.100 906.600 21.300 907.500 ;
        RECT 26.100 906.600 27.300 907.500 ;
        RECT 47.100 907.500 52.800 908.400 ;
        RECT 17.100 900.000 18.900 906.600 ;
        RECT 20.100 900.600 21.900 906.600 ;
        RECT 23.100 900.000 24.900 906.600 ;
        RECT 26.100 900.600 27.900 906.600 ;
        RECT 29.100 900.000 30.900 906.600 ;
        RECT 47.100 903.600 48.300 907.500 ;
        RECT 53.700 906.600 54.900 913.950 ;
        RECT 47.100 900.600 48.900 903.600 ;
        RECT 50.100 900.000 51.900 906.600 ;
        RECT 53.100 900.600 54.900 906.600 ;
        RECT 71.100 923.400 72.900 935.400 ;
        RECT 74.100 925.200 75.900 936.000 ;
        RECT 77.100 929.400 78.900 935.400 ;
        RECT 71.100 916.050 72.300 923.400 ;
        RECT 77.700 922.500 78.900 929.400 ;
        RECT 95.100 923.400 96.900 936.000 ;
        RECT 100.200 924.600 102.000 935.400 ;
        RECT 119.700 929.400 121.500 936.000 ;
        RECT 120.000 926.100 121.800 927.900 ;
        RECT 122.700 924.900 124.500 935.400 ;
        RECT 98.400 923.400 102.000 924.600 ;
        RECT 122.100 923.400 124.500 924.900 ;
        RECT 127.800 923.400 129.600 936.000 ;
        RECT 146.700 929.400 148.500 936.000 ;
        RECT 147.000 926.100 148.800 927.900 ;
        RECT 149.700 924.900 151.500 935.400 ;
        RECT 149.100 923.400 151.500 924.900 ;
        RECT 154.800 923.400 156.600 936.000 ;
        RECT 158.700 929.400 160.500 936.000 ;
        RECT 161.700 930.300 163.500 935.400 ;
        RECT 161.400 929.400 163.500 930.300 ;
        RECT 164.700 929.400 166.500 936.000 ;
        RECT 161.400 928.500 162.300 929.400 ;
        RECT 158.700 927.600 162.300 928.500 ;
        RECT 73.200 921.600 78.900 922.500 ;
        RECT 73.200 920.700 75.000 921.600 ;
        RECT 71.100 913.950 73.200 916.050 ;
        RECT 71.100 906.600 72.300 913.950 ;
        RECT 74.100 909.300 75.000 920.700 ;
        RECT 76.800 916.050 78.600 917.850 ;
        RECT 95.250 916.050 97.050 917.850 ;
        RECT 98.400 916.050 99.300 923.400 ;
        RECT 101.100 916.050 102.900 917.850 ;
        RECT 122.100 916.050 123.300 923.400 ;
        RECT 128.100 916.050 129.900 917.850 ;
        RECT 149.100 916.050 150.300 923.400 ;
        RECT 155.100 916.050 156.900 917.850 ;
        RECT 76.500 913.950 78.600 916.050 ;
        RECT 94.950 913.950 97.050 916.050 ;
        RECT 97.950 913.950 100.050 916.050 ;
        RECT 100.950 913.950 103.050 916.050 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 121.950 913.950 124.050 916.050 ;
        RECT 124.950 913.950 127.050 916.050 ;
        RECT 127.950 913.950 130.050 916.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 148.950 913.950 151.050 916.050 ;
        RECT 151.950 913.950 154.050 916.050 ;
        RECT 154.950 913.950 157.050 916.050 ;
        RECT 73.200 908.400 75.000 909.300 ;
        RECT 73.200 907.500 78.900 908.400 ;
        RECT 71.100 900.600 72.900 906.600 ;
        RECT 74.100 900.000 75.900 906.600 ;
        RECT 77.700 903.600 78.900 907.500 ;
        RECT 98.400 903.600 99.300 913.950 ;
        RECT 119.100 912.150 120.900 913.950 ;
        RECT 122.100 909.600 123.300 913.950 ;
        RECT 125.100 912.150 126.900 913.950 ;
        RECT 146.100 912.150 147.900 913.950 ;
        RECT 149.100 909.600 150.300 913.950 ;
        RECT 152.100 912.150 153.900 913.950 ;
        RECT 119.700 908.700 123.300 909.600 ;
        RECT 146.700 908.700 150.300 909.600 ;
        RECT 158.700 911.400 159.900 927.600 ;
        RECT 163.200 926.400 165.000 926.700 ;
        RECT 167.700 926.400 169.500 935.400 ;
        RECT 170.700 929.400 172.500 936.000 ;
        RECT 174.300 932.400 176.100 935.400 ;
        RECT 177.300 932.400 179.100 935.400 ;
        RECT 174.300 930.300 176.400 932.400 ;
        RECT 177.300 930.300 179.400 932.400 ;
        RECT 180.300 929.400 182.100 935.400 ;
        RECT 183.300 929.400 185.100 936.000 ;
        RECT 179.700 927.300 181.800 929.400 ;
        RECT 187.200 927.900 189.000 935.400 ;
        RECT 190.200 929.400 192.000 936.000 ;
        RECT 193.200 929.400 195.000 935.400 ;
        RECT 196.200 932.400 198.000 935.400 ;
        RECT 199.200 932.400 201.000 935.400 ;
        RECT 202.200 932.400 204.000 935.400 ;
        RECT 196.200 930.300 198.300 932.400 ;
        RECT 199.200 930.300 201.300 932.400 ;
        RECT 202.200 930.300 204.300 932.400 ;
        RECT 205.200 929.400 207.000 936.000 ;
        RECT 208.200 929.400 210.000 935.400 ;
        RECT 211.200 929.400 213.000 936.000 ;
        RECT 214.200 929.400 216.000 935.400 ;
        RECT 217.200 929.400 219.000 936.000 ;
        RECT 220.500 929.400 222.300 935.400 ;
        RECT 223.500 929.400 225.300 936.000 ;
        RECT 163.200 925.200 182.400 926.400 ;
        RECT 187.200 925.800 190.500 927.900 ;
        RECT 193.200 925.500 195.900 929.400 ;
        RECT 199.200 928.500 201.300 929.400 ;
        RECT 199.200 927.300 207.300 928.500 ;
        RECT 205.500 926.700 207.300 927.300 ;
        RECT 208.200 926.400 209.400 929.400 ;
        RECT 214.800 928.500 216.000 929.400 ;
        RECT 214.800 927.600 218.700 928.500 ;
        RECT 212.100 926.400 213.900 927.000 ;
        RECT 163.200 924.900 165.000 925.200 ;
        RECT 181.200 924.600 182.400 925.200 ;
        RECT 196.800 924.600 198.900 925.500 ;
        RECT 166.500 923.700 168.300 924.300 ;
        RECT 176.400 923.700 178.500 924.300 ;
        RECT 166.500 922.500 178.500 923.700 ;
        RECT 181.200 923.400 198.900 924.600 ;
        RECT 202.200 924.300 204.300 925.500 ;
        RECT 208.200 925.200 213.900 926.400 ;
        RECT 217.800 924.300 218.700 927.600 ;
        RECT 202.200 923.400 218.700 924.300 ;
        RECT 176.400 922.200 178.500 922.500 ;
        RECT 181.200 921.300 216.900 922.500 ;
        RECT 181.200 920.700 182.400 921.300 ;
        RECT 215.100 920.700 216.900 921.300 ;
        RECT 168.900 919.800 182.400 920.700 ;
        RECT 193.800 919.800 195.900 920.100 ;
        RECT 168.900 919.050 170.700 919.800 ;
        RECT 160.800 916.950 162.900 919.050 ;
        RECT 166.800 917.250 170.700 919.050 ;
        RECT 188.400 918.300 190.500 919.200 ;
        RECT 166.800 916.950 168.900 917.250 ;
        RECT 179.400 917.100 190.500 918.300 ;
        RECT 192.000 918.000 195.900 919.800 ;
        RECT 200.100 918.300 201.900 920.100 ;
        RECT 201.000 917.100 201.900 918.300 ;
        RECT 161.100 915.300 162.900 916.950 ;
        RECT 179.400 916.500 181.200 917.100 ;
        RECT 188.400 916.200 201.900 917.100 ;
        RECT 204.600 916.800 209.700 918.600 ;
        RECT 211.800 916.950 213.900 919.050 ;
        RECT 204.600 915.300 205.500 916.800 ;
        RECT 161.100 914.100 205.500 915.300 ;
        RECT 211.800 914.100 213.300 916.950 ;
        RECT 176.400 911.400 178.200 913.200 ;
        RECT 184.800 912.000 186.900 913.050 ;
        RECT 206.700 912.600 213.300 914.100 ;
        RECT 158.700 910.200 175.500 911.400 ;
        RECT 119.700 906.600 120.900 908.700 ;
        RECT 77.100 900.600 78.900 903.600 ;
        RECT 95.100 900.000 96.900 903.600 ;
        RECT 98.100 900.600 99.900 903.600 ;
        RECT 101.100 900.000 102.900 903.600 ;
        RECT 119.100 900.600 120.900 906.600 ;
        RECT 122.100 905.700 129.900 907.050 ;
        RECT 146.700 906.600 147.900 908.700 ;
        RECT 122.100 900.600 123.900 905.700 ;
        RECT 125.100 900.000 126.900 904.800 ;
        RECT 128.100 900.600 129.900 905.700 ;
        RECT 146.100 900.600 147.900 906.600 ;
        RECT 149.100 905.700 156.900 907.050 ;
        RECT 149.100 900.600 150.900 905.700 ;
        RECT 152.100 900.000 153.900 904.800 ;
        RECT 155.100 900.600 156.900 905.700 ;
        RECT 158.700 906.600 159.900 910.200 ;
        RECT 173.400 909.300 175.500 910.200 ;
        RECT 162.900 908.700 164.700 909.300 ;
        RECT 162.900 907.500 171.300 908.700 ;
        RECT 169.800 906.600 171.300 907.500 ;
        RECT 176.400 908.400 177.300 911.400 ;
        RECT 181.800 911.100 186.900 912.000 ;
        RECT 181.800 910.200 183.600 911.100 ;
        RECT 184.800 910.950 186.900 911.100 ;
        RECT 191.100 911.100 208.200 912.600 ;
        RECT 191.100 910.500 193.200 911.100 ;
        RECT 191.100 908.700 192.900 910.500 ;
        RECT 209.100 909.900 216.900 911.700 ;
        RECT 176.400 907.200 183.600 908.400 ;
        RECT 178.800 906.600 180.600 907.200 ;
        RECT 182.700 906.600 183.600 907.200 ;
        RECT 198.300 906.600 204.900 908.400 ;
        RECT 209.100 906.600 210.600 909.900 ;
        RECT 217.800 906.600 218.700 923.400 ;
        RECT 158.700 900.600 160.500 906.600 ;
        RECT 164.100 900.000 165.900 906.600 ;
        RECT 169.500 900.600 171.300 906.600 ;
        RECT 173.700 903.600 175.800 905.700 ;
        RECT 176.700 903.600 178.800 905.700 ;
        RECT 179.700 903.600 181.800 905.700 ;
        RECT 182.700 905.400 185.400 906.600 ;
        RECT 183.600 904.500 185.400 905.400 ;
        RECT 187.200 904.500 189.900 906.600 ;
        RECT 173.700 900.600 175.500 903.600 ;
        RECT 176.700 900.600 178.500 903.600 ;
        RECT 179.700 900.600 181.500 903.600 ;
        RECT 182.700 900.000 184.500 903.600 ;
        RECT 187.200 900.600 189.000 904.500 ;
        RECT 193.200 903.600 195.300 905.700 ;
        RECT 196.200 903.600 198.300 905.700 ;
        RECT 199.200 903.600 201.300 905.700 ;
        RECT 202.200 903.600 204.300 905.700 ;
        RECT 206.400 905.400 210.600 906.600 ;
        RECT 190.200 900.000 192.000 903.600 ;
        RECT 193.200 900.600 195.000 903.600 ;
        RECT 196.200 900.600 198.000 903.600 ;
        RECT 199.200 900.600 201.000 903.600 ;
        RECT 202.200 900.600 204.000 903.600 ;
        RECT 206.400 900.600 208.200 905.400 ;
        RECT 211.500 900.000 213.300 906.600 ;
        RECT 216.900 900.600 218.700 906.600 ;
        RECT 220.500 919.050 222.000 929.400 ;
        RECT 242.400 923.400 244.200 936.000 ;
        RECT 247.500 924.900 249.300 935.400 ;
        RECT 250.500 929.400 252.300 936.000 ;
        RECT 269.700 929.400 271.500 936.000 ;
        RECT 250.200 926.100 252.000 927.900 ;
        RECT 270.000 926.100 271.800 927.900 ;
        RECT 272.700 924.900 274.500 935.400 ;
        RECT 247.500 923.400 249.900 924.900 ;
        RECT 220.500 916.950 222.900 919.050 ;
        RECT 220.500 903.600 222.000 916.950 ;
        RECT 242.100 916.050 243.900 917.850 ;
        RECT 248.700 916.050 249.900 923.400 ;
        RECT 272.100 923.400 274.500 924.900 ;
        RECT 277.800 923.400 279.600 936.000 ;
        RECT 296.400 923.400 298.200 936.000 ;
        RECT 301.500 924.900 303.300 935.400 ;
        RECT 304.500 929.400 306.300 936.000 ;
        RECT 323.100 929.400 324.900 935.400 ;
        RECT 326.100 930.000 327.900 936.000 ;
        RECT 324.000 929.100 324.900 929.400 ;
        RECT 329.100 929.400 330.900 935.400 ;
        RECT 332.100 929.400 333.900 936.000 ;
        RECT 350.100 929.400 351.900 936.000 ;
        RECT 353.100 929.400 354.900 935.400 ;
        RECT 371.100 929.400 372.900 935.400 ;
        RECT 374.100 930.000 375.900 936.000 ;
        RECT 329.100 929.100 330.600 929.400 ;
        RECT 324.000 928.200 330.600 929.100 ;
        RECT 304.200 926.100 306.000 927.900 ;
        RECT 301.500 923.400 303.900 924.900 ;
        RECT 250.950 921.450 253.050 922.050 ;
        RECT 259.950 921.450 262.050 922.050 ;
        RECT 250.950 920.550 262.050 921.450 ;
        RECT 250.950 919.950 253.050 920.550 ;
        RECT 259.950 919.950 262.050 920.550 ;
        RECT 272.100 916.050 273.300 923.400 ;
        RECT 278.100 916.050 279.900 917.850 ;
        RECT 296.100 916.050 297.900 917.850 ;
        RECT 302.700 916.050 303.900 923.400 ;
        RECT 324.000 916.050 324.900 928.200 ;
        RECT 329.100 916.050 330.900 917.850 ;
        RECT 350.100 916.050 351.900 917.850 ;
        RECT 353.100 916.050 354.300 929.400 ;
        RECT 372.000 929.100 372.900 929.400 ;
        RECT 377.100 929.400 378.900 935.400 ;
        RECT 380.100 929.400 381.900 936.000 ;
        RECT 377.100 929.100 378.600 929.400 ;
        RECT 372.000 928.200 378.600 929.100 ;
        RECT 372.000 916.050 372.900 928.200 ;
        RECT 398.100 925.500 399.900 935.400 ;
        RECT 401.100 926.400 402.900 936.000 ;
        RECT 404.100 934.500 411.900 935.400 ;
        RECT 404.100 925.500 405.900 934.500 ;
        RECT 398.100 924.600 405.900 925.500 ;
        RECT 407.100 925.800 408.900 933.600 ;
        RECT 410.100 926.700 411.900 934.500 ;
        RECT 413.100 934.500 420.900 935.400 ;
        RECT 413.100 925.800 414.900 934.500 ;
        RECT 407.100 924.900 414.900 925.800 ;
        RECT 416.100 925.800 417.900 933.600 ;
        RECT 373.950 921.450 376.050 922.050 ;
        RECT 388.950 921.450 391.050 922.050 ;
        RECT 373.950 920.550 391.050 921.450 ;
        RECT 373.950 919.950 376.050 920.550 ;
        RECT 388.950 919.950 391.050 920.550 ;
        RECT 377.100 916.050 378.900 917.850 ;
        RECT 401.100 916.050 402.900 917.850 ;
        RECT 410.250 916.050 412.050 917.850 ;
        RECT 416.100 916.050 417.300 925.800 ;
        RECT 419.100 925.200 420.900 934.500 ;
        RECT 437.100 929.400 438.900 936.000 ;
        RECT 440.100 929.400 441.900 935.400 ;
        RECT 458.100 929.400 459.900 935.400 ;
        RECT 461.100 930.000 462.900 936.000 ;
        RECT 437.100 916.050 438.900 917.850 ;
        RECT 440.100 916.050 441.300 929.400 ;
        RECT 459.000 929.100 459.900 929.400 ;
        RECT 464.100 929.400 465.900 935.400 ;
        RECT 467.100 929.400 468.900 936.000 ;
        RECT 485.100 929.400 486.900 936.000 ;
        RECT 488.100 929.400 489.900 935.400 ;
        RECT 491.100 929.400 492.900 936.000 ;
        RECT 464.100 929.100 465.600 929.400 ;
        RECT 459.000 928.200 465.600 929.100 ;
        RECT 459.000 916.050 459.900 928.200 ;
        RECT 460.950 921.450 463.050 922.050 ;
        RECT 484.950 921.450 487.050 922.050 ;
        RECT 460.950 920.550 487.050 921.450 ;
        RECT 460.950 919.950 463.050 920.550 ;
        RECT 484.950 919.950 487.050 920.550 ;
        RECT 464.100 916.050 465.900 917.850 ;
        RECT 488.700 916.050 489.900 929.400 ;
        RECT 510.000 924.600 511.800 935.400 ;
        RECT 510.000 923.400 513.600 924.600 ;
        RECT 515.100 923.400 516.900 936.000 ;
        RECT 533.700 929.400 535.500 936.000 ;
        RECT 534.000 926.100 535.800 927.900 ;
        RECT 536.700 924.900 538.500 935.400 ;
        RECT 536.100 923.400 538.500 924.900 ;
        RECT 541.800 923.400 543.600 936.000 ;
        RECT 561.000 924.600 562.800 935.400 ;
        RECT 561.000 923.400 564.600 924.600 ;
        RECT 566.100 923.400 567.900 936.000 ;
        RECT 584.100 929.400 585.900 936.000 ;
        RECT 587.100 929.400 588.900 935.400 ;
        RECT 590.100 929.400 591.900 936.000 ;
        RECT 509.100 916.050 510.900 917.850 ;
        RECT 512.700 916.050 513.600 923.400 ;
        RECT 514.950 916.050 516.750 917.850 ;
        RECT 536.100 916.050 537.300 923.400 ;
        RECT 542.100 916.050 543.900 917.850 ;
        RECT 560.100 916.050 561.900 917.850 ;
        RECT 563.700 916.050 564.600 923.400 ;
        RECT 565.950 916.050 567.750 917.850 ;
        RECT 587.700 916.050 588.900 929.400 ;
        RECT 609.000 924.600 610.800 935.400 ;
        RECT 609.000 923.400 612.600 924.600 ;
        RECT 614.100 923.400 615.900 936.000 ;
        RECT 632.100 923.400 633.900 936.000 ;
        RECT 637.200 924.600 639.000 935.400 ;
        RECT 635.400 923.400 639.000 924.600 ;
        RECT 656.100 923.400 657.900 935.400 ;
        RECT 659.100 924.300 660.900 935.400 ;
        RECT 662.100 925.200 663.900 936.000 ;
        RECT 665.100 924.300 666.900 935.400 ;
        RECT 659.100 923.400 666.900 924.300 ;
        RECT 683.100 934.500 690.900 935.400 ;
        RECT 683.100 923.400 684.900 934.500 ;
        RECT 608.100 916.050 609.900 917.850 ;
        RECT 611.700 916.050 612.600 923.400 ;
        RECT 613.950 916.050 615.750 917.850 ;
        RECT 632.250 916.050 634.050 917.850 ;
        RECT 635.400 916.050 636.300 923.400 ;
        RECT 638.100 916.050 639.900 917.850 ;
        RECT 656.400 916.050 657.300 923.400 ;
        RECT 686.100 922.500 687.900 933.600 ;
        RECT 689.100 924.600 690.900 934.500 ;
        RECT 692.100 925.500 693.900 936.000 ;
        RECT 695.100 924.600 696.900 935.400 ;
        RECT 689.100 923.700 696.900 924.600 ;
        RECT 713.100 923.400 714.900 936.000 ;
        RECT 718.200 924.600 720.000 935.400 ;
        RECT 737.100 929.400 738.900 936.000 ;
        RECT 740.100 929.400 741.900 935.400 ;
        RECT 716.400 923.400 720.000 924.600 ;
        RECT 664.950 921.450 667.050 922.050 ;
        RECT 676.950 921.450 679.050 922.050 ;
        RECT 686.100 921.600 690.900 922.500 ;
        RECT 664.950 920.550 679.050 921.450 ;
        RECT 664.950 919.950 667.050 920.550 ;
        RECT 676.950 919.950 679.050 920.550 ;
        RECT 661.950 916.050 663.750 917.850 ;
        RECT 686.100 916.050 687.900 917.850 ;
        RECT 690.000 916.050 690.900 921.600 ;
        RECT 691.950 916.050 693.750 917.850 ;
        RECT 713.250 916.050 715.050 917.850 ;
        RECT 716.400 916.050 717.300 923.400 ;
        RECT 719.100 916.050 720.900 917.850 ;
        RECT 737.100 916.050 738.900 917.850 ;
        RECT 740.100 916.050 741.300 929.400 ;
        RECT 758.400 923.400 760.200 936.000 ;
        RECT 763.500 924.900 765.300 935.400 ;
        RECT 766.500 929.400 768.300 936.000 ;
        RECT 785.100 929.400 786.900 936.000 ;
        RECT 788.100 929.400 789.900 935.400 ;
        RECT 791.100 929.400 792.900 936.000 ;
        RECT 809.100 929.400 810.900 936.000 ;
        RECT 812.100 929.400 813.900 935.400 ;
        RECT 766.200 926.100 768.000 927.900 ;
        RECT 763.500 923.400 765.900 924.900 ;
        RECT 758.100 916.050 759.900 917.850 ;
        RECT 764.700 916.050 765.900 923.400 ;
        RECT 788.100 916.050 789.300 929.400 ;
        RECT 241.950 913.950 244.050 916.050 ;
        RECT 244.950 913.950 247.050 916.050 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 301.950 913.950 304.050 916.050 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 322.950 913.950 325.050 916.050 ;
        RECT 325.950 913.950 328.050 916.050 ;
        RECT 328.950 913.950 331.050 916.050 ;
        RECT 331.950 913.950 334.050 916.050 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 373.950 913.950 376.050 916.050 ;
        RECT 376.950 913.950 379.050 916.050 ;
        RECT 379.950 913.950 382.050 916.050 ;
        RECT 400.800 913.950 402.900 916.050 ;
        RECT 406.950 913.950 409.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 415.500 913.950 417.600 916.050 ;
        RECT 436.950 913.950 439.050 916.050 ;
        RECT 439.950 913.950 442.050 916.050 ;
        RECT 457.950 913.950 460.050 916.050 ;
        RECT 460.950 913.950 463.050 916.050 ;
        RECT 463.950 913.950 466.050 916.050 ;
        RECT 466.950 913.950 469.050 916.050 ;
        RECT 484.950 913.950 487.050 916.050 ;
        RECT 487.950 913.950 490.050 916.050 ;
        RECT 490.950 913.950 493.050 916.050 ;
        RECT 508.950 913.950 511.050 916.050 ;
        RECT 511.950 913.950 514.050 916.050 ;
        RECT 514.950 913.950 517.050 916.050 ;
        RECT 532.950 913.950 535.050 916.050 ;
        RECT 535.950 913.950 538.050 916.050 ;
        RECT 538.950 913.950 541.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 559.950 913.950 562.050 916.050 ;
        RECT 562.950 913.950 565.050 916.050 ;
        RECT 565.950 913.950 568.050 916.050 ;
        RECT 583.950 913.950 586.050 916.050 ;
        RECT 586.950 913.950 589.050 916.050 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 607.950 913.950 610.050 916.050 ;
        RECT 610.950 913.950 613.050 916.050 ;
        RECT 613.950 913.950 616.050 916.050 ;
        RECT 631.950 913.950 634.050 916.050 ;
        RECT 634.950 913.950 637.050 916.050 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 655.950 913.950 658.050 916.050 ;
        RECT 658.950 913.950 661.050 916.050 ;
        RECT 661.950 913.950 664.050 916.050 ;
        RECT 664.950 913.950 667.050 916.050 ;
        RECT 682.950 913.950 685.050 916.050 ;
        RECT 685.950 913.950 688.050 916.050 ;
        RECT 688.950 913.950 691.050 916.050 ;
        RECT 691.950 913.950 694.050 916.050 ;
        RECT 694.950 913.950 697.050 916.050 ;
        RECT 712.950 913.950 715.050 916.050 ;
        RECT 715.950 913.950 718.050 916.050 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 736.950 913.950 739.050 916.050 ;
        RECT 739.950 913.950 742.050 916.050 ;
        RECT 757.950 913.950 760.050 916.050 ;
        RECT 760.950 913.950 763.050 916.050 ;
        RECT 763.950 913.950 766.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 809.100 913.950 811.200 916.050 ;
        RECT 245.100 912.150 246.900 913.950 ;
        RECT 248.700 909.600 249.900 913.950 ;
        RECT 251.100 912.150 252.900 913.950 ;
        RECT 269.100 912.150 270.900 913.950 ;
        RECT 272.100 909.600 273.300 913.950 ;
        RECT 275.100 912.150 276.900 913.950 ;
        RECT 299.100 912.150 300.900 913.950 ;
        RECT 248.700 908.700 252.300 909.600 ;
        RECT 242.100 905.700 249.900 907.050 ;
        RECT 220.500 900.600 222.300 903.600 ;
        RECT 223.500 900.000 225.300 903.600 ;
        RECT 242.100 900.600 243.900 905.700 ;
        RECT 245.100 900.000 246.900 904.800 ;
        RECT 248.100 900.600 249.900 905.700 ;
        RECT 251.100 906.600 252.300 908.700 ;
        RECT 269.700 908.700 273.300 909.600 ;
        RECT 302.700 909.600 303.900 913.950 ;
        RECT 305.100 912.150 306.900 913.950 ;
        RECT 324.000 910.200 324.900 913.950 ;
        RECT 326.100 912.150 327.900 913.950 ;
        RECT 332.100 912.150 333.900 913.950 ;
        RECT 302.700 908.700 306.300 909.600 ;
        RECT 324.000 909.000 327.300 910.200 ;
        RECT 269.700 906.600 270.900 908.700 ;
        RECT 251.100 900.600 252.900 906.600 ;
        RECT 269.100 900.600 270.900 906.600 ;
        RECT 272.100 905.700 279.900 907.050 ;
        RECT 272.100 900.600 273.900 905.700 ;
        RECT 275.100 900.000 276.900 904.800 ;
        RECT 278.100 900.600 279.900 905.700 ;
        RECT 296.100 905.700 303.900 907.050 ;
        RECT 296.100 900.600 297.900 905.700 ;
        RECT 299.100 900.000 300.900 904.800 ;
        RECT 302.100 900.600 303.900 905.700 ;
        RECT 305.100 906.600 306.300 908.700 ;
        RECT 305.100 900.600 306.900 906.600 ;
        RECT 325.500 900.600 327.300 909.000 ;
        RECT 332.100 900.000 333.900 909.600 ;
        RECT 353.100 903.600 354.300 913.950 ;
        RECT 372.000 910.200 372.900 913.950 ;
        RECT 374.100 912.150 375.900 913.950 ;
        RECT 380.100 912.150 381.900 913.950 ;
        RECT 406.950 912.150 408.750 913.950 ;
        RECT 372.000 909.000 375.300 910.200 ;
        RECT 350.100 900.000 351.900 903.600 ;
        RECT 353.100 900.600 354.900 903.600 ;
        RECT 373.500 900.600 375.300 909.000 ;
        RECT 380.100 900.000 381.900 909.600 ;
        RECT 397.950 909.450 400.050 910.050 ;
        RECT 409.950 909.450 412.050 910.050 ;
        RECT 397.950 908.550 412.050 909.450 ;
        RECT 397.950 907.950 400.050 908.550 ;
        RECT 409.950 907.950 412.050 908.550 ;
        RECT 416.100 905.400 417.300 913.950 ;
        RECT 404.700 904.500 417.300 905.400 ;
        RECT 404.700 903.600 405.600 904.500 ;
        RECT 411.900 903.600 412.800 904.500 ;
        RECT 440.100 903.600 441.300 913.950 ;
        RECT 459.000 910.200 459.900 913.950 ;
        RECT 461.100 912.150 462.900 913.950 ;
        RECT 467.100 912.150 468.900 913.950 ;
        RECT 485.100 912.150 486.900 913.950 ;
        RECT 459.000 909.000 462.300 910.200 ;
        RECT 400.800 900.000 402.900 903.600 ;
        RECT 404.100 900.600 405.900 903.600 ;
        RECT 407.100 900.000 408.900 903.600 ;
        RECT 410.100 900.600 412.800 903.600 ;
        RECT 437.100 900.000 438.900 903.600 ;
        RECT 440.100 900.600 441.900 903.600 ;
        RECT 460.500 900.600 462.300 909.000 ;
        RECT 467.100 900.000 468.900 909.600 ;
        RECT 488.700 908.700 489.900 913.950 ;
        RECT 490.950 912.150 492.750 913.950 ;
        RECT 485.700 907.800 489.900 908.700 ;
        RECT 485.700 900.600 487.500 907.800 ;
        RECT 490.800 900.000 492.600 906.600 ;
        RECT 512.700 903.600 513.600 913.950 ;
        RECT 533.100 912.150 534.900 913.950 ;
        RECT 536.100 909.600 537.300 913.950 ;
        RECT 539.100 912.150 540.900 913.950 ;
        RECT 533.700 908.700 537.300 909.600 ;
        RECT 533.700 906.600 534.900 908.700 ;
        RECT 509.100 900.000 510.900 903.600 ;
        RECT 512.100 900.600 513.900 903.600 ;
        RECT 515.100 900.000 516.900 903.600 ;
        RECT 533.100 900.600 534.900 906.600 ;
        RECT 536.100 905.700 543.900 907.050 ;
        RECT 536.100 900.600 537.900 905.700 ;
        RECT 539.100 900.000 540.900 904.800 ;
        RECT 542.100 900.600 543.900 905.700 ;
        RECT 563.700 903.600 564.600 913.950 ;
        RECT 584.100 912.150 585.900 913.950 ;
        RECT 587.700 908.700 588.900 913.950 ;
        RECT 589.950 912.150 591.750 913.950 ;
        RECT 584.700 907.800 588.900 908.700 ;
        RECT 589.950 909.450 592.050 910.050 ;
        RECT 595.950 909.450 598.050 910.050 ;
        RECT 589.950 908.550 598.050 909.450 ;
        RECT 589.950 907.950 592.050 908.550 ;
        RECT 595.950 907.950 598.050 908.550 ;
        RECT 560.100 900.000 561.900 903.600 ;
        RECT 563.100 900.600 564.900 903.600 ;
        RECT 566.100 900.000 567.900 903.600 ;
        RECT 584.700 900.600 586.500 907.800 ;
        RECT 589.800 900.000 591.600 906.600 ;
        RECT 611.700 903.600 612.600 913.950 ;
        RECT 635.400 903.600 636.300 913.950 ;
        RECT 656.400 906.600 657.300 913.950 ;
        RECT 658.950 912.150 660.750 913.950 ;
        RECT 665.100 912.150 666.900 913.950 ;
        RECT 683.100 912.150 684.900 913.950 ;
        RECT 689.700 906.600 690.900 913.950 ;
        RECT 694.950 912.150 696.750 913.950 ;
        RECT 656.400 905.400 661.500 906.600 ;
        RECT 608.100 900.000 609.900 903.600 ;
        RECT 611.100 900.600 612.900 903.600 ;
        RECT 614.100 900.000 615.900 903.600 ;
        RECT 632.100 900.000 633.900 903.600 ;
        RECT 635.100 900.600 636.900 903.600 ;
        RECT 638.100 900.000 639.900 903.600 ;
        RECT 656.700 900.000 658.500 903.600 ;
        RECT 659.700 900.600 661.500 905.400 ;
        RECT 664.200 900.000 666.000 906.600 ;
        RECT 685.500 900.000 687.300 906.600 ;
        RECT 690.000 900.600 691.800 906.600 ;
        RECT 694.500 900.000 696.300 906.600 ;
        RECT 716.400 903.600 717.300 913.950 ;
        RECT 721.950 906.450 724.050 907.050 ;
        RECT 730.950 906.450 733.050 907.050 ;
        RECT 721.950 905.550 733.050 906.450 ;
        RECT 721.950 904.950 724.050 905.550 ;
        RECT 730.950 904.950 733.050 905.550 ;
        RECT 740.100 903.600 741.300 913.950 ;
        RECT 761.100 912.150 762.900 913.950 ;
        RECT 764.700 909.600 765.900 913.950 ;
        RECT 767.100 912.150 768.900 913.950 ;
        RECT 785.250 912.150 787.050 913.950 ;
        RECT 764.700 908.700 768.300 909.600 ;
        RECT 758.100 905.700 765.900 907.050 ;
        RECT 713.100 900.000 714.900 903.600 ;
        RECT 716.100 900.600 717.900 903.600 ;
        RECT 719.100 900.000 720.900 903.600 ;
        RECT 737.100 900.000 738.900 903.600 ;
        RECT 740.100 900.600 741.900 903.600 ;
        RECT 758.100 900.600 759.900 905.700 ;
        RECT 761.100 900.000 762.900 904.800 ;
        RECT 764.100 900.600 765.900 905.700 ;
        RECT 767.100 906.600 768.300 908.700 ;
        RECT 788.100 908.700 789.300 913.950 ;
        RECT 791.100 912.150 792.900 913.950 ;
        RECT 809.250 912.150 811.050 913.950 ;
        RECT 812.100 909.300 813.000 929.400 ;
        RECT 815.100 924.000 816.900 936.000 ;
        RECT 818.100 923.400 819.900 935.400 ;
        RECT 836.100 929.400 837.900 936.000 ;
        RECT 839.100 929.400 840.900 935.400 ;
        RECT 842.100 930.000 843.900 936.000 ;
        RECT 839.400 929.100 840.900 929.400 ;
        RECT 845.100 929.400 846.900 935.400 ;
        RECT 863.100 929.400 864.900 936.000 ;
        RECT 866.100 929.400 867.900 935.400 ;
        RECT 869.100 930.000 870.900 936.000 ;
        RECT 845.100 929.100 846.000 929.400 ;
        RECT 839.400 928.200 846.000 929.100 ;
        RECT 866.400 929.100 867.900 929.400 ;
        RECT 872.100 929.400 873.900 935.400 ;
        RECT 872.100 929.100 873.000 929.400 ;
        RECT 866.400 928.200 873.000 929.100 ;
        RECT 823.950 924.450 826.050 925.050 ;
        RECT 841.950 924.450 844.050 925.050 ;
        RECT 823.950 923.550 844.050 924.450 ;
        RECT 814.200 916.050 816.000 917.850 ;
        RECT 818.400 916.050 819.300 923.400 ;
        RECT 823.950 922.950 826.050 923.550 ;
        RECT 841.950 922.950 844.050 923.550 ;
        RECT 839.100 916.050 840.900 917.850 ;
        RECT 845.100 916.050 846.000 928.200 ;
        RECT 853.950 918.450 856.050 919.050 ;
        RECT 859.950 918.450 862.050 919.050 ;
        RECT 853.950 917.550 862.050 918.450 ;
        RECT 853.950 916.950 856.050 917.550 ;
        RECT 859.950 916.950 862.050 917.550 ;
        RECT 866.100 916.050 867.900 917.850 ;
        RECT 872.100 916.050 873.000 928.200 ;
        RECT 890.100 924.300 891.900 935.400 ;
        RECT 893.100 925.200 894.900 936.000 ;
        RECT 896.100 924.300 897.900 935.400 ;
        RECT 890.100 923.400 897.900 924.300 ;
        RECT 899.100 923.400 900.900 935.400 ;
        RECT 917.100 929.400 918.900 936.000 ;
        RECT 920.100 929.400 921.900 935.400 ;
        RECT 923.100 930.000 924.900 936.000 ;
        RECT 920.400 929.100 921.900 929.400 ;
        RECT 926.100 929.400 927.900 935.400 ;
        RECT 941.100 929.400 942.900 936.000 ;
        RECT 944.100 929.400 945.900 935.400 ;
        RECT 947.100 929.400 948.900 936.000 ;
        RECT 926.100 929.100 927.000 929.400 ;
        RECT 920.400 928.200 927.000 929.100 ;
        RECT 893.250 916.050 895.050 917.850 ;
        RECT 899.700 916.050 900.600 923.400 ;
        RECT 907.950 921.450 910.050 922.050 ;
        RECT 916.950 921.450 919.050 922.050 ;
        RECT 907.950 920.550 919.050 921.450 ;
        RECT 907.950 919.950 910.050 920.550 ;
        RECT 916.950 919.950 919.050 920.550 ;
        RECT 920.100 916.050 921.900 917.850 ;
        RECT 926.100 916.050 927.000 928.200 ;
        RECT 944.700 916.050 945.900 929.400 ;
        RECT 965.100 923.400 966.900 935.400 ;
        RECT 968.100 924.300 969.900 935.400 ;
        RECT 971.100 925.200 972.900 936.000 ;
        RECT 974.100 924.300 975.900 935.400 ;
        RECT 992.100 929.400 993.900 936.000 ;
        RECT 995.100 929.400 996.900 935.400 ;
        RECT 998.100 930.000 999.900 936.000 ;
        RECT 995.400 929.100 996.900 929.400 ;
        RECT 1001.100 929.400 1002.900 935.400 ;
        RECT 1001.100 929.100 1002.000 929.400 ;
        RECT 995.400 928.200 1002.000 929.100 ;
        RECT 968.100 923.400 975.900 924.300 ;
        RECT 965.400 916.050 966.300 923.400 ;
        RECT 970.950 916.050 972.750 917.850 ;
        RECT 995.100 916.050 996.900 917.850 ;
        RECT 1001.100 916.050 1002.000 928.200 ;
        RECT 1019.100 923.400 1020.900 936.000 ;
        RECT 1024.200 924.600 1026.000 935.400 ;
        RECT 1022.400 923.400 1026.000 924.600 ;
        RECT 1019.250 916.050 1021.050 917.850 ;
        RECT 1022.400 916.050 1023.300 923.400 ;
        RECT 1025.100 916.050 1026.900 917.850 ;
        RECT 814.500 913.950 816.600 916.050 ;
        RECT 817.800 913.950 819.900 916.050 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 838.950 913.950 841.050 916.050 ;
        RECT 841.950 913.950 844.050 916.050 ;
        RECT 844.950 913.950 847.050 916.050 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 865.950 913.950 868.050 916.050 ;
        RECT 868.950 913.950 871.050 916.050 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 892.950 913.950 895.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 916.950 913.950 919.050 916.050 ;
        RECT 919.950 913.950 922.050 916.050 ;
        RECT 922.950 913.950 925.050 916.050 ;
        RECT 925.950 913.950 928.050 916.050 ;
        RECT 940.950 913.950 943.050 916.050 ;
        RECT 943.950 913.950 946.050 916.050 ;
        RECT 946.950 913.950 949.050 916.050 ;
        RECT 964.950 913.950 967.050 916.050 ;
        RECT 967.950 913.950 970.050 916.050 ;
        RECT 970.950 913.950 973.050 916.050 ;
        RECT 973.950 913.950 976.050 916.050 ;
        RECT 991.950 913.950 994.050 916.050 ;
        RECT 994.950 913.950 997.050 916.050 ;
        RECT 997.950 913.950 1000.050 916.050 ;
        RECT 1000.950 913.950 1003.050 916.050 ;
        RECT 1018.950 913.950 1021.050 916.050 ;
        RECT 1021.950 913.950 1024.050 916.050 ;
        RECT 1024.950 913.950 1027.050 916.050 ;
        RECT 788.100 907.800 792.300 908.700 ;
        RECT 767.100 900.600 768.900 906.600 ;
        RECT 785.400 900.000 787.200 906.600 ;
        RECT 790.500 900.600 792.300 907.800 ;
        RECT 809.100 908.400 817.500 909.300 ;
        RECT 809.100 900.600 810.900 908.400 ;
        RECT 815.700 907.500 817.500 908.400 ;
        RECT 818.400 906.600 819.300 913.950 ;
        RECT 836.100 912.150 837.900 913.950 ;
        RECT 842.100 912.150 843.900 913.950 ;
        RECT 845.100 910.200 846.000 913.950 ;
        RECT 863.100 912.150 864.900 913.950 ;
        RECT 869.100 912.150 870.900 913.950 ;
        RECT 872.100 910.200 873.000 913.950 ;
        RECT 890.100 912.150 891.900 913.950 ;
        RECT 896.250 912.150 898.050 913.950 ;
        RECT 813.600 900.000 815.400 906.600 ;
        RECT 816.600 904.800 819.300 906.600 ;
        RECT 816.600 900.600 818.400 904.800 ;
        RECT 836.100 900.000 837.900 909.600 ;
        RECT 842.700 909.000 846.000 910.200 ;
        RECT 842.700 900.600 844.500 909.000 ;
        RECT 863.100 900.000 864.900 909.600 ;
        RECT 869.700 909.000 873.000 910.200 ;
        RECT 869.700 900.600 871.500 909.000 ;
        RECT 899.700 906.600 900.600 913.950 ;
        RECT 917.100 912.150 918.900 913.950 ;
        RECT 923.100 912.150 924.900 913.950 ;
        RECT 926.100 910.200 927.000 913.950 ;
        RECT 941.100 912.150 942.900 913.950 ;
        RECT 891.000 900.000 892.800 906.600 ;
        RECT 895.500 905.400 900.600 906.600 ;
        RECT 895.500 900.600 897.300 905.400 ;
        RECT 898.500 900.000 900.300 903.600 ;
        RECT 917.100 900.000 918.900 909.600 ;
        RECT 923.700 909.000 927.000 910.200 ;
        RECT 923.700 900.600 925.500 909.000 ;
        RECT 944.700 908.700 945.900 913.950 ;
        RECT 946.950 912.150 948.750 913.950 ;
        RECT 941.700 907.800 945.900 908.700 ;
        RECT 946.950 909.450 949.050 910.050 ;
        RECT 958.950 909.450 961.050 910.050 ;
        RECT 946.950 908.550 961.050 909.450 ;
        RECT 946.950 907.950 949.050 908.550 ;
        RECT 958.950 907.950 961.050 908.550 ;
        RECT 941.700 900.600 943.500 907.800 ;
        RECT 965.400 906.600 966.300 913.950 ;
        RECT 967.950 912.150 969.750 913.950 ;
        RECT 974.100 912.150 975.900 913.950 ;
        RECT 992.100 912.150 993.900 913.950 ;
        RECT 998.100 912.150 999.900 913.950 ;
        RECT 1001.100 910.200 1002.000 913.950 ;
        RECT 946.800 900.000 948.600 906.600 ;
        RECT 965.400 905.400 970.500 906.600 ;
        RECT 965.700 900.000 967.500 903.600 ;
        RECT 968.700 900.600 970.500 905.400 ;
        RECT 973.200 900.000 975.000 906.600 ;
        RECT 992.100 900.000 993.900 909.600 ;
        RECT 998.700 909.000 1002.000 910.200 ;
        RECT 998.700 900.600 1000.500 909.000 ;
        RECT 1022.400 903.600 1023.300 913.950 ;
        RECT 1019.100 900.000 1020.900 903.600 ;
        RECT 1022.100 900.600 1023.900 903.600 ;
        RECT 1025.100 900.000 1026.900 903.600 ;
        RECT 17.100 890.400 18.900 896.400 ;
        RECT 20.100 890.400 21.900 897.000 ;
        RECT 23.100 893.400 24.900 896.400 ;
        RECT 17.100 883.050 18.300 890.400 ;
        RECT 23.700 889.500 24.900 893.400 ;
        RECT 19.200 888.600 24.900 889.500 ;
        RECT 26.700 890.400 28.500 896.400 ;
        RECT 32.100 890.400 33.900 897.000 ;
        RECT 37.500 890.400 39.300 896.400 ;
        RECT 41.700 893.400 43.500 896.400 ;
        RECT 44.700 893.400 46.500 896.400 ;
        RECT 47.700 893.400 49.500 896.400 ;
        RECT 50.700 893.400 52.500 897.000 ;
        RECT 41.700 891.300 43.800 893.400 ;
        RECT 44.700 891.300 46.800 893.400 ;
        RECT 47.700 891.300 49.800 893.400 ;
        RECT 55.200 892.500 57.000 896.400 ;
        RECT 58.200 893.400 60.000 897.000 ;
        RECT 61.200 893.400 63.000 896.400 ;
        RECT 64.200 893.400 66.000 896.400 ;
        RECT 67.200 893.400 69.000 896.400 ;
        RECT 70.200 893.400 72.000 896.400 ;
        RECT 51.600 891.600 53.400 892.500 ;
        RECT 50.700 890.400 53.400 891.600 ;
        RECT 55.200 890.400 57.900 892.500 ;
        RECT 61.200 891.300 63.300 893.400 ;
        RECT 64.200 891.300 66.300 893.400 ;
        RECT 67.200 891.300 69.300 893.400 ;
        RECT 70.200 891.300 72.300 893.400 ;
        RECT 74.400 891.600 76.200 896.400 ;
        RECT 74.400 890.400 78.600 891.600 ;
        RECT 79.500 890.400 81.300 897.000 ;
        RECT 84.900 890.400 86.700 896.400 ;
        RECT 19.200 887.700 21.000 888.600 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 17.100 873.600 18.300 880.950 ;
        RECT 20.100 876.300 21.000 887.700 ;
        RECT 26.700 886.800 27.900 890.400 ;
        RECT 37.800 889.500 39.300 890.400 ;
        RECT 46.800 889.800 48.600 890.400 ;
        RECT 50.700 889.800 51.600 890.400 ;
        RECT 30.900 888.300 39.300 889.500 ;
        RECT 44.400 888.600 51.600 889.800 ;
        RECT 66.300 888.600 72.900 890.400 ;
        RECT 30.900 887.700 32.700 888.300 ;
        RECT 41.400 886.800 43.500 887.700 ;
        RECT 26.700 885.600 43.500 886.800 ;
        RECT 44.400 885.600 45.300 888.600 ;
        RECT 49.800 885.900 51.600 886.800 ;
        RECT 59.100 886.500 60.900 888.300 ;
        RECT 77.100 887.100 78.600 890.400 ;
        RECT 52.800 885.900 54.900 886.050 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 22.800 879.150 24.600 880.950 ;
        RECT 19.200 875.400 21.000 876.300 ;
        RECT 19.200 874.500 24.900 875.400 ;
        RECT 17.100 861.600 18.900 873.600 ;
        RECT 20.100 861.000 21.900 871.800 ;
        RECT 23.700 867.600 24.900 874.500 ;
        RECT 26.700 869.400 27.900 885.600 ;
        RECT 44.400 883.800 46.200 885.600 ;
        RECT 49.800 885.000 54.900 885.900 ;
        RECT 52.800 883.950 54.900 885.000 ;
        RECT 59.100 885.900 61.200 886.500 ;
        RECT 59.100 884.400 76.200 885.900 ;
        RECT 77.100 885.300 84.900 887.100 ;
        RECT 74.700 882.900 81.300 884.400 ;
        RECT 29.100 881.700 73.500 882.900 ;
        RECT 29.100 880.050 30.900 881.700 ;
        RECT 28.800 877.950 30.900 880.050 ;
        RECT 34.800 879.750 36.900 880.050 ;
        RECT 47.400 879.900 49.200 880.500 ;
        RECT 56.400 879.900 69.900 880.800 ;
        RECT 34.800 877.950 38.700 879.750 ;
        RECT 47.400 878.700 58.500 879.900 ;
        RECT 36.900 877.200 38.700 877.950 ;
        RECT 56.400 877.800 58.500 878.700 ;
        RECT 60.000 877.200 63.900 879.000 ;
        RECT 69.000 878.700 69.900 879.900 ;
        RECT 36.900 876.300 50.400 877.200 ;
        RECT 61.800 876.900 63.900 877.200 ;
        RECT 68.100 876.900 69.900 878.700 ;
        RECT 72.600 880.200 73.500 881.700 ;
        RECT 72.600 878.400 77.700 880.200 ;
        RECT 79.800 880.050 81.300 882.900 ;
        RECT 79.800 877.950 81.900 880.050 ;
        RECT 49.200 875.700 50.400 876.300 ;
        RECT 83.100 875.700 84.900 876.300 ;
        RECT 44.400 874.500 46.500 874.800 ;
        RECT 49.200 874.500 84.900 875.700 ;
        RECT 34.500 873.300 46.500 874.500 ;
        RECT 85.800 873.600 86.700 890.400 ;
        RECT 34.500 872.700 36.300 873.300 ;
        RECT 44.400 872.700 46.500 873.300 ;
        RECT 49.200 872.400 66.900 873.600 ;
        RECT 31.200 871.800 33.000 872.100 ;
        RECT 49.200 871.800 50.400 872.400 ;
        RECT 31.200 870.600 50.400 871.800 ;
        RECT 64.800 871.500 66.900 872.400 ;
        RECT 70.200 872.700 86.700 873.600 ;
        RECT 70.200 871.500 72.300 872.700 ;
        RECT 31.200 870.300 33.000 870.600 ;
        RECT 26.700 868.500 30.300 869.400 ;
        RECT 29.400 867.600 30.300 868.500 ;
        RECT 23.100 861.600 24.900 867.600 ;
        RECT 26.700 861.000 28.500 867.600 ;
        RECT 29.400 866.700 31.500 867.600 ;
        RECT 29.700 861.600 31.500 866.700 ;
        RECT 32.700 861.000 34.500 867.600 ;
        RECT 35.700 861.600 37.500 870.600 ;
        RECT 47.700 867.600 49.800 869.700 ;
        RECT 55.200 869.100 58.500 871.200 ;
        RECT 38.700 861.000 40.500 867.600 ;
        RECT 42.300 864.600 44.400 866.700 ;
        RECT 45.300 864.600 47.400 866.700 ;
        RECT 42.300 861.600 44.100 864.600 ;
        RECT 45.300 861.600 47.100 864.600 ;
        RECT 48.300 861.600 50.100 867.600 ;
        RECT 51.300 861.000 53.100 867.600 ;
        RECT 55.200 861.600 57.000 869.100 ;
        RECT 61.200 867.600 63.900 871.500 ;
        RECT 76.200 870.600 81.900 871.800 ;
        RECT 73.500 869.700 75.300 870.300 ;
        RECT 67.200 868.500 75.300 869.700 ;
        RECT 67.200 867.600 69.300 868.500 ;
        RECT 76.200 867.600 77.400 870.600 ;
        RECT 80.100 870.000 81.900 870.600 ;
        RECT 85.800 869.400 86.700 872.700 ;
        RECT 82.800 868.500 86.700 869.400 ;
        RECT 88.500 893.400 90.300 896.400 ;
        RECT 91.500 893.400 93.300 897.000 ;
        RECT 88.500 880.050 90.000 893.400 ;
        RECT 110.100 890.400 111.900 896.400 ;
        RECT 113.100 891.000 114.900 897.000 ;
        RECT 119.700 896.400 120.900 897.000 ;
        RECT 116.100 893.400 117.900 896.400 ;
        RECT 119.100 893.400 120.900 896.400 ;
        RECT 110.100 883.050 111.000 890.400 ;
        RECT 116.700 889.200 117.600 893.400 ;
        RECT 112.200 888.300 117.600 889.200 ;
        RECT 137.700 889.200 139.500 896.400 ;
        RECT 142.800 890.400 144.600 897.000 ;
        RECT 161.100 890.400 162.900 897.000 ;
        RECT 164.100 890.400 165.900 896.400 ;
        RECT 167.700 890.400 169.500 896.400 ;
        RECT 173.100 890.400 174.900 897.000 ;
        RECT 178.500 890.400 180.300 896.400 ;
        RECT 182.700 893.400 184.500 896.400 ;
        RECT 185.700 893.400 187.500 896.400 ;
        RECT 188.700 893.400 190.500 896.400 ;
        RECT 191.700 893.400 193.500 897.000 ;
        RECT 182.700 891.300 184.800 893.400 ;
        RECT 185.700 891.300 187.800 893.400 ;
        RECT 188.700 891.300 190.800 893.400 ;
        RECT 196.200 892.500 198.000 896.400 ;
        RECT 199.200 893.400 201.000 897.000 ;
        RECT 202.200 893.400 204.000 896.400 ;
        RECT 205.200 893.400 207.000 896.400 ;
        RECT 208.200 893.400 210.000 896.400 ;
        RECT 211.200 893.400 213.000 896.400 ;
        RECT 192.600 891.600 194.400 892.500 ;
        RECT 191.700 890.400 194.400 891.600 ;
        RECT 196.200 890.400 198.900 892.500 ;
        RECT 202.200 891.300 204.300 893.400 ;
        RECT 205.200 891.300 207.300 893.400 ;
        RECT 208.200 891.300 210.300 893.400 ;
        RECT 211.200 891.300 213.300 893.400 ;
        RECT 215.400 891.600 217.200 896.400 ;
        RECT 215.400 890.400 219.600 891.600 ;
        RECT 220.500 890.400 222.300 897.000 ;
        RECT 225.900 890.400 227.700 896.400 ;
        RECT 137.700 888.300 141.900 889.200 ;
        RECT 112.200 887.400 114.300 888.300 ;
        RECT 110.100 880.950 112.200 883.050 ;
        RECT 88.500 877.950 90.900 880.050 ;
        RECT 82.800 867.600 84.000 868.500 ;
        RECT 88.500 867.600 90.000 877.950 ;
        RECT 111.000 873.600 112.200 880.950 ;
        RECT 113.400 876.900 114.300 887.400 ;
        RECT 118.800 883.050 120.600 884.850 ;
        RECT 137.100 883.050 138.900 884.850 ;
        RECT 140.700 883.050 141.900 888.300 ;
        RECT 142.950 883.050 144.750 884.850 ;
        RECT 161.100 883.050 162.900 884.850 ;
        RECT 164.100 883.050 165.300 890.400 ;
        RECT 167.700 886.800 168.900 890.400 ;
        RECT 178.800 889.500 180.300 890.400 ;
        RECT 187.800 889.800 189.600 890.400 ;
        RECT 191.700 889.800 192.600 890.400 ;
        RECT 171.900 888.300 180.300 889.500 ;
        RECT 185.400 888.600 192.600 889.800 ;
        RECT 207.300 888.600 213.900 890.400 ;
        RECT 171.900 887.700 173.700 888.300 ;
        RECT 182.400 886.800 184.500 887.700 ;
        RECT 167.700 885.600 184.500 886.800 ;
        RECT 185.400 885.600 186.300 888.600 ;
        RECT 190.800 885.900 192.600 886.800 ;
        RECT 200.100 886.500 201.900 888.300 ;
        RECT 218.100 887.100 219.600 890.400 ;
        RECT 193.800 885.900 195.900 886.050 ;
        RECT 115.500 880.950 117.600 883.050 ;
        RECT 118.800 880.950 120.900 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 142.950 880.950 145.050 883.050 ;
        RECT 160.950 880.950 163.050 883.050 ;
        RECT 163.950 880.950 166.050 883.050 ;
        RECT 115.200 879.150 117.000 880.950 ;
        RECT 113.100 876.300 114.900 876.900 ;
        RECT 113.100 875.100 120.900 876.300 ;
        RECT 119.700 873.600 120.900 875.100 ;
        RECT 111.000 872.100 113.400 873.600 ;
        RECT 58.200 861.000 60.000 867.600 ;
        RECT 61.200 861.600 63.000 867.600 ;
        RECT 64.200 864.600 66.300 866.700 ;
        RECT 67.200 864.600 69.300 866.700 ;
        RECT 70.200 864.600 72.300 866.700 ;
        RECT 64.200 861.600 66.000 864.600 ;
        RECT 67.200 861.600 69.000 864.600 ;
        RECT 70.200 861.600 72.000 864.600 ;
        RECT 73.200 861.000 75.000 867.600 ;
        RECT 76.200 861.600 78.000 867.600 ;
        RECT 79.200 861.000 81.000 867.600 ;
        RECT 82.200 861.600 84.000 867.600 ;
        RECT 85.200 861.000 87.000 867.600 ;
        RECT 88.500 861.600 90.300 867.600 ;
        RECT 91.500 861.000 93.300 867.600 ;
        RECT 111.600 861.600 113.400 872.100 ;
        RECT 114.600 861.000 116.400 873.600 ;
        RECT 119.100 861.600 120.900 873.600 ;
        RECT 140.700 867.600 141.900 880.950 ;
        RECT 164.100 873.600 165.300 880.950 ;
        RECT 137.100 861.000 138.900 867.600 ;
        RECT 140.100 861.600 141.900 867.600 ;
        RECT 143.100 861.000 144.900 867.600 ;
        RECT 161.100 861.000 162.900 873.600 ;
        RECT 164.100 861.600 165.900 873.600 ;
        RECT 167.700 869.400 168.900 885.600 ;
        RECT 185.400 883.800 187.200 885.600 ;
        RECT 190.800 885.000 195.900 885.900 ;
        RECT 193.800 883.950 195.900 885.000 ;
        RECT 200.100 885.900 202.200 886.500 ;
        RECT 200.100 884.400 217.200 885.900 ;
        RECT 218.100 885.300 225.900 887.100 ;
        RECT 215.700 882.900 222.300 884.400 ;
        RECT 170.100 881.700 214.500 882.900 ;
        RECT 170.100 880.050 171.900 881.700 ;
        RECT 169.800 877.950 171.900 880.050 ;
        RECT 175.800 879.750 177.900 880.050 ;
        RECT 188.400 879.900 190.200 880.500 ;
        RECT 197.400 879.900 210.900 880.800 ;
        RECT 175.800 877.950 179.700 879.750 ;
        RECT 188.400 878.700 199.500 879.900 ;
        RECT 177.900 877.200 179.700 877.950 ;
        RECT 197.400 877.800 199.500 878.700 ;
        RECT 201.000 877.200 204.900 879.000 ;
        RECT 210.000 878.700 210.900 879.900 ;
        RECT 177.900 876.300 191.400 877.200 ;
        RECT 202.800 876.900 204.900 877.200 ;
        RECT 209.100 876.900 210.900 878.700 ;
        RECT 213.600 880.200 214.500 881.700 ;
        RECT 213.600 878.400 218.700 880.200 ;
        RECT 220.800 880.050 222.300 882.900 ;
        RECT 220.800 877.950 222.900 880.050 ;
        RECT 190.200 875.700 191.400 876.300 ;
        RECT 224.100 875.700 225.900 876.300 ;
        RECT 185.400 874.500 187.500 874.800 ;
        RECT 190.200 874.500 225.900 875.700 ;
        RECT 175.500 873.300 187.500 874.500 ;
        RECT 226.800 873.600 227.700 890.400 ;
        RECT 175.500 872.700 177.300 873.300 ;
        RECT 185.400 872.700 187.500 873.300 ;
        RECT 190.200 872.400 207.900 873.600 ;
        RECT 172.200 871.800 174.000 872.100 ;
        RECT 190.200 871.800 191.400 872.400 ;
        RECT 172.200 870.600 191.400 871.800 ;
        RECT 205.800 871.500 207.900 872.400 ;
        RECT 211.200 872.700 227.700 873.600 ;
        RECT 211.200 871.500 213.300 872.700 ;
        RECT 172.200 870.300 174.000 870.600 ;
        RECT 167.700 868.500 171.300 869.400 ;
        RECT 170.400 867.600 171.300 868.500 ;
        RECT 167.700 861.000 169.500 867.600 ;
        RECT 170.400 866.700 172.500 867.600 ;
        RECT 170.700 861.600 172.500 866.700 ;
        RECT 173.700 861.000 175.500 867.600 ;
        RECT 176.700 861.600 178.500 870.600 ;
        RECT 188.700 867.600 190.800 869.700 ;
        RECT 196.200 869.100 199.500 871.200 ;
        RECT 179.700 861.000 181.500 867.600 ;
        RECT 183.300 864.600 185.400 866.700 ;
        RECT 186.300 864.600 188.400 866.700 ;
        RECT 183.300 861.600 185.100 864.600 ;
        RECT 186.300 861.600 188.100 864.600 ;
        RECT 189.300 861.600 191.100 867.600 ;
        RECT 192.300 861.000 194.100 867.600 ;
        RECT 196.200 861.600 198.000 869.100 ;
        RECT 202.200 867.600 204.900 871.500 ;
        RECT 217.200 870.600 222.900 871.800 ;
        RECT 214.500 869.700 216.300 870.300 ;
        RECT 208.200 868.500 216.300 869.700 ;
        RECT 208.200 867.600 210.300 868.500 ;
        RECT 217.200 867.600 218.400 870.600 ;
        RECT 221.100 870.000 222.900 870.600 ;
        RECT 226.800 869.400 227.700 872.700 ;
        RECT 223.800 868.500 227.700 869.400 ;
        RECT 229.500 893.400 231.300 896.400 ;
        RECT 232.500 893.400 234.300 897.000 ;
        RECT 229.500 880.050 231.000 893.400 ;
        RECT 251.100 891.300 252.900 896.400 ;
        RECT 254.100 892.200 255.900 897.000 ;
        RECT 257.100 891.300 258.900 896.400 ;
        RECT 251.100 889.950 258.900 891.300 ;
        RECT 260.100 890.400 261.900 896.400 ;
        RECT 278.100 891.300 279.900 896.400 ;
        RECT 281.100 892.200 282.900 897.000 ;
        RECT 284.100 891.300 285.900 896.400 ;
        RECT 260.100 888.300 261.300 890.400 ;
        RECT 278.100 889.950 285.900 891.300 ;
        RECT 287.100 890.400 288.900 896.400 ;
        RECT 305.100 893.400 306.900 897.000 ;
        RECT 308.100 893.400 309.900 896.400 ;
        RECT 287.100 888.300 288.300 890.400 ;
        RECT 257.700 887.400 261.300 888.300 ;
        RECT 284.700 887.400 288.300 888.300 ;
        RECT 254.100 883.050 255.900 884.850 ;
        RECT 257.700 883.050 258.900 887.400 ;
        RECT 260.100 883.050 261.900 884.850 ;
        RECT 281.100 883.050 282.900 884.850 ;
        RECT 284.700 883.050 285.900 887.400 ;
        RECT 287.100 883.050 288.900 884.850 ;
        RECT 308.100 883.050 309.300 893.400 ;
        RECT 326.100 891.300 327.900 896.400 ;
        RECT 329.100 892.200 330.900 897.000 ;
        RECT 332.100 891.300 333.900 896.400 ;
        RECT 326.100 889.950 333.900 891.300 ;
        RECT 335.100 890.400 336.900 896.400 ;
        RECT 353.100 890.400 354.900 896.400 ;
        RECT 335.100 888.300 336.300 890.400 ;
        RECT 332.700 887.400 336.300 888.300 ;
        RECT 353.700 888.300 354.900 890.400 ;
        RECT 356.100 891.300 357.900 896.400 ;
        RECT 359.100 892.200 360.900 897.000 ;
        RECT 362.100 891.300 363.900 896.400 ;
        RECT 356.100 889.950 363.900 891.300 ;
        RECT 353.700 887.400 357.300 888.300 ;
        RECT 382.500 888.000 384.300 896.400 ;
        RECT 329.100 883.050 330.900 884.850 ;
        RECT 332.700 883.050 333.900 887.400 ;
        RECT 335.100 883.050 336.900 884.850 ;
        RECT 353.100 883.050 354.900 884.850 ;
        RECT 356.100 883.050 357.300 887.400 ;
        RECT 381.000 886.800 384.300 888.000 ;
        RECT 389.100 887.400 390.900 897.000 ;
        RECT 407.100 891.300 408.900 896.400 ;
        RECT 410.100 892.200 411.900 897.000 ;
        RECT 413.100 891.300 414.900 896.400 ;
        RECT 407.100 889.950 414.900 891.300 ;
        RECT 416.100 890.400 417.900 896.400 ;
        RECT 431.100 890.400 432.900 896.400 ;
        RECT 416.100 888.300 417.300 890.400 ;
        RECT 413.700 887.400 417.300 888.300 ;
        RECT 431.700 888.300 432.900 890.400 ;
        RECT 434.100 891.300 435.900 896.400 ;
        RECT 437.100 892.200 438.900 897.000 ;
        RECT 440.100 891.300 441.900 896.400 ;
        RECT 458.100 893.400 459.900 896.400 ;
        RECT 461.100 893.400 462.900 897.000 ;
        RECT 434.100 889.950 441.900 891.300 ;
        RECT 431.700 887.400 435.300 888.300 ;
        RECT 359.100 883.050 360.900 884.850 ;
        RECT 381.000 883.050 381.900 886.800 ;
        RECT 383.100 883.050 384.900 884.850 ;
        RECT 389.100 883.050 390.900 884.850 ;
        RECT 410.100 883.050 411.900 884.850 ;
        RECT 413.700 883.050 414.900 887.400 ;
        RECT 416.100 883.050 417.900 884.850 ;
        RECT 431.100 883.050 432.900 884.850 ;
        RECT 434.100 883.050 435.300 887.400 ;
        RECT 445.950 885.450 448.050 886.050 ;
        RECT 454.950 885.450 457.050 886.050 ;
        RECT 437.100 883.050 438.900 884.850 ;
        RECT 445.950 884.550 457.050 885.450 ;
        RECT 445.950 883.950 448.050 884.550 ;
        RECT 454.950 883.950 457.050 884.550 ;
        RECT 458.700 883.050 459.900 893.400 ;
        RECT 479.700 889.200 481.500 896.400 ;
        RECT 484.800 890.400 486.600 897.000 ;
        RECT 503.100 893.400 504.900 897.000 ;
        RECT 506.100 893.400 507.900 896.400 ;
        RECT 509.100 893.400 510.900 897.000 ;
        RECT 524.100 893.400 525.900 897.000 ;
        RECT 527.100 893.400 528.900 896.400 ;
        RECT 530.100 893.400 531.900 897.000 ;
        RECT 479.700 888.300 483.900 889.200 ;
        RECT 479.100 883.050 480.900 884.850 ;
        RECT 482.700 883.050 483.900 888.300 ;
        RECT 490.950 885.450 493.050 886.050 ;
        RECT 499.950 885.450 502.050 886.050 ;
        RECT 484.950 883.050 486.750 884.850 ;
        RECT 490.950 884.550 502.050 885.450 ;
        RECT 490.950 883.950 493.050 884.550 ;
        RECT 499.950 883.950 502.050 884.550 ;
        RECT 506.400 883.050 507.300 893.400 ;
        RECT 508.950 888.450 511.050 888.900 ;
        RECT 517.950 888.450 520.050 889.050 ;
        RECT 508.950 887.550 520.050 888.450 ;
        RECT 508.950 886.800 511.050 887.550 ;
        RECT 517.950 886.950 520.050 887.550 ;
        RECT 511.950 885.450 516.000 886.050 ;
        RECT 511.950 883.950 516.450 885.450 ;
        RECT 232.950 882.450 235.050 883.050 ;
        RECT 244.950 882.450 247.050 883.050 ;
        RECT 232.950 881.550 247.050 882.450 ;
        RECT 232.950 880.950 235.050 881.550 ;
        RECT 244.950 880.950 247.050 881.550 ;
        RECT 250.950 880.950 253.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 277.950 880.950 280.050 883.050 ;
        RECT 280.950 880.950 283.050 883.050 ;
        RECT 283.950 880.950 286.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 304.950 880.950 307.050 883.050 ;
        RECT 307.950 880.950 310.050 883.050 ;
        RECT 325.950 880.950 328.050 883.050 ;
        RECT 328.950 880.950 331.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 361.950 880.950 364.050 883.050 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 382.950 880.950 385.050 883.050 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 430.950 880.950 433.050 883.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 481.950 880.950 484.050 883.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 502.950 880.950 505.050 883.050 ;
        RECT 505.950 880.950 508.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 229.500 877.950 231.900 880.050 ;
        RECT 251.100 879.150 252.900 880.950 ;
        RECT 223.800 867.600 225.000 868.500 ;
        RECT 229.500 867.600 231.000 877.950 ;
        RECT 257.700 873.600 258.900 880.950 ;
        RECT 278.100 879.150 279.900 880.950 ;
        RECT 284.700 873.600 285.900 880.950 ;
        RECT 305.100 879.150 306.900 880.950 ;
        RECT 199.200 861.000 201.000 867.600 ;
        RECT 202.200 861.600 204.000 867.600 ;
        RECT 205.200 864.600 207.300 866.700 ;
        RECT 208.200 864.600 210.300 866.700 ;
        RECT 211.200 864.600 213.300 866.700 ;
        RECT 205.200 861.600 207.000 864.600 ;
        RECT 208.200 861.600 210.000 864.600 ;
        RECT 211.200 861.600 213.000 864.600 ;
        RECT 214.200 861.000 216.000 867.600 ;
        RECT 217.200 861.600 219.000 867.600 ;
        RECT 220.200 861.000 222.000 867.600 ;
        RECT 223.200 861.600 225.000 867.600 ;
        RECT 226.200 861.000 228.000 867.600 ;
        RECT 229.500 861.600 231.300 867.600 ;
        RECT 232.500 861.000 234.300 867.600 ;
        RECT 251.400 861.000 253.200 873.600 ;
        RECT 256.500 872.100 258.900 873.600 ;
        RECT 256.500 861.600 258.300 872.100 ;
        RECT 259.200 869.100 261.000 870.900 ;
        RECT 259.500 861.000 261.300 867.600 ;
        RECT 278.400 861.000 280.200 873.600 ;
        RECT 283.500 872.100 285.900 873.600 ;
        RECT 283.500 861.600 285.300 872.100 ;
        RECT 286.200 869.100 288.000 870.900 ;
        RECT 308.100 867.600 309.300 880.950 ;
        RECT 326.100 879.150 327.900 880.950 ;
        RECT 332.700 873.600 333.900 880.950 ;
        RECT 286.500 861.000 288.300 867.600 ;
        RECT 305.100 861.000 306.900 867.600 ;
        RECT 308.100 861.600 309.900 867.600 ;
        RECT 326.400 861.000 328.200 873.600 ;
        RECT 331.500 872.100 333.900 873.600 ;
        RECT 356.100 873.600 357.300 880.950 ;
        RECT 362.100 879.150 363.900 880.950 ;
        RECT 356.100 872.100 358.500 873.600 ;
        RECT 331.500 861.600 333.300 872.100 ;
        RECT 334.200 869.100 336.000 870.900 ;
        RECT 354.000 869.100 355.800 870.900 ;
        RECT 334.500 861.000 336.300 867.600 ;
        RECT 353.700 861.000 355.500 867.600 ;
        RECT 356.700 861.600 358.500 872.100 ;
        RECT 361.800 861.000 363.600 873.600 ;
        RECT 381.000 868.800 381.900 880.950 ;
        RECT 386.100 879.150 387.900 880.950 ;
        RECT 407.100 879.150 408.900 880.950 ;
        RECT 413.700 873.600 414.900 880.950 ;
        RECT 381.000 867.900 387.600 868.800 ;
        RECT 381.000 867.600 381.900 867.900 ;
        RECT 380.100 861.600 381.900 867.600 ;
        RECT 386.100 867.600 387.600 867.900 ;
        RECT 383.100 861.000 384.900 867.000 ;
        RECT 386.100 861.600 387.900 867.600 ;
        RECT 389.100 861.000 390.900 867.600 ;
        RECT 407.400 861.000 409.200 873.600 ;
        RECT 412.500 872.100 414.900 873.600 ;
        RECT 434.100 873.600 435.300 880.950 ;
        RECT 440.100 879.150 441.900 880.950 ;
        RECT 434.100 872.100 436.500 873.600 ;
        RECT 412.500 861.600 414.300 872.100 ;
        RECT 415.200 869.100 417.000 870.900 ;
        RECT 432.000 869.100 433.800 870.900 ;
        RECT 415.500 861.000 417.300 867.600 ;
        RECT 431.700 861.000 433.500 867.600 ;
        RECT 434.700 861.600 436.500 872.100 ;
        RECT 439.800 861.000 441.600 873.600 ;
        RECT 458.700 867.600 459.900 880.950 ;
        RECT 461.100 879.150 462.900 880.950 ;
        RECT 482.700 867.600 483.900 880.950 ;
        RECT 503.250 879.150 505.050 880.950 ;
        RECT 506.400 873.600 507.300 880.950 ;
        RECT 509.100 879.150 510.900 880.950 ;
        RECT 515.550 880.050 516.450 883.950 ;
        RECT 527.700 883.050 528.600 893.400 ;
        RECT 548.100 887.400 549.900 897.000 ;
        RECT 554.700 888.000 556.500 896.400 ;
        RECT 575.400 890.400 577.200 897.000 ;
        RECT 580.500 889.200 582.300 896.400 ;
        RECT 599.700 893.400 601.500 897.000 ;
        RECT 602.700 891.600 604.500 896.400 ;
        RECT 578.100 888.300 582.300 889.200 ;
        RECT 599.400 890.400 604.500 891.600 ;
        RECT 607.200 890.400 609.000 897.000 ;
        RECT 626.100 893.400 627.900 897.000 ;
        RECT 629.100 893.400 630.900 896.400 ;
        RECT 632.100 893.400 633.900 897.000 ;
        RECT 554.700 886.800 558.000 888.000 ;
        RECT 548.100 883.050 549.900 884.850 ;
        RECT 554.100 883.050 555.900 884.850 ;
        RECT 557.100 883.050 558.000 886.800 ;
        RECT 575.250 883.050 577.050 884.850 ;
        RECT 578.100 883.050 579.300 888.300 ;
        RECT 581.100 883.050 582.900 884.850 ;
        RECT 599.400 883.050 600.300 890.400 ;
        RECT 601.950 883.050 603.750 884.850 ;
        RECT 608.100 883.050 609.900 884.850 ;
        RECT 629.400 883.050 630.300 893.400 ;
        RECT 650.100 891.000 651.900 896.400 ;
        RECT 653.100 891.900 654.900 897.000 ;
        RECT 656.100 895.500 663.900 896.400 ;
        RECT 656.100 891.000 657.900 895.500 ;
        RECT 650.100 890.100 657.900 891.000 ;
        RECT 659.100 890.400 660.900 894.600 ;
        RECT 662.100 890.400 663.900 895.500 ;
        RECT 680.100 893.400 681.900 897.000 ;
        RECT 683.100 893.400 684.900 896.400 ;
        RECT 686.100 893.400 687.900 897.000 ;
        RECT 704.100 893.400 705.900 897.000 ;
        RECT 707.100 893.400 708.900 896.400 ;
        RECT 710.100 893.400 711.900 897.000 ;
        RECT 659.400 888.900 660.300 890.400 ;
        RECT 655.950 887.700 660.300 888.900 ;
        RECT 634.950 885.450 637.050 886.050 ;
        RECT 640.950 885.450 643.050 886.050 ;
        RECT 634.950 884.550 643.050 885.450 ;
        RECT 634.950 883.950 637.050 884.550 ;
        RECT 640.950 883.950 643.050 884.550 ;
        RECT 653.250 883.050 655.050 884.850 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 529.950 880.950 532.050 883.050 ;
        RECT 547.950 880.950 550.050 883.050 ;
        RECT 550.950 880.950 553.050 883.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 604.950 880.950 607.050 883.050 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 652.950 880.950 655.050 883.050 ;
        RECT 655.950 883.050 657.000 887.700 ;
        RECT 658.950 883.050 660.750 884.850 ;
        RECT 683.400 883.050 684.300 893.400 ;
        RECT 691.950 891.450 694.050 892.050 ;
        RECT 703.950 891.450 706.050 892.050 ;
        RECT 691.950 890.550 706.050 891.450 ;
        RECT 691.950 889.950 694.050 890.550 ;
        RECT 703.950 889.950 706.050 890.550 ;
        RECT 707.400 883.050 708.300 893.400 ;
        RECT 728.700 889.200 730.500 896.400 ;
        RECT 733.800 890.400 735.600 897.000 ;
        RECT 739.950 894.450 742.050 895.050 ;
        RECT 748.950 894.450 751.050 895.050 ;
        RECT 739.950 893.550 751.050 894.450 ;
        RECT 739.950 892.950 742.050 893.550 ;
        RECT 748.950 892.950 751.050 893.550 ;
        RECT 728.700 888.300 732.900 889.200 ;
        RECT 728.100 883.050 729.900 884.850 ;
        RECT 731.700 883.050 732.900 888.300 ;
        RECT 754.500 888.000 756.300 896.400 ;
        RECT 753.000 886.800 756.300 888.000 ;
        RECT 761.100 887.400 762.900 897.000 ;
        RECT 769.950 891.450 772.050 892.050 ;
        RECT 775.950 891.450 778.050 892.050 ;
        RECT 769.950 890.550 778.050 891.450 ;
        RECT 769.950 889.950 772.050 890.550 ;
        RECT 775.950 889.950 778.050 890.550 ;
        RECT 779.100 890.400 780.900 896.400 ;
        RECT 779.700 888.300 780.900 890.400 ;
        RECT 782.100 891.300 783.900 896.400 ;
        RECT 785.100 892.200 786.900 897.000 ;
        RECT 788.100 891.300 789.900 896.400 ;
        RECT 782.100 889.950 789.900 891.300 ;
        RECT 779.700 887.400 783.300 888.300 ;
        RECT 806.100 887.400 807.900 897.000 ;
        RECT 812.700 888.000 814.500 896.400 ;
        RECT 834.000 890.400 835.800 897.000 ;
        RECT 838.500 891.600 840.300 896.400 ;
        RECT 841.500 893.400 843.300 897.000 ;
        RECT 838.500 890.400 843.600 891.600 ;
        RECT 733.950 883.050 735.750 884.850 ;
        RECT 753.000 883.050 753.900 886.800 ;
        RECT 755.100 883.050 756.900 884.850 ;
        RECT 761.100 883.050 762.900 884.850 ;
        RECT 779.100 883.050 780.900 884.850 ;
        RECT 782.100 883.050 783.300 887.400 ;
        RECT 812.700 886.800 816.000 888.000 ;
        RECT 785.100 883.050 786.900 884.850 ;
        RECT 806.100 883.050 807.900 884.850 ;
        RECT 812.100 883.050 813.900 884.850 ;
        RECT 815.100 883.050 816.000 886.800 ;
        RECT 833.100 883.050 834.900 884.850 ;
        RECT 839.250 883.050 841.050 884.850 ;
        RECT 842.700 883.050 843.600 890.400 ;
        RECT 857.700 889.200 859.500 896.400 ;
        RECT 862.800 890.400 864.600 897.000 ;
        RECT 857.700 888.300 861.900 889.200 ;
        RECT 857.100 883.050 858.900 884.850 ;
        RECT 860.700 883.050 861.900 888.300 ;
        RECT 881.100 888.600 882.900 896.400 ;
        RECT 885.600 890.400 887.400 897.000 ;
        RECT 888.600 892.200 890.400 896.400 ;
        RECT 888.600 890.400 891.300 892.200 ;
        RECT 887.700 888.600 889.500 889.500 ;
        RECT 881.100 887.700 889.500 888.600 ;
        RECT 862.950 883.050 864.750 884.850 ;
        RECT 881.250 883.050 883.050 884.850 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 881.100 880.950 883.200 883.050 ;
        RECT 511.950 878.550 516.450 880.050 ;
        RECT 524.100 879.150 525.900 880.950 ;
        RECT 511.950 877.950 516.000 878.550 ;
        RECT 527.700 873.600 528.600 880.950 ;
        RECT 529.950 879.150 531.750 880.950 ;
        RECT 551.100 879.150 552.900 880.950 ;
        RECT 529.950 876.450 532.050 877.050 ;
        RECT 553.950 876.450 556.050 877.050 ;
        RECT 529.950 875.550 556.050 876.450 ;
        RECT 529.950 874.950 532.050 875.550 ;
        RECT 553.950 874.950 556.050 875.550 ;
        RECT 458.100 861.600 459.900 867.600 ;
        RECT 461.100 861.000 462.900 867.600 ;
        RECT 479.100 861.000 480.900 867.600 ;
        RECT 482.100 861.600 483.900 867.600 ;
        RECT 485.100 861.000 486.900 867.600 ;
        RECT 503.100 861.000 504.900 873.600 ;
        RECT 506.400 872.400 510.000 873.600 ;
        RECT 508.200 861.600 510.000 872.400 ;
        RECT 525.000 872.400 528.600 873.600 ;
        RECT 525.000 861.600 526.800 872.400 ;
        RECT 530.100 861.000 531.900 873.600 ;
        RECT 557.100 868.800 558.000 880.950 ;
        RECT 551.400 867.900 558.000 868.800 ;
        RECT 551.400 867.600 552.900 867.900 ;
        RECT 548.100 861.000 549.900 867.600 ;
        RECT 551.100 861.600 552.900 867.600 ;
        RECT 557.100 867.600 558.000 867.900 ;
        RECT 578.100 867.600 579.300 880.950 ;
        RECT 580.950 876.450 583.050 877.050 ;
        RECT 589.950 876.450 592.050 877.050 ;
        RECT 580.950 875.550 592.050 876.450 ;
        RECT 580.950 874.950 583.050 875.550 ;
        RECT 589.950 874.950 592.050 875.550 ;
        RECT 599.400 873.600 600.300 880.950 ;
        RECT 604.950 879.150 606.750 880.950 ;
        RECT 626.250 879.150 628.050 880.950 ;
        RECT 601.950 876.450 604.050 877.050 ;
        RECT 613.950 876.450 616.050 877.050 ;
        RECT 601.950 875.550 616.050 876.450 ;
        RECT 601.950 874.950 604.050 875.550 ;
        RECT 613.950 874.950 616.050 875.550 ;
        RECT 629.400 873.600 630.300 880.950 ;
        RECT 632.100 879.150 633.900 880.950 ;
        RECT 650.100 879.150 651.900 880.950 ;
        RECT 631.950 876.450 634.050 877.050 ;
        RECT 649.950 876.450 652.050 877.050 ;
        RECT 631.950 875.550 652.050 876.450 ;
        RECT 631.950 874.950 634.050 875.550 ;
        RECT 649.950 874.950 652.050 875.550 ;
        RECT 655.950 873.600 657.000 880.950 ;
        RECT 661.950 879.150 663.750 880.950 ;
        RECT 680.250 879.150 682.050 880.950 ;
        RECT 683.400 873.600 684.300 880.950 ;
        RECT 686.100 879.150 687.900 880.950 ;
        RECT 704.250 879.150 706.050 880.950 ;
        RECT 685.950 876.450 688.050 877.050 ;
        RECT 703.950 876.450 706.050 877.050 ;
        RECT 685.950 875.550 706.050 876.450 ;
        RECT 685.950 874.950 688.050 875.550 ;
        RECT 703.950 874.950 706.050 875.550 ;
        RECT 707.400 873.600 708.300 880.950 ;
        RECT 710.100 879.150 711.900 880.950 ;
        RECT 715.950 879.450 718.050 880.050 ;
        RECT 724.950 879.450 727.050 880.050 ;
        RECT 715.950 878.550 727.050 879.450 ;
        RECT 715.950 877.950 718.050 878.550 ;
        RECT 724.950 877.950 727.050 878.550 ;
        RECT 554.100 861.000 555.900 867.000 ;
        RECT 557.100 861.600 558.900 867.600 ;
        RECT 575.100 861.000 576.900 867.600 ;
        RECT 578.100 861.600 579.900 867.600 ;
        RECT 581.100 861.000 582.900 867.600 ;
        RECT 599.100 861.600 600.900 873.600 ;
        RECT 602.100 872.700 609.900 873.600 ;
        RECT 602.100 861.600 603.900 872.700 ;
        RECT 605.100 861.000 606.900 871.800 ;
        RECT 608.100 861.600 609.900 872.700 ;
        RECT 626.100 861.000 627.900 873.600 ;
        RECT 629.400 872.400 633.000 873.600 ;
        RECT 631.200 861.600 633.000 872.400 ;
        RECT 650.100 861.000 651.900 873.600 ;
        RECT 654.600 861.600 657.900 873.600 ;
        RECT 660.600 861.000 662.400 873.600 ;
        RECT 680.100 861.000 681.900 873.600 ;
        RECT 683.400 872.400 687.000 873.600 ;
        RECT 685.200 861.600 687.000 872.400 ;
        RECT 704.100 861.000 705.900 873.600 ;
        RECT 707.400 872.400 711.000 873.600 ;
        RECT 709.200 861.600 711.000 872.400 ;
        RECT 731.700 867.600 732.900 880.950 ;
        RECT 753.000 868.800 753.900 880.950 ;
        RECT 758.100 879.150 759.900 880.950 ;
        RECT 782.100 873.600 783.300 880.950 ;
        RECT 788.100 879.150 789.900 880.950 ;
        RECT 809.100 879.150 810.900 880.950 ;
        RECT 784.950 876.450 787.050 877.050 ;
        RECT 790.800 876.450 792.900 877.050 ;
        RECT 784.950 875.550 792.900 876.450 ;
        RECT 784.950 874.950 787.050 875.550 ;
        RECT 790.800 874.950 792.900 875.550 ;
        RECT 793.950 876.450 796.050 877.050 ;
        RECT 805.950 876.450 808.050 877.050 ;
        RECT 793.950 875.550 808.050 876.450 ;
        RECT 793.950 874.950 796.050 875.550 ;
        RECT 805.950 874.950 808.050 875.550 ;
        RECT 782.100 872.100 784.500 873.600 ;
        RECT 780.000 869.100 781.800 870.900 ;
        RECT 753.000 867.900 759.600 868.800 ;
        RECT 753.000 867.600 753.900 867.900 ;
        RECT 728.100 861.000 729.900 867.600 ;
        RECT 731.100 861.600 732.900 867.600 ;
        RECT 734.100 861.000 735.900 867.600 ;
        RECT 752.100 861.600 753.900 867.600 ;
        RECT 758.100 867.600 759.600 867.900 ;
        RECT 755.100 861.000 756.900 867.000 ;
        RECT 758.100 861.600 759.900 867.600 ;
        RECT 761.100 861.000 762.900 867.600 ;
        RECT 779.700 861.000 781.500 867.600 ;
        RECT 782.700 861.600 784.500 872.100 ;
        RECT 787.800 861.000 789.600 873.600 ;
        RECT 815.100 868.800 816.000 880.950 ;
        RECT 836.250 879.150 838.050 880.950 ;
        RECT 842.700 873.600 843.600 880.950 ;
        RECT 793.950 867.450 796.050 868.050 ;
        RECT 809.400 867.900 816.000 868.800 ;
        RECT 799.950 867.450 802.050 867.900 ;
        RECT 809.400 867.600 810.900 867.900 ;
        RECT 793.950 866.550 802.050 867.450 ;
        RECT 793.950 865.950 796.050 866.550 ;
        RECT 799.950 865.800 802.050 866.550 ;
        RECT 806.100 861.000 807.900 867.600 ;
        RECT 809.100 861.600 810.900 867.600 ;
        RECT 815.100 867.600 816.000 867.900 ;
        RECT 833.100 872.700 840.900 873.600 ;
        RECT 812.100 861.000 813.900 867.000 ;
        RECT 815.100 861.600 816.900 867.600 ;
        RECT 833.100 861.600 834.900 872.700 ;
        RECT 836.100 861.000 837.900 871.800 ;
        RECT 839.100 861.600 840.900 872.700 ;
        RECT 842.100 861.600 843.900 873.600 ;
        RECT 860.700 867.600 861.900 880.950 ;
        RECT 884.100 867.600 885.000 887.700 ;
        RECT 890.400 883.050 891.300 890.400 ;
        RECT 908.100 887.400 909.900 897.000 ;
        RECT 914.700 888.000 916.500 896.400 ;
        RECT 937.500 888.000 939.300 896.400 ;
        RECT 914.700 886.800 918.000 888.000 ;
        RECT 908.100 883.050 909.900 884.850 ;
        RECT 914.100 883.050 915.900 884.850 ;
        RECT 917.100 883.050 918.000 886.800 ;
        RECT 936.000 886.800 939.300 888.000 ;
        RECT 944.100 887.400 945.900 897.000 ;
        RECT 962.100 887.400 963.900 897.000 ;
        RECT 968.700 888.000 970.500 896.400 ;
        RECT 989.100 888.600 990.900 896.400 ;
        RECT 993.600 890.400 995.400 897.000 ;
        RECT 996.600 892.200 998.400 896.400 ;
        RECT 996.600 890.400 999.300 892.200 ;
        RECT 995.700 888.600 997.500 889.500 ;
        RECT 968.700 886.800 972.000 888.000 ;
        RECT 989.100 887.700 997.500 888.600 ;
        RECT 936.000 883.050 936.900 886.800 ;
        RECT 938.100 883.050 939.900 884.850 ;
        RECT 944.100 883.050 945.900 884.850 ;
        RECT 962.100 883.050 963.900 884.850 ;
        RECT 968.100 883.050 969.900 884.850 ;
        RECT 971.100 883.050 972.000 886.800 ;
        RECT 989.250 883.050 991.050 884.850 ;
        RECT 886.500 880.950 888.600 883.050 ;
        RECT 889.800 880.950 891.900 883.050 ;
        RECT 907.950 880.950 910.050 883.050 ;
        RECT 910.950 880.950 913.050 883.050 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 934.950 880.950 937.050 883.050 ;
        RECT 937.950 880.950 940.050 883.050 ;
        RECT 940.950 880.950 943.050 883.050 ;
        RECT 943.950 880.950 946.050 883.050 ;
        RECT 961.950 880.950 964.050 883.050 ;
        RECT 964.950 880.950 967.050 883.050 ;
        RECT 967.950 880.950 970.050 883.050 ;
        RECT 970.950 880.950 973.050 883.050 ;
        RECT 989.100 880.950 991.200 883.050 ;
        RECT 886.200 879.150 888.000 880.950 ;
        RECT 890.400 873.600 891.300 880.950 ;
        RECT 911.100 879.150 912.900 880.950 ;
        RECT 892.950 876.450 895.050 877.050 ;
        RECT 907.950 876.450 910.050 877.050 ;
        RECT 892.950 875.550 910.050 876.450 ;
        RECT 892.950 874.950 895.050 875.550 ;
        RECT 907.950 874.950 910.050 875.550 ;
        RECT 857.100 861.000 858.900 867.600 ;
        RECT 860.100 861.600 861.900 867.600 ;
        RECT 863.100 861.000 864.900 867.600 ;
        RECT 881.100 861.000 882.900 867.600 ;
        RECT 884.100 861.600 885.900 867.600 ;
        RECT 887.100 861.000 888.900 873.000 ;
        RECT 890.100 861.600 891.900 873.600 ;
        RECT 917.100 868.800 918.000 880.950 ;
        RECT 911.400 867.900 918.000 868.800 ;
        RECT 911.400 867.600 912.900 867.900 ;
        RECT 908.100 861.000 909.900 867.600 ;
        RECT 911.100 861.600 912.900 867.600 ;
        RECT 917.100 867.600 918.000 867.900 ;
        RECT 936.000 868.800 936.900 880.950 ;
        RECT 941.100 879.150 942.900 880.950 ;
        RECT 965.100 879.150 966.900 880.950 ;
        RECT 949.950 873.450 952.050 874.050 ;
        RECT 967.950 873.450 970.050 874.050 ;
        RECT 949.950 872.550 970.050 873.450 ;
        RECT 949.950 871.950 952.050 872.550 ;
        RECT 967.950 871.950 970.050 872.550 ;
        RECT 943.950 870.450 946.050 871.050 ;
        RECT 961.950 870.450 964.050 871.050 ;
        RECT 943.950 869.550 964.050 870.450 ;
        RECT 943.950 868.950 946.050 869.550 ;
        RECT 961.950 868.950 964.050 869.550 ;
        RECT 971.100 868.800 972.000 880.950 ;
        RECT 976.950 876.450 979.050 877.050 ;
        RECT 988.950 876.450 991.050 877.050 ;
        RECT 976.950 875.550 991.050 876.450 ;
        RECT 976.950 874.950 979.050 875.550 ;
        RECT 988.950 874.950 991.050 875.550 ;
        RECT 936.000 867.900 942.600 868.800 ;
        RECT 936.000 867.600 936.900 867.900 ;
        RECT 914.100 861.000 915.900 867.000 ;
        RECT 917.100 861.600 918.900 867.600 ;
        RECT 935.100 861.600 936.900 867.600 ;
        RECT 941.100 867.600 942.600 867.900 ;
        RECT 965.400 867.900 972.000 868.800 ;
        RECT 965.400 867.600 966.900 867.900 ;
        RECT 938.100 861.000 939.900 867.000 ;
        RECT 941.100 861.600 942.900 867.600 ;
        RECT 944.100 861.000 945.900 867.600 ;
        RECT 962.100 861.000 963.900 867.600 ;
        RECT 965.100 861.600 966.900 867.600 ;
        RECT 971.100 867.600 972.000 867.900 ;
        RECT 992.100 867.600 993.000 887.700 ;
        RECT 998.400 883.050 999.300 890.400 ;
        RECT 1016.700 889.200 1018.500 896.400 ;
        RECT 1021.800 890.400 1023.600 897.000 ;
        RECT 1016.700 888.300 1020.900 889.200 ;
        RECT 1016.100 883.050 1017.900 884.850 ;
        RECT 1019.700 883.050 1020.900 888.300 ;
        RECT 1021.950 883.050 1023.750 884.850 ;
        RECT 994.500 880.950 996.600 883.050 ;
        RECT 997.800 880.950 999.900 883.050 ;
        RECT 1015.950 880.950 1018.050 883.050 ;
        RECT 1018.950 880.950 1021.050 883.050 ;
        RECT 1021.950 880.950 1024.050 883.050 ;
        RECT 994.200 879.150 996.000 880.950 ;
        RECT 998.400 873.600 999.300 880.950 ;
        RECT 968.100 861.000 969.900 867.000 ;
        RECT 971.100 861.600 972.900 867.600 ;
        RECT 989.100 861.000 990.900 867.600 ;
        RECT 992.100 861.600 993.900 867.600 ;
        RECT 995.100 861.000 996.900 873.000 ;
        RECT 998.100 861.600 999.900 873.600 ;
        RECT 1019.700 867.600 1020.900 880.950 ;
        RECT 1016.100 861.000 1017.900 867.600 ;
        RECT 1019.100 861.600 1020.900 867.600 ;
        RECT 1022.100 861.000 1023.900 867.600 ;
        RECT 17.100 845.400 18.900 857.400 ;
        RECT 20.100 847.200 21.900 858.000 ;
        RECT 23.100 851.400 24.900 857.400 ;
        RECT 26.700 851.400 28.500 858.000 ;
        RECT 29.700 852.300 31.500 857.400 ;
        RECT 29.400 851.400 31.500 852.300 ;
        RECT 32.700 851.400 34.500 858.000 ;
        RECT 17.100 838.050 18.300 845.400 ;
        RECT 23.700 844.500 24.900 851.400 ;
        RECT 29.400 850.500 30.300 851.400 ;
        RECT 19.200 843.600 24.900 844.500 ;
        RECT 26.700 849.600 30.300 850.500 ;
        RECT 19.200 842.700 21.000 843.600 ;
        RECT 17.100 835.950 19.200 838.050 ;
        RECT 17.100 828.600 18.300 835.950 ;
        RECT 20.100 831.300 21.000 842.700 ;
        RECT 22.800 838.050 24.600 839.850 ;
        RECT 22.500 835.950 24.600 838.050 ;
        RECT 19.200 830.400 21.000 831.300 ;
        RECT 26.700 833.400 27.900 849.600 ;
        RECT 31.200 848.400 33.000 848.700 ;
        RECT 35.700 848.400 37.500 857.400 ;
        RECT 38.700 851.400 40.500 858.000 ;
        RECT 42.300 854.400 44.100 857.400 ;
        RECT 45.300 854.400 47.100 857.400 ;
        RECT 42.300 852.300 44.400 854.400 ;
        RECT 45.300 852.300 47.400 854.400 ;
        RECT 48.300 851.400 50.100 857.400 ;
        RECT 51.300 851.400 53.100 858.000 ;
        RECT 47.700 849.300 49.800 851.400 ;
        RECT 55.200 849.900 57.000 857.400 ;
        RECT 58.200 851.400 60.000 858.000 ;
        RECT 61.200 851.400 63.000 857.400 ;
        RECT 64.200 854.400 66.000 857.400 ;
        RECT 67.200 854.400 69.000 857.400 ;
        RECT 70.200 854.400 72.000 857.400 ;
        RECT 64.200 852.300 66.300 854.400 ;
        RECT 67.200 852.300 69.300 854.400 ;
        RECT 70.200 852.300 72.300 854.400 ;
        RECT 73.200 851.400 75.000 858.000 ;
        RECT 76.200 851.400 78.000 857.400 ;
        RECT 79.200 851.400 81.000 858.000 ;
        RECT 82.200 851.400 84.000 857.400 ;
        RECT 85.200 851.400 87.000 858.000 ;
        RECT 88.500 851.400 90.300 857.400 ;
        RECT 91.500 851.400 93.300 858.000 ;
        RECT 31.200 847.200 50.400 848.400 ;
        RECT 55.200 847.800 58.500 849.900 ;
        RECT 61.200 847.500 63.900 851.400 ;
        RECT 67.200 850.500 69.300 851.400 ;
        RECT 67.200 849.300 75.300 850.500 ;
        RECT 73.500 848.700 75.300 849.300 ;
        RECT 76.200 848.400 77.400 851.400 ;
        RECT 82.800 850.500 84.000 851.400 ;
        RECT 82.800 849.600 86.700 850.500 ;
        RECT 80.100 848.400 81.900 849.000 ;
        RECT 31.200 846.900 33.000 847.200 ;
        RECT 49.200 846.600 50.400 847.200 ;
        RECT 64.800 846.600 66.900 847.500 ;
        RECT 34.500 845.700 36.300 846.300 ;
        RECT 44.400 845.700 46.500 846.300 ;
        RECT 34.500 844.500 46.500 845.700 ;
        RECT 49.200 845.400 66.900 846.600 ;
        RECT 70.200 846.300 72.300 847.500 ;
        RECT 76.200 847.200 81.900 848.400 ;
        RECT 85.800 846.300 86.700 849.600 ;
        RECT 70.200 845.400 86.700 846.300 ;
        RECT 44.400 844.200 46.500 844.500 ;
        RECT 49.200 843.300 84.900 844.500 ;
        RECT 49.200 842.700 50.400 843.300 ;
        RECT 83.100 842.700 84.900 843.300 ;
        RECT 36.900 841.800 50.400 842.700 ;
        RECT 61.800 841.800 63.900 842.100 ;
        RECT 36.900 841.050 38.700 841.800 ;
        RECT 28.800 838.950 30.900 841.050 ;
        RECT 34.800 839.250 38.700 841.050 ;
        RECT 56.400 840.300 58.500 841.200 ;
        RECT 34.800 838.950 36.900 839.250 ;
        RECT 47.400 839.100 58.500 840.300 ;
        RECT 60.000 840.000 63.900 841.800 ;
        RECT 68.100 840.300 69.900 842.100 ;
        RECT 69.000 839.100 69.900 840.300 ;
        RECT 29.100 837.300 30.900 838.950 ;
        RECT 47.400 838.500 49.200 839.100 ;
        RECT 56.400 838.200 69.900 839.100 ;
        RECT 72.600 838.800 77.700 840.600 ;
        RECT 79.800 838.950 81.900 841.050 ;
        RECT 72.600 837.300 73.500 838.800 ;
        RECT 29.100 836.100 73.500 837.300 ;
        RECT 79.800 836.100 81.300 838.950 ;
        RECT 44.400 833.400 46.200 835.200 ;
        RECT 52.800 834.000 54.900 835.050 ;
        RECT 74.700 834.600 81.300 836.100 ;
        RECT 26.700 832.200 43.500 833.400 ;
        RECT 19.200 829.500 24.900 830.400 ;
        RECT 17.100 822.600 18.900 828.600 ;
        RECT 20.100 822.000 21.900 828.600 ;
        RECT 23.700 825.600 24.900 829.500 ;
        RECT 23.100 822.600 24.900 825.600 ;
        RECT 26.700 828.600 27.900 832.200 ;
        RECT 41.400 831.300 43.500 832.200 ;
        RECT 30.900 830.700 32.700 831.300 ;
        RECT 30.900 829.500 39.300 830.700 ;
        RECT 37.800 828.600 39.300 829.500 ;
        RECT 44.400 830.400 45.300 833.400 ;
        RECT 49.800 833.100 54.900 834.000 ;
        RECT 49.800 832.200 51.600 833.100 ;
        RECT 52.800 832.950 54.900 833.100 ;
        RECT 59.100 833.100 76.200 834.600 ;
        RECT 59.100 832.500 61.200 833.100 ;
        RECT 59.100 830.700 60.900 832.500 ;
        RECT 77.100 831.900 84.900 833.700 ;
        RECT 44.400 829.200 51.600 830.400 ;
        RECT 46.800 828.600 48.600 829.200 ;
        RECT 50.700 828.600 51.600 829.200 ;
        RECT 66.300 828.600 72.900 830.400 ;
        RECT 77.100 828.600 78.600 831.900 ;
        RECT 85.800 828.600 86.700 845.400 ;
        RECT 26.700 822.600 28.500 828.600 ;
        RECT 32.100 822.000 33.900 828.600 ;
        RECT 37.500 822.600 39.300 828.600 ;
        RECT 41.700 825.600 43.800 827.700 ;
        RECT 44.700 825.600 46.800 827.700 ;
        RECT 47.700 825.600 49.800 827.700 ;
        RECT 50.700 827.400 53.400 828.600 ;
        RECT 51.600 826.500 53.400 827.400 ;
        RECT 55.200 826.500 57.900 828.600 ;
        RECT 41.700 822.600 43.500 825.600 ;
        RECT 44.700 822.600 46.500 825.600 ;
        RECT 47.700 822.600 49.500 825.600 ;
        RECT 50.700 822.000 52.500 825.600 ;
        RECT 55.200 822.600 57.000 826.500 ;
        RECT 61.200 825.600 63.300 827.700 ;
        RECT 64.200 825.600 66.300 827.700 ;
        RECT 67.200 825.600 69.300 827.700 ;
        RECT 70.200 825.600 72.300 827.700 ;
        RECT 74.400 827.400 78.600 828.600 ;
        RECT 58.200 822.000 60.000 825.600 ;
        RECT 61.200 822.600 63.000 825.600 ;
        RECT 64.200 822.600 66.000 825.600 ;
        RECT 67.200 822.600 69.000 825.600 ;
        RECT 70.200 822.600 72.000 825.600 ;
        RECT 74.400 822.600 76.200 827.400 ;
        RECT 79.500 822.000 81.300 828.600 ;
        RECT 84.900 822.600 86.700 828.600 ;
        RECT 88.500 841.050 90.000 851.400 ;
        RECT 111.000 846.600 112.800 857.400 ;
        RECT 111.000 845.400 114.600 846.600 ;
        RECT 116.100 845.400 117.900 858.000 ;
        RECT 134.100 851.400 135.900 858.000 ;
        RECT 137.100 851.400 138.900 857.400 ;
        RECT 88.500 838.950 90.900 841.050 ;
        RECT 88.500 825.600 90.000 838.950 ;
        RECT 110.100 838.050 111.900 839.850 ;
        RECT 113.700 838.050 114.600 845.400 ;
        RECT 115.950 838.050 117.750 839.850 ;
        RECT 134.100 838.050 135.900 839.850 ;
        RECT 137.100 838.050 138.300 851.400 ;
        RECT 156.600 845.400 158.400 858.000 ;
        RECT 161.100 845.400 164.400 857.400 ;
        RECT 167.100 845.400 168.900 858.000 ;
        RECT 186.000 846.600 187.800 857.400 ;
        RECT 186.000 845.400 189.600 846.600 ;
        RECT 191.100 845.400 192.900 858.000 ;
        RECT 209.100 851.400 210.900 857.400 ;
        RECT 212.100 852.000 213.900 858.000 ;
        RECT 210.000 851.100 210.900 851.400 ;
        RECT 215.100 851.400 216.900 857.400 ;
        RECT 218.100 851.400 219.900 858.000 ;
        RECT 236.100 851.400 237.900 858.000 ;
        RECT 239.100 851.400 240.900 857.400 ;
        RECT 257.100 851.400 258.900 857.400 ;
        RECT 260.100 852.000 261.900 858.000 ;
        RECT 215.100 851.100 216.600 851.400 ;
        RECT 210.000 850.200 216.600 851.100 ;
        RECT 155.250 838.050 157.050 839.850 ;
        RECT 162.000 838.050 163.050 845.400 ;
        RECT 167.100 838.050 168.900 839.850 ;
        RECT 185.100 838.050 186.900 839.850 ;
        RECT 188.700 838.050 189.600 845.400 ;
        RECT 190.950 838.050 192.750 839.850 ;
        RECT 210.000 838.050 210.900 850.200 ;
        RECT 215.100 838.050 216.900 839.850 ;
        RECT 236.100 838.050 237.900 839.850 ;
        RECT 239.100 838.050 240.300 851.400 ;
        RECT 258.000 851.100 258.900 851.400 ;
        RECT 263.100 851.400 264.900 857.400 ;
        RECT 266.100 851.400 267.900 858.000 ;
        RECT 284.100 851.400 285.900 857.400 ;
        RECT 287.100 852.000 288.900 858.000 ;
        RECT 263.100 851.100 264.600 851.400 ;
        RECT 258.000 850.200 264.600 851.100 ;
        RECT 285.000 851.100 285.900 851.400 ;
        RECT 290.100 851.400 291.900 857.400 ;
        RECT 293.100 851.400 294.900 858.000 ;
        RECT 311.100 851.400 312.900 858.000 ;
        RECT 314.100 851.400 315.900 857.400 ;
        RECT 317.100 851.400 318.900 858.000 ;
        RECT 335.700 851.400 337.500 858.000 ;
        RECT 290.100 851.100 291.600 851.400 ;
        RECT 285.000 850.200 291.600 851.100 ;
        RECT 258.000 838.050 258.900 850.200 ;
        RECT 263.100 838.050 264.900 839.850 ;
        RECT 285.000 838.050 285.900 850.200 ;
        RECT 286.950 846.450 289.050 847.050 ;
        RECT 310.950 846.450 313.050 847.050 ;
        RECT 286.950 845.550 313.050 846.450 ;
        RECT 286.950 844.950 289.050 845.550 ;
        RECT 310.950 844.950 313.050 845.550 ;
        RECT 290.100 838.050 291.900 839.850 ;
        RECT 314.100 838.050 315.300 851.400 ;
        RECT 336.000 848.100 337.800 849.900 ;
        RECT 316.950 846.450 319.050 847.050 ;
        RECT 338.700 846.900 340.500 857.400 ;
        RECT 334.950 846.450 337.050 846.900 ;
        RECT 316.950 845.550 337.050 846.450 ;
        RECT 316.950 844.950 319.050 845.550 ;
        RECT 334.950 844.800 337.050 845.550 ;
        RECT 338.100 845.400 340.500 846.900 ;
        RECT 343.800 845.400 345.600 858.000 ;
        RECT 363.000 846.600 364.800 857.400 ;
        RECT 363.000 845.400 366.600 846.600 ;
        RECT 368.100 845.400 369.900 858.000 ;
        RECT 386.100 851.400 387.900 857.400 ;
        RECT 389.100 851.400 390.900 858.000 ;
        RECT 316.950 843.450 319.050 843.900 ;
        RECT 328.950 843.450 331.050 844.050 ;
        RECT 316.950 842.550 331.050 843.450 ;
        RECT 316.950 841.800 319.050 842.550 ;
        RECT 328.950 841.950 331.050 842.550 ;
        RECT 338.100 838.050 339.300 845.400 ;
        RECT 344.100 838.050 345.900 839.850 ;
        RECT 362.100 838.050 363.900 839.850 ;
        RECT 365.700 838.050 366.600 845.400 ;
        RECT 367.950 838.050 369.750 839.850 ;
        RECT 386.700 838.050 387.900 851.400 ;
        RECT 407.100 845.400 408.900 857.400 ;
        RECT 410.100 845.400 411.900 858.000 ;
        RECT 428.100 846.300 429.900 857.400 ;
        RECT 431.100 847.200 432.900 858.000 ;
        RECT 434.100 846.300 435.900 857.400 ;
        RECT 428.100 845.400 435.900 846.300 ;
        RECT 437.100 845.400 438.900 857.400 ;
        RECT 455.100 845.400 456.900 858.000 ;
        RECT 460.200 846.600 462.000 857.400 ;
        RECT 458.400 845.400 462.000 846.600 ;
        RECT 479.100 845.400 480.900 858.000 ;
        RECT 483.600 845.400 486.900 857.400 ;
        RECT 489.600 845.400 491.400 858.000 ;
        RECT 510.000 846.600 511.800 857.400 ;
        RECT 510.000 845.400 513.600 846.600 ;
        RECT 515.100 845.400 516.900 858.000 ;
        RECT 533.400 845.400 535.200 858.000 ;
        RECT 538.500 846.900 540.300 857.400 ;
        RECT 541.500 851.400 543.300 858.000 ;
        RECT 560.100 851.400 561.900 858.000 ;
        RECT 563.100 851.400 564.900 857.400 ;
        RECT 566.100 851.400 567.900 858.000 ;
        RECT 541.200 848.100 543.000 849.900 ;
        RECT 538.500 845.400 540.900 846.900 ;
        RECT 389.100 838.050 390.900 839.850 ;
        RECT 407.700 838.050 408.900 845.400 ;
        RECT 409.950 843.450 412.050 844.050 ;
        RECT 418.950 843.450 421.050 844.050 ;
        RECT 409.950 842.550 421.050 843.450 ;
        RECT 409.950 841.950 412.050 842.550 ;
        RECT 418.950 841.950 421.050 842.550 ;
        RECT 431.250 838.050 433.050 839.850 ;
        RECT 437.700 838.050 438.600 845.400 ;
        RECT 455.250 838.050 457.050 839.850 ;
        RECT 458.400 838.050 459.300 845.400 ;
        RECT 463.950 840.450 468.000 841.050 ;
        RECT 461.100 838.050 462.900 839.850 ;
        RECT 463.950 838.950 468.450 840.450 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 112.950 835.950 115.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 157.950 835.950 160.050 838.050 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 113.700 825.600 114.600 835.950 ;
        RECT 127.950 828.450 130.050 829.050 ;
        RECT 133.950 828.450 136.050 829.050 ;
        RECT 127.950 827.550 136.050 828.450 ;
        RECT 127.950 826.950 130.050 827.550 ;
        RECT 133.950 826.950 136.050 827.550 ;
        RECT 137.100 825.600 138.300 835.950 ;
        RECT 158.250 834.150 160.050 835.950 ;
        RECT 162.000 831.300 163.050 835.950 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 166.950 835.950 169.050 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 292.950 835.950 295.050 838.050 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 316.950 835.950 319.050 838.050 ;
        RECT 334.950 835.950 337.050 838.050 ;
        RECT 337.950 835.950 340.050 838.050 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 427.950 835.950 430.050 838.050 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 163.950 834.150 165.750 835.950 ;
        RECT 158.700 830.100 163.050 831.300 ;
        RECT 158.700 828.600 159.600 830.100 ;
        RECT 88.500 822.600 90.300 825.600 ;
        RECT 91.500 822.000 93.300 825.600 ;
        RECT 110.100 822.000 111.900 825.600 ;
        RECT 113.100 822.600 114.900 825.600 ;
        RECT 116.100 822.000 117.900 825.600 ;
        RECT 134.100 822.000 135.900 825.600 ;
        RECT 137.100 822.600 138.900 825.600 ;
        RECT 155.100 823.500 156.900 828.600 ;
        RECT 158.100 824.400 159.900 828.600 ;
        RECT 161.100 828.000 168.900 828.900 ;
        RECT 161.100 823.500 162.900 828.000 ;
        RECT 155.100 822.600 162.900 823.500 ;
        RECT 164.100 822.000 165.900 827.100 ;
        RECT 167.100 822.600 168.900 828.000 ;
        RECT 188.700 825.600 189.600 835.950 ;
        RECT 210.000 832.200 210.900 835.950 ;
        RECT 212.100 834.150 213.900 835.950 ;
        RECT 218.100 834.150 219.900 835.950 ;
        RECT 210.000 831.000 213.300 832.200 ;
        RECT 185.100 822.000 186.900 825.600 ;
        RECT 188.100 822.600 189.900 825.600 ;
        RECT 191.100 822.000 192.900 825.600 ;
        RECT 211.500 822.600 213.300 831.000 ;
        RECT 218.100 822.000 219.900 831.600 ;
        RECT 239.100 825.600 240.300 835.950 ;
        RECT 258.000 832.200 258.900 835.950 ;
        RECT 260.100 834.150 261.900 835.950 ;
        RECT 266.100 834.150 267.900 835.950 ;
        RECT 285.000 832.200 285.900 835.950 ;
        RECT 287.100 834.150 288.900 835.950 ;
        RECT 293.100 834.150 294.900 835.950 ;
        RECT 311.250 834.150 313.050 835.950 ;
        RECT 258.000 831.000 261.300 832.200 ;
        RECT 236.100 822.000 237.900 825.600 ;
        RECT 239.100 822.600 240.900 825.600 ;
        RECT 259.500 822.600 261.300 831.000 ;
        RECT 266.100 822.000 267.900 831.600 ;
        RECT 285.000 831.000 288.300 832.200 ;
        RECT 286.500 822.600 288.300 831.000 ;
        RECT 293.100 822.000 294.900 831.600 ;
        RECT 314.100 830.700 315.300 835.950 ;
        RECT 317.100 834.150 318.900 835.950 ;
        RECT 335.100 834.150 336.900 835.950 ;
        RECT 338.100 831.600 339.300 835.950 ;
        RECT 341.100 834.150 342.900 835.950 ;
        RECT 335.700 830.700 339.300 831.600 ;
        RECT 314.100 829.800 318.300 830.700 ;
        RECT 311.400 822.000 313.200 828.600 ;
        RECT 316.500 822.600 318.300 829.800 ;
        RECT 335.700 828.600 336.900 830.700 ;
        RECT 335.100 822.600 336.900 828.600 ;
        RECT 338.100 827.700 345.900 829.050 ;
        RECT 338.100 822.600 339.900 827.700 ;
        RECT 341.100 822.000 342.900 826.800 ;
        RECT 344.100 822.600 345.900 827.700 ;
        RECT 365.700 825.600 366.600 835.950 ;
        RECT 386.700 825.600 387.900 835.950 ;
        RECT 407.700 828.600 408.900 835.950 ;
        RECT 410.100 834.150 411.900 835.950 ;
        RECT 428.100 834.150 429.900 835.950 ;
        RECT 434.250 834.150 436.050 835.950 ;
        RECT 437.700 828.600 438.600 835.950 ;
        RECT 362.100 822.000 363.900 825.600 ;
        RECT 365.100 822.600 366.900 825.600 ;
        RECT 368.100 822.000 369.900 825.600 ;
        RECT 386.100 822.600 387.900 825.600 ;
        RECT 389.100 822.000 390.900 825.600 ;
        RECT 407.100 822.600 408.900 828.600 ;
        RECT 410.100 822.000 411.900 828.600 ;
        RECT 429.000 822.000 430.800 828.600 ;
        RECT 433.500 827.400 438.600 828.600 ;
        RECT 433.500 822.600 435.300 827.400 ;
        RECT 458.400 825.600 459.300 835.950 ;
        RECT 467.550 835.050 468.450 838.950 ;
        RECT 479.100 838.050 480.900 839.850 ;
        RECT 484.950 838.050 486.000 845.400 ;
        RECT 490.950 838.050 492.750 839.850 ;
        RECT 509.100 838.050 510.900 839.850 ;
        RECT 512.700 838.050 513.600 845.400 ;
        RECT 514.950 838.050 516.750 839.850 ;
        RECT 533.100 838.050 534.900 839.850 ;
        RECT 539.700 838.050 540.900 845.400 ;
        RECT 563.100 838.050 564.300 851.400 ;
        RECT 584.100 845.400 585.900 857.400 ;
        RECT 587.100 846.300 588.900 857.400 ;
        RECT 590.100 847.200 591.900 858.000 ;
        RECT 593.100 846.300 594.900 857.400 ;
        RECT 587.100 845.400 594.900 846.300 ;
        RECT 611.100 845.400 612.900 858.000 ;
        RECT 616.200 846.600 618.000 857.400 ;
        RECT 614.400 845.400 618.000 846.600 ;
        RECT 636.000 846.600 637.800 857.400 ;
        RECT 636.000 845.400 639.600 846.600 ;
        RECT 641.100 845.400 642.900 858.000 ;
        RECT 659.100 851.400 660.900 857.400 ;
        RECT 662.100 852.000 663.900 858.000 ;
        RECT 660.000 851.100 660.900 851.400 ;
        RECT 665.100 851.400 666.900 857.400 ;
        RECT 668.100 851.400 669.900 858.000 ;
        RECT 686.100 851.400 687.900 858.000 ;
        RECT 689.100 851.400 690.900 857.400 ;
        RECT 692.100 851.400 693.900 858.000 ;
        RECT 665.100 851.100 666.600 851.400 ;
        RECT 660.000 850.200 666.600 851.100 ;
        RECT 584.400 838.050 585.300 845.400 ;
        RECT 589.950 838.050 591.750 839.850 ;
        RECT 611.250 838.050 613.050 839.850 ;
        RECT 614.400 838.050 615.300 845.400 ;
        RECT 617.100 838.050 618.900 839.850 ;
        RECT 635.100 838.050 636.900 839.850 ;
        RECT 638.700 838.050 639.600 845.400 ;
        RECT 640.950 838.050 642.750 839.850 ;
        RECT 660.000 838.050 660.900 850.200 ;
        RECT 665.100 838.050 666.900 839.850 ;
        RECT 689.700 838.050 690.900 851.400 ;
        RECT 711.000 846.600 712.800 857.400 ;
        RECT 711.000 845.400 714.600 846.600 ;
        RECT 716.100 845.400 717.900 858.000 ;
        RECT 734.100 847.500 735.900 857.400 ;
        RECT 737.100 848.400 738.900 858.000 ;
        RECT 740.100 856.500 747.900 857.400 ;
        RECT 740.100 847.500 741.900 856.500 ;
        RECT 734.100 846.600 741.900 847.500 ;
        RECT 743.100 847.800 744.900 855.600 ;
        RECT 746.100 848.700 747.900 856.500 ;
        RECT 749.100 856.500 756.900 857.400 ;
        RECT 749.100 847.800 750.900 856.500 ;
        RECT 743.100 846.900 750.900 847.800 ;
        RECT 752.100 847.800 753.900 855.600 ;
        RECT 691.950 843.450 694.050 844.050 ;
        RECT 700.950 843.450 703.050 844.050 ;
        RECT 691.950 842.550 703.050 843.450 ;
        RECT 691.950 841.950 694.050 842.550 ;
        RECT 700.950 841.950 703.050 842.550 ;
        RECT 710.100 838.050 711.900 839.850 ;
        RECT 713.700 838.050 714.600 845.400 ;
        RECT 715.950 843.450 718.050 844.050 ;
        RECT 730.950 843.450 733.050 844.050 ;
        RECT 715.950 842.550 733.050 843.450 ;
        RECT 715.950 841.950 718.050 842.550 ;
        RECT 730.950 841.950 733.050 842.550 ;
        RECT 715.950 838.050 717.750 839.850 ;
        RECT 737.100 838.050 738.900 839.850 ;
        RECT 746.250 838.050 748.050 839.850 ;
        RECT 752.100 838.050 753.300 847.800 ;
        RECT 755.100 847.200 756.900 856.500 ;
        RECT 773.100 846.300 774.900 857.400 ;
        RECT 776.100 847.200 777.900 858.000 ;
        RECT 779.100 846.300 780.900 857.400 ;
        RECT 773.100 845.400 780.900 846.300 ;
        RECT 782.100 845.400 783.900 857.400 ;
        RECT 800.100 851.400 801.900 858.000 ;
        RECT 803.100 851.400 804.900 857.400 ;
        RECT 806.100 852.000 807.900 858.000 ;
        RECT 803.400 851.100 804.900 851.400 ;
        RECT 809.100 851.400 810.900 857.400 ;
        RECT 827.700 851.400 829.500 858.000 ;
        RECT 809.100 851.100 810.000 851.400 ;
        RECT 803.400 850.200 810.000 851.100 ;
        RECT 776.250 838.050 778.050 839.850 ;
        RECT 782.700 838.050 783.600 845.400 ;
        RECT 803.100 838.050 804.900 839.850 ;
        RECT 809.100 838.050 810.000 850.200 ;
        RECT 828.000 848.100 829.800 849.900 ;
        RECT 830.700 846.900 832.500 857.400 ;
        RECT 830.100 845.400 832.500 846.900 ;
        RECT 835.800 845.400 837.600 858.000 ;
        RECT 854.100 845.400 855.900 858.000 ;
        RECT 859.200 846.600 861.000 857.400 ;
        RECT 857.400 845.400 861.000 846.600 ;
        RECT 878.400 845.400 880.200 858.000 ;
        RECT 883.500 846.900 885.300 857.400 ;
        RECT 886.500 851.400 888.300 858.000 ;
        RECT 886.200 848.100 888.000 849.900 ;
        RECT 883.500 845.400 885.900 846.900 ;
        RECT 905.400 845.400 907.200 858.000 ;
        RECT 910.500 846.900 912.300 857.400 ;
        RECT 913.500 851.400 915.300 858.000 ;
        RECT 932.100 851.400 933.900 858.000 ;
        RECT 935.100 851.400 936.900 857.400 ;
        RECT 938.100 851.400 939.900 858.000 ;
        RECT 956.100 851.400 957.900 858.000 ;
        RECT 959.100 851.400 960.900 857.400 ;
        RECT 962.100 852.000 963.900 858.000 ;
        RECT 913.200 848.100 915.000 849.900 ;
        RECT 910.500 845.400 912.900 846.900 ;
        RECT 830.100 838.050 831.300 845.400 ;
        RECT 836.100 838.050 837.900 839.850 ;
        RECT 854.250 838.050 856.050 839.850 ;
        RECT 857.400 838.050 858.300 845.400 ;
        RECT 860.100 838.050 861.900 839.850 ;
        RECT 878.100 838.050 879.900 839.850 ;
        RECT 884.700 838.050 885.900 845.400 ;
        RECT 905.100 838.050 906.900 839.850 ;
        RECT 911.700 838.050 912.900 845.400 ;
        RECT 922.950 843.450 925.050 844.050 ;
        RECT 931.950 843.450 934.050 844.050 ;
        RECT 922.950 842.550 934.050 843.450 ;
        RECT 922.950 841.950 925.050 842.550 ;
        RECT 931.950 841.950 934.050 842.550 ;
        RECT 935.100 838.050 936.300 851.400 ;
        RECT 959.400 851.100 960.900 851.400 ;
        RECT 965.100 851.400 966.900 857.400 ;
        RECT 983.100 851.400 984.900 858.000 ;
        RECT 986.100 851.400 987.900 857.400 ;
        RECT 989.100 851.400 990.900 858.000 ;
        RECT 1007.100 851.400 1008.900 858.000 ;
        RECT 1010.100 851.400 1011.900 857.400 ;
        RECT 1013.100 851.400 1014.900 858.000 ;
        RECT 1031.700 851.400 1033.500 858.000 ;
        RECT 965.100 851.100 966.000 851.400 ;
        RECT 959.400 850.200 966.000 851.100 ;
        RECT 959.100 838.050 960.900 839.850 ;
        RECT 965.100 838.050 966.000 850.200 ;
        RECT 982.950 844.050 985.050 844.200 ;
        RECT 981.000 843.450 985.050 844.050 ;
        RECT 980.550 842.100 985.050 843.450 ;
        RECT 980.550 841.950 984.000 842.100 ;
        RECT 967.950 840.450 972.000 841.050 ;
        RECT 980.550 840.450 981.450 841.950 ;
        RECT 967.950 838.950 972.450 840.450 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 463.950 833.550 468.450 835.050 ;
        RECT 482.250 834.150 484.050 835.950 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 487.950 835.950 490.050 838.050 ;
        RECT 490.950 835.950 493.050 838.050 ;
        RECT 508.950 835.950 511.050 838.050 ;
        RECT 511.950 835.950 514.050 838.050 ;
        RECT 514.950 835.950 517.050 838.050 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 592.950 835.950 595.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 661.950 835.950 664.050 838.050 ;
        RECT 664.950 835.950 667.050 838.050 ;
        RECT 667.950 835.950 670.050 838.050 ;
        RECT 685.950 835.950 688.050 838.050 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 736.800 835.950 738.900 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 751.500 835.950 753.600 838.050 ;
        RECT 772.950 835.950 775.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 805.950 835.950 808.050 838.050 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 829.950 835.950 832.050 838.050 ;
        RECT 832.950 835.950 835.050 838.050 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 907.950 835.950 910.050 838.050 ;
        RECT 910.950 835.950 913.050 838.050 ;
        RECT 913.950 835.950 916.050 838.050 ;
        RECT 931.950 835.950 934.050 838.050 ;
        RECT 934.950 835.950 937.050 838.050 ;
        RECT 937.950 835.950 940.050 838.050 ;
        RECT 955.950 835.950 958.050 838.050 ;
        RECT 958.950 835.950 961.050 838.050 ;
        RECT 961.950 835.950 964.050 838.050 ;
        RECT 964.950 835.950 967.050 838.050 ;
        RECT 463.950 832.950 468.000 833.550 ;
        RECT 484.950 831.300 486.000 835.950 ;
        RECT 487.950 834.150 489.750 835.950 ;
        RECT 484.950 830.100 489.300 831.300 ;
        RECT 479.100 828.000 486.900 828.900 ;
        RECT 488.400 828.600 489.300 830.100 ;
        RECT 436.500 822.000 438.300 825.600 ;
        RECT 455.100 822.000 456.900 825.600 ;
        RECT 458.100 822.600 459.900 825.600 ;
        RECT 461.100 822.000 462.900 825.600 ;
        RECT 479.100 822.600 480.900 828.000 ;
        RECT 482.100 822.000 483.900 827.100 ;
        RECT 485.100 823.500 486.900 828.000 ;
        RECT 488.100 824.400 489.900 828.600 ;
        RECT 491.100 823.500 492.900 828.600 ;
        RECT 512.700 825.600 513.600 835.950 ;
        RECT 536.100 834.150 537.900 835.950 ;
        RECT 539.700 831.600 540.900 835.950 ;
        RECT 542.100 834.150 543.900 835.950 ;
        RECT 560.250 834.150 562.050 835.950 ;
        RECT 539.700 830.700 543.300 831.600 ;
        RECT 533.100 827.700 540.900 829.050 ;
        RECT 485.100 822.600 492.900 823.500 ;
        RECT 509.100 822.000 510.900 825.600 ;
        RECT 512.100 822.600 513.900 825.600 ;
        RECT 515.100 822.000 516.900 825.600 ;
        RECT 533.100 822.600 534.900 827.700 ;
        RECT 536.100 822.000 537.900 826.800 ;
        RECT 539.100 822.600 540.900 827.700 ;
        RECT 542.100 828.600 543.300 830.700 ;
        RECT 563.100 830.700 564.300 835.950 ;
        RECT 566.100 834.150 567.900 835.950 ;
        RECT 563.100 829.800 567.300 830.700 ;
        RECT 542.100 822.600 543.900 828.600 ;
        RECT 560.400 822.000 562.200 828.600 ;
        RECT 565.500 822.600 567.300 829.800 ;
        RECT 584.400 828.600 585.300 835.950 ;
        RECT 586.950 834.150 588.750 835.950 ;
        RECT 593.100 834.150 594.900 835.950 ;
        RECT 589.950 831.450 592.050 832.050 ;
        RECT 601.950 831.450 604.050 832.050 ;
        RECT 589.950 830.550 604.050 831.450 ;
        RECT 589.950 829.950 592.050 830.550 ;
        RECT 601.950 829.950 604.050 830.550 ;
        RECT 584.400 827.400 589.500 828.600 ;
        RECT 584.700 822.000 586.500 825.600 ;
        RECT 587.700 822.600 589.500 827.400 ;
        RECT 592.200 822.000 594.000 828.600 ;
        RECT 614.400 825.600 615.300 835.950 ;
        RECT 616.950 831.450 619.050 832.050 ;
        RECT 625.950 831.450 628.050 832.050 ;
        RECT 616.950 830.550 628.050 831.450 ;
        RECT 616.950 829.950 619.050 830.550 ;
        RECT 625.950 829.950 628.050 830.550 ;
        RECT 638.700 825.600 639.600 835.950 ;
        RECT 660.000 832.200 660.900 835.950 ;
        RECT 662.100 834.150 663.900 835.950 ;
        RECT 668.100 834.150 669.900 835.950 ;
        RECT 686.100 834.150 687.900 835.950 ;
        RECT 660.000 831.000 663.300 832.200 ;
        RECT 611.100 822.000 612.900 825.600 ;
        RECT 614.100 822.600 615.900 825.600 ;
        RECT 617.100 822.000 618.900 825.600 ;
        RECT 635.100 822.000 636.900 825.600 ;
        RECT 638.100 822.600 639.900 825.600 ;
        RECT 641.100 822.000 642.900 825.600 ;
        RECT 661.500 822.600 663.300 831.000 ;
        RECT 668.100 822.000 669.900 831.600 ;
        RECT 689.700 830.700 690.900 835.950 ;
        RECT 691.950 834.150 693.750 835.950 ;
        RECT 686.700 829.800 690.900 830.700 ;
        RECT 686.700 822.600 688.500 829.800 ;
        RECT 691.800 822.000 693.600 828.600 ;
        RECT 713.700 825.600 714.600 835.950 ;
        RECT 724.950 834.450 727.050 835.050 ;
        RECT 733.950 834.450 736.050 835.050 ;
        RECT 724.950 833.550 736.050 834.450 ;
        RECT 742.950 834.150 744.750 835.950 ;
        RECT 724.950 832.950 727.050 833.550 ;
        RECT 733.950 832.950 736.050 833.550 ;
        RECT 724.950 831.450 727.050 831.900 ;
        RECT 748.950 831.450 751.050 832.050 ;
        RECT 724.950 830.550 751.050 831.450 ;
        RECT 724.950 829.800 727.050 830.550 ;
        RECT 748.950 829.950 751.050 830.550 ;
        RECT 752.100 827.400 753.300 835.950 ;
        RECT 773.100 834.150 774.900 835.950 ;
        RECT 779.250 834.150 781.050 835.950 ;
        RECT 782.700 828.600 783.600 835.950 ;
        RECT 800.100 834.150 801.900 835.950 ;
        RECT 806.100 834.150 807.900 835.950 ;
        RECT 809.100 832.200 810.000 835.950 ;
        RECT 827.100 834.150 828.900 835.950 ;
        RECT 740.700 826.500 753.300 827.400 ;
        RECT 740.700 825.600 741.600 826.500 ;
        RECT 747.900 825.600 748.800 826.500 ;
        RECT 710.100 822.000 711.900 825.600 ;
        RECT 713.100 822.600 714.900 825.600 ;
        RECT 716.100 822.000 717.900 825.600 ;
        RECT 736.800 822.000 738.900 825.600 ;
        RECT 740.100 822.600 741.900 825.600 ;
        RECT 743.100 822.000 744.900 825.600 ;
        RECT 746.100 822.600 748.800 825.600 ;
        RECT 774.000 822.000 775.800 828.600 ;
        RECT 778.500 827.400 783.600 828.600 ;
        RECT 778.500 822.600 780.300 827.400 ;
        RECT 781.500 822.000 783.300 825.600 ;
        RECT 800.100 822.000 801.900 831.600 ;
        RECT 806.700 831.000 810.000 832.200 ;
        RECT 830.100 831.600 831.300 835.950 ;
        RECT 833.100 834.150 834.900 835.950 ;
        RECT 844.950 834.450 847.050 835.050 ;
        RECT 850.950 834.450 853.050 835.050 ;
        RECT 844.950 833.550 853.050 834.450 ;
        RECT 844.950 832.950 847.050 833.550 ;
        RECT 850.950 832.950 853.050 833.550 ;
        RECT 806.700 822.600 808.500 831.000 ;
        RECT 827.700 830.700 831.300 831.600 ;
        RECT 827.700 828.600 828.900 830.700 ;
        RECT 827.100 822.600 828.900 828.600 ;
        RECT 830.100 827.700 837.900 829.050 ;
        RECT 830.100 822.600 831.900 827.700 ;
        RECT 833.100 822.000 834.900 826.800 ;
        RECT 836.100 822.600 837.900 827.700 ;
        RECT 857.400 825.600 858.300 835.950 ;
        RECT 862.950 834.450 865.050 835.050 ;
        RECT 868.950 834.450 871.050 835.050 ;
        RECT 862.950 833.550 871.050 834.450 ;
        RECT 881.100 834.150 882.900 835.950 ;
        RECT 862.950 832.950 865.050 833.550 ;
        RECT 868.950 832.950 871.050 833.550 ;
        RECT 884.700 831.600 885.900 835.950 ;
        RECT 887.100 834.150 888.900 835.950 ;
        RECT 908.100 834.150 909.900 835.950 ;
        RECT 911.700 831.600 912.900 835.950 ;
        RECT 914.100 834.150 915.900 835.950 ;
        RECT 932.250 834.150 934.050 835.950 ;
        RECT 884.700 830.700 888.300 831.600 ;
        RECT 911.700 830.700 915.300 831.600 ;
        RECT 878.100 827.700 885.900 829.050 ;
        RECT 854.100 822.000 855.900 825.600 ;
        RECT 857.100 822.600 858.900 825.600 ;
        RECT 860.100 822.000 861.900 825.600 ;
        RECT 878.100 822.600 879.900 827.700 ;
        RECT 881.100 822.000 882.900 826.800 ;
        RECT 884.100 822.600 885.900 827.700 ;
        RECT 887.100 828.600 888.300 830.700 ;
        RECT 887.100 822.600 888.900 828.600 ;
        RECT 905.100 827.700 912.900 829.050 ;
        RECT 905.100 822.600 906.900 827.700 ;
        RECT 908.100 822.000 909.900 826.800 ;
        RECT 911.100 822.600 912.900 827.700 ;
        RECT 914.100 828.600 915.300 830.700 ;
        RECT 935.100 830.700 936.300 835.950 ;
        RECT 938.100 834.150 939.900 835.950 ;
        RECT 956.100 834.150 957.900 835.950 ;
        RECT 962.100 834.150 963.900 835.950 ;
        RECT 965.100 832.200 966.000 835.950 ;
        RECT 971.550 835.050 972.450 838.950 ;
        RECT 967.950 833.550 972.450 835.050 ;
        RECT 977.550 839.550 981.450 840.450 ;
        RECT 977.550 835.050 978.450 839.550 ;
        RECT 986.100 838.050 987.300 851.400 ;
        RECT 1010.700 838.050 1011.900 851.400 ;
        RECT 1032.000 848.100 1033.800 849.900 ;
        RECT 1034.700 846.900 1036.500 857.400 ;
        RECT 1034.100 845.400 1036.500 846.900 ;
        RECT 1039.800 845.400 1041.600 858.000 ;
        RECT 1034.100 838.050 1035.300 845.400 ;
        RECT 1040.100 838.050 1041.900 839.850 ;
        RECT 982.950 835.950 985.050 838.050 ;
        RECT 985.950 835.950 988.050 838.050 ;
        RECT 988.950 835.950 991.050 838.050 ;
        RECT 1006.950 835.950 1009.050 838.050 ;
        RECT 1009.950 835.950 1012.050 838.050 ;
        RECT 1012.950 835.950 1015.050 838.050 ;
        RECT 1030.950 835.950 1033.050 838.050 ;
        RECT 1033.950 835.950 1036.050 838.050 ;
        RECT 1036.950 835.950 1039.050 838.050 ;
        RECT 1039.950 835.950 1042.050 838.050 ;
        RECT 977.550 833.550 982.050 835.050 ;
        RECT 983.250 834.150 985.050 835.950 ;
        RECT 967.950 832.950 972.000 833.550 ;
        RECT 978.000 832.950 982.050 833.550 ;
        RECT 935.100 829.800 939.300 830.700 ;
        RECT 914.100 822.600 915.900 828.600 ;
        RECT 932.400 822.000 934.200 828.600 ;
        RECT 937.500 822.600 939.300 829.800 ;
        RECT 956.100 822.000 957.900 831.600 ;
        RECT 962.700 831.000 966.000 832.200 ;
        RECT 962.700 822.600 964.500 831.000 ;
        RECT 986.100 830.700 987.300 835.950 ;
        RECT 989.100 834.150 990.900 835.950 ;
        RECT 1007.100 834.150 1008.900 835.950 ;
        RECT 1010.700 830.700 1011.900 835.950 ;
        RECT 1012.950 834.150 1014.750 835.950 ;
        RECT 1031.100 834.150 1032.900 835.950 ;
        RECT 1034.100 831.600 1035.300 835.950 ;
        RECT 1037.100 834.150 1038.900 835.950 ;
        RECT 986.100 829.800 990.300 830.700 ;
        RECT 983.400 822.000 985.200 828.600 ;
        RECT 988.500 822.600 990.300 829.800 ;
        RECT 1007.700 829.800 1011.900 830.700 ;
        RECT 1031.700 830.700 1035.300 831.600 ;
        RECT 1007.700 822.600 1009.500 829.800 ;
        RECT 1031.700 828.600 1032.900 830.700 ;
        RECT 1012.800 822.000 1014.600 828.600 ;
        RECT 1031.100 822.600 1032.900 828.600 ;
        RECT 1034.100 827.700 1041.900 829.050 ;
        RECT 1034.100 822.600 1035.900 827.700 ;
        RECT 1037.100 822.000 1038.900 826.800 ;
        RECT 1040.100 822.600 1041.900 827.700 ;
        RECT 2.700 812.400 4.500 818.400 ;
        RECT 8.100 812.400 9.900 819.000 ;
        RECT 13.500 812.400 15.300 818.400 ;
        RECT 17.700 815.400 19.500 818.400 ;
        RECT 20.700 815.400 22.500 818.400 ;
        RECT 23.700 815.400 25.500 818.400 ;
        RECT 26.700 815.400 28.500 819.000 ;
        RECT 17.700 813.300 19.800 815.400 ;
        RECT 20.700 813.300 22.800 815.400 ;
        RECT 23.700 813.300 25.800 815.400 ;
        RECT 31.200 814.500 33.000 818.400 ;
        RECT 34.200 815.400 36.000 819.000 ;
        RECT 37.200 815.400 39.000 818.400 ;
        RECT 40.200 815.400 42.000 818.400 ;
        RECT 43.200 815.400 45.000 818.400 ;
        RECT 46.200 815.400 48.000 818.400 ;
        RECT 27.600 813.600 29.400 814.500 ;
        RECT 26.700 812.400 29.400 813.600 ;
        RECT 31.200 812.400 33.900 814.500 ;
        RECT 37.200 813.300 39.300 815.400 ;
        RECT 40.200 813.300 42.300 815.400 ;
        RECT 43.200 813.300 45.300 815.400 ;
        RECT 46.200 813.300 48.300 815.400 ;
        RECT 50.400 813.600 52.200 818.400 ;
        RECT 50.400 812.400 54.600 813.600 ;
        RECT 55.500 812.400 57.300 819.000 ;
        RECT 60.900 812.400 62.700 818.400 ;
        RECT 2.700 808.800 3.900 812.400 ;
        RECT 13.800 811.500 15.300 812.400 ;
        RECT 22.800 811.800 24.600 812.400 ;
        RECT 26.700 811.800 27.600 812.400 ;
        RECT 6.900 810.300 15.300 811.500 ;
        RECT 20.400 810.600 27.600 811.800 ;
        RECT 42.300 810.600 48.900 812.400 ;
        RECT 6.900 809.700 8.700 810.300 ;
        RECT 17.400 808.800 19.500 809.700 ;
        RECT 2.700 807.600 19.500 808.800 ;
        RECT 20.400 807.600 21.300 810.600 ;
        RECT 25.800 807.900 27.600 808.800 ;
        RECT 35.100 808.500 36.900 810.300 ;
        RECT 53.100 809.100 54.600 812.400 ;
        RECT 28.800 807.900 30.900 808.050 ;
        RECT 2.700 791.400 3.900 807.600 ;
        RECT 20.400 805.800 22.200 807.600 ;
        RECT 25.800 807.000 30.900 807.900 ;
        RECT 28.800 805.950 30.900 807.000 ;
        RECT 35.100 807.900 37.200 808.500 ;
        RECT 35.100 806.400 52.200 807.900 ;
        RECT 53.100 807.300 60.900 809.100 ;
        RECT 50.700 804.900 57.300 806.400 ;
        RECT 5.100 803.700 49.500 804.900 ;
        RECT 5.100 802.050 6.900 803.700 ;
        RECT 4.800 799.950 6.900 802.050 ;
        RECT 10.800 801.750 12.900 802.050 ;
        RECT 23.400 801.900 25.200 802.500 ;
        RECT 32.400 801.900 45.900 802.800 ;
        RECT 10.800 799.950 14.700 801.750 ;
        RECT 23.400 800.700 34.500 801.900 ;
        RECT 12.900 799.200 14.700 799.950 ;
        RECT 32.400 799.800 34.500 800.700 ;
        RECT 36.000 799.200 39.900 801.000 ;
        RECT 45.000 800.700 45.900 801.900 ;
        RECT 12.900 798.300 26.400 799.200 ;
        RECT 37.800 798.900 39.900 799.200 ;
        RECT 44.100 798.900 45.900 800.700 ;
        RECT 48.600 802.200 49.500 803.700 ;
        RECT 48.600 800.400 53.700 802.200 ;
        RECT 55.800 802.050 57.300 804.900 ;
        RECT 55.800 799.950 57.900 802.050 ;
        RECT 25.200 797.700 26.400 798.300 ;
        RECT 59.100 797.700 60.900 798.300 ;
        RECT 20.400 796.500 22.500 796.800 ;
        RECT 25.200 796.500 60.900 797.700 ;
        RECT 10.500 795.300 22.500 796.500 ;
        RECT 61.800 795.600 62.700 812.400 ;
        RECT 10.500 794.700 12.300 795.300 ;
        RECT 20.400 794.700 22.500 795.300 ;
        RECT 25.200 794.400 42.900 795.600 ;
        RECT 7.200 793.800 9.000 794.100 ;
        RECT 25.200 793.800 26.400 794.400 ;
        RECT 7.200 792.600 26.400 793.800 ;
        RECT 40.800 793.500 42.900 794.400 ;
        RECT 46.200 794.700 62.700 795.600 ;
        RECT 46.200 793.500 48.300 794.700 ;
        RECT 7.200 792.300 9.000 792.600 ;
        RECT 2.700 790.500 6.300 791.400 ;
        RECT 5.400 789.600 6.300 790.500 ;
        RECT 2.700 783.000 4.500 789.600 ;
        RECT 5.400 788.700 7.500 789.600 ;
        RECT 5.700 783.600 7.500 788.700 ;
        RECT 8.700 783.000 10.500 789.600 ;
        RECT 11.700 783.600 13.500 792.600 ;
        RECT 23.700 789.600 25.800 791.700 ;
        RECT 31.200 791.100 34.500 793.200 ;
        RECT 14.700 783.000 16.500 789.600 ;
        RECT 18.300 786.600 20.400 788.700 ;
        RECT 21.300 786.600 23.400 788.700 ;
        RECT 18.300 783.600 20.100 786.600 ;
        RECT 21.300 783.600 23.100 786.600 ;
        RECT 24.300 783.600 26.100 789.600 ;
        RECT 27.300 783.000 29.100 789.600 ;
        RECT 31.200 783.600 33.000 791.100 ;
        RECT 37.200 789.600 39.900 793.500 ;
        RECT 52.200 792.600 57.900 793.800 ;
        RECT 49.500 791.700 51.300 792.300 ;
        RECT 43.200 790.500 51.300 791.700 ;
        RECT 43.200 789.600 45.300 790.500 ;
        RECT 52.200 789.600 53.400 792.600 ;
        RECT 56.100 792.000 57.900 792.600 ;
        RECT 61.800 791.400 62.700 794.700 ;
        RECT 58.800 790.500 62.700 791.400 ;
        RECT 64.500 815.400 66.300 818.400 ;
        RECT 67.500 815.400 69.300 819.000 ;
        RECT 64.500 802.050 66.000 815.400 ;
        RECT 86.100 812.400 87.900 818.400 ;
        RECT 86.700 810.300 87.900 812.400 ;
        RECT 89.100 813.300 90.900 818.400 ;
        RECT 92.100 814.200 93.900 819.000 ;
        RECT 95.100 813.300 96.900 818.400 ;
        RECT 89.100 811.950 96.900 813.300 ;
        RECT 86.700 809.400 90.300 810.300 ;
        RECT 115.500 810.000 117.300 818.400 ;
        RECT 86.100 805.050 87.900 806.850 ;
        RECT 89.100 805.050 90.300 809.400 ;
        RECT 114.000 808.800 117.300 810.000 ;
        RECT 122.100 809.400 123.900 819.000 ;
        RECT 137.400 812.400 139.200 819.000 ;
        RECT 142.500 811.200 144.300 818.400 ;
        RECT 140.100 810.300 144.300 811.200 ;
        RECT 146.700 812.400 148.500 818.400 ;
        RECT 152.100 812.400 153.900 819.000 ;
        RECT 157.500 812.400 159.300 818.400 ;
        RECT 161.700 815.400 163.500 818.400 ;
        RECT 164.700 815.400 166.500 818.400 ;
        RECT 167.700 815.400 169.500 818.400 ;
        RECT 170.700 815.400 172.500 819.000 ;
        RECT 161.700 813.300 163.800 815.400 ;
        RECT 164.700 813.300 166.800 815.400 ;
        RECT 167.700 813.300 169.800 815.400 ;
        RECT 175.200 814.500 177.000 818.400 ;
        RECT 178.200 815.400 180.000 819.000 ;
        RECT 181.200 815.400 183.000 818.400 ;
        RECT 184.200 815.400 186.000 818.400 ;
        RECT 187.200 815.400 189.000 818.400 ;
        RECT 190.200 815.400 192.000 818.400 ;
        RECT 171.600 813.600 173.400 814.500 ;
        RECT 170.700 812.400 173.400 813.600 ;
        RECT 175.200 812.400 177.900 814.500 ;
        RECT 181.200 813.300 183.300 815.400 ;
        RECT 184.200 813.300 186.300 815.400 ;
        RECT 187.200 813.300 189.300 815.400 ;
        RECT 190.200 813.300 192.300 815.400 ;
        RECT 194.400 813.600 196.200 818.400 ;
        RECT 194.400 812.400 198.600 813.600 ;
        RECT 199.500 812.400 201.300 819.000 ;
        RECT 204.900 812.400 206.700 818.400 ;
        RECT 97.950 807.450 102.000 808.050 ;
        RECT 92.100 805.050 93.900 806.850 ;
        RECT 97.950 805.950 102.450 807.450 ;
        RECT 85.950 802.950 88.050 805.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 64.500 799.950 66.900 802.050 ;
        RECT 58.800 789.600 60.000 790.500 ;
        RECT 64.500 789.600 66.000 799.950 ;
        RECT 89.100 795.600 90.300 802.950 ;
        RECT 95.100 801.150 96.900 802.950 ;
        RECT 101.550 801.450 102.450 805.950 ;
        RECT 114.000 805.050 114.900 808.800 ;
        RECT 116.100 805.050 117.900 806.850 ;
        RECT 122.100 805.050 123.900 806.850 ;
        RECT 137.250 805.050 139.050 806.850 ;
        RECT 140.100 805.050 141.300 810.300 ;
        RECT 146.700 808.800 147.900 812.400 ;
        RECT 157.800 811.500 159.300 812.400 ;
        RECT 166.800 811.800 168.600 812.400 ;
        RECT 170.700 811.800 171.600 812.400 ;
        RECT 150.900 810.300 159.300 811.500 ;
        RECT 164.400 810.600 171.600 811.800 ;
        RECT 186.300 810.600 192.900 812.400 ;
        RECT 150.900 809.700 152.700 810.300 ;
        RECT 161.400 808.800 163.500 809.700 ;
        RECT 146.700 807.600 163.500 808.800 ;
        RECT 164.400 807.600 165.300 810.600 ;
        RECT 169.800 807.900 171.600 808.800 ;
        RECT 179.100 808.500 180.900 810.300 ;
        RECT 197.100 809.100 198.600 812.400 ;
        RECT 172.800 807.900 174.900 808.050 ;
        RECT 143.100 805.050 144.900 806.850 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 142.950 802.950 145.050 805.050 ;
        RECT 109.950 801.450 112.050 802.050 ;
        RECT 101.550 800.550 112.050 801.450 ;
        RECT 109.950 799.950 112.050 800.550 ;
        RECT 89.100 794.100 91.500 795.600 ;
        RECT 87.000 791.100 88.800 792.900 ;
        RECT 34.200 783.000 36.000 789.600 ;
        RECT 37.200 783.600 39.000 789.600 ;
        RECT 40.200 786.600 42.300 788.700 ;
        RECT 43.200 786.600 45.300 788.700 ;
        RECT 46.200 786.600 48.300 788.700 ;
        RECT 40.200 783.600 42.000 786.600 ;
        RECT 43.200 783.600 45.000 786.600 ;
        RECT 46.200 783.600 48.000 786.600 ;
        RECT 49.200 783.000 51.000 789.600 ;
        RECT 52.200 783.600 54.000 789.600 ;
        RECT 55.200 783.000 57.000 789.600 ;
        RECT 58.200 783.600 60.000 789.600 ;
        RECT 61.200 783.000 63.000 789.600 ;
        RECT 64.500 783.600 66.300 789.600 ;
        RECT 67.500 783.000 69.300 789.600 ;
        RECT 86.700 783.000 88.500 789.600 ;
        RECT 89.700 783.600 91.500 794.100 ;
        RECT 94.800 783.000 96.600 795.600 ;
        RECT 114.000 790.800 114.900 802.950 ;
        RECT 119.100 801.150 120.900 802.950 ;
        RECT 114.000 789.900 120.600 790.800 ;
        RECT 114.000 789.600 114.900 789.900 ;
        RECT 113.100 783.600 114.900 789.600 ;
        RECT 119.100 789.600 120.600 789.900 ;
        RECT 140.100 789.600 141.300 802.950 ;
        RECT 146.700 791.400 147.900 807.600 ;
        RECT 164.400 805.800 166.200 807.600 ;
        RECT 169.800 807.000 174.900 807.900 ;
        RECT 172.800 805.950 174.900 807.000 ;
        RECT 179.100 807.900 181.200 808.500 ;
        RECT 179.100 806.400 196.200 807.900 ;
        RECT 197.100 807.300 204.900 809.100 ;
        RECT 194.700 804.900 201.300 806.400 ;
        RECT 149.100 803.700 193.500 804.900 ;
        RECT 149.100 802.050 150.900 803.700 ;
        RECT 148.800 799.950 150.900 802.050 ;
        RECT 154.800 801.750 156.900 802.050 ;
        RECT 167.400 801.900 169.200 802.500 ;
        RECT 176.400 801.900 189.900 802.800 ;
        RECT 154.800 799.950 158.700 801.750 ;
        RECT 167.400 800.700 178.500 801.900 ;
        RECT 156.900 799.200 158.700 799.950 ;
        RECT 176.400 799.800 178.500 800.700 ;
        RECT 180.000 799.200 183.900 801.000 ;
        RECT 189.000 800.700 189.900 801.900 ;
        RECT 156.900 798.300 170.400 799.200 ;
        RECT 181.800 798.900 183.900 799.200 ;
        RECT 188.100 798.900 189.900 800.700 ;
        RECT 192.600 802.200 193.500 803.700 ;
        RECT 192.600 800.400 197.700 802.200 ;
        RECT 199.800 802.050 201.300 804.900 ;
        RECT 199.800 799.950 201.900 802.050 ;
        RECT 169.200 797.700 170.400 798.300 ;
        RECT 203.100 797.700 204.900 798.300 ;
        RECT 164.400 796.500 166.500 796.800 ;
        RECT 169.200 796.500 204.900 797.700 ;
        RECT 154.500 795.300 166.500 796.500 ;
        RECT 205.800 795.600 206.700 812.400 ;
        RECT 154.500 794.700 156.300 795.300 ;
        RECT 164.400 794.700 166.500 795.300 ;
        RECT 169.200 794.400 186.900 795.600 ;
        RECT 151.200 793.800 153.000 794.100 ;
        RECT 169.200 793.800 170.400 794.400 ;
        RECT 151.200 792.600 170.400 793.800 ;
        RECT 184.800 793.500 186.900 794.400 ;
        RECT 190.200 794.700 206.700 795.600 ;
        RECT 190.200 793.500 192.300 794.700 ;
        RECT 151.200 792.300 153.000 792.600 ;
        RECT 146.700 790.500 150.300 791.400 ;
        RECT 149.400 789.600 150.300 790.500 ;
        RECT 116.100 783.000 117.900 789.000 ;
        RECT 119.100 783.600 120.900 789.600 ;
        RECT 122.100 783.000 123.900 789.600 ;
        RECT 137.100 783.000 138.900 789.600 ;
        RECT 140.100 783.600 141.900 789.600 ;
        RECT 143.100 783.000 144.900 789.600 ;
        RECT 146.700 783.000 148.500 789.600 ;
        RECT 149.400 788.700 151.500 789.600 ;
        RECT 149.700 783.600 151.500 788.700 ;
        RECT 152.700 783.000 154.500 789.600 ;
        RECT 155.700 783.600 157.500 792.600 ;
        RECT 167.700 789.600 169.800 791.700 ;
        RECT 175.200 791.100 178.500 793.200 ;
        RECT 158.700 783.000 160.500 789.600 ;
        RECT 162.300 786.600 164.400 788.700 ;
        RECT 165.300 786.600 167.400 788.700 ;
        RECT 162.300 783.600 164.100 786.600 ;
        RECT 165.300 783.600 167.100 786.600 ;
        RECT 168.300 783.600 170.100 789.600 ;
        RECT 171.300 783.000 173.100 789.600 ;
        RECT 175.200 783.600 177.000 791.100 ;
        RECT 181.200 789.600 183.900 793.500 ;
        RECT 196.200 792.600 201.900 793.800 ;
        RECT 193.500 791.700 195.300 792.300 ;
        RECT 187.200 790.500 195.300 791.700 ;
        RECT 187.200 789.600 189.300 790.500 ;
        RECT 196.200 789.600 197.400 792.600 ;
        RECT 200.100 792.000 201.900 792.600 ;
        RECT 205.800 791.400 206.700 794.700 ;
        RECT 202.800 790.500 206.700 791.400 ;
        RECT 208.500 815.400 210.300 818.400 ;
        RECT 211.500 815.400 213.300 819.000 ;
        RECT 208.500 802.050 210.000 815.400 ;
        RECT 232.500 810.000 234.300 818.400 ;
        RECT 231.000 808.800 234.300 810.000 ;
        RECT 239.100 809.400 240.900 819.000 ;
        RECT 257.100 815.400 258.900 818.400 ;
        RECT 260.100 815.400 261.900 819.000 ;
        RECT 231.000 805.050 231.900 808.800 ;
        RECT 233.100 805.050 234.900 806.850 ;
        RECT 239.100 805.050 240.900 806.850 ;
        RECT 257.700 805.050 258.900 815.400 ;
        RECT 278.700 811.200 280.500 818.400 ;
        RECT 283.800 812.400 285.600 819.000 ;
        RECT 302.100 813.300 303.900 818.400 ;
        RECT 305.100 814.200 306.900 819.000 ;
        RECT 308.100 813.300 309.900 818.400 ;
        RECT 302.100 811.950 309.900 813.300 ;
        RECT 311.100 812.400 312.900 818.400 ;
        RECT 329.100 815.400 330.900 819.000 ;
        RECT 332.100 815.400 333.900 818.400 ;
        RECT 335.100 815.400 336.900 819.000 ;
        RECT 278.700 810.300 282.900 811.200 ;
        RECT 311.100 810.300 312.300 812.400 ;
        RECT 278.100 805.050 279.900 806.850 ;
        RECT 281.700 805.050 282.900 810.300 ;
        RECT 308.700 809.400 312.300 810.300 ;
        RECT 283.950 805.050 285.750 806.850 ;
        RECT 305.100 805.050 306.900 806.850 ;
        RECT 308.700 805.050 309.900 809.400 ;
        RECT 311.100 805.050 312.900 806.850 ;
        RECT 332.400 805.050 333.300 815.400 ;
        RECT 353.100 809.400 354.900 819.000 ;
        RECT 359.700 810.000 361.500 818.400 ;
        RECT 359.700 808.800 363.000 810.000 ;
        RECT 380.100 809.400 381.900 819.000 ;
        RECT 386.700 810.000 388.500 818.400 ;
        RECT 391.950 813.450 394.050 814.050 ;
        RECT 397.950 813.450 400.050 814.050 ;
        RECT 391.950 812.550 400.050 813.450 ;
        RECT 391.950 811.950 394.050 812.550 ;
        RECT 397.950 811.950 400.050 812.550 ;
        RECT 407.100 812.400 408.900 818.400 ;
        RECT 407.700 810.300 408.900 812.400 ;
        RECT 410.100 813.300 411.900 818.400 ;
        RECT 413.100 814.200 414.900 819.000 ;
        RECT 416.100 813.300 417.900 818.400 ;
        RECT 434.100 815.400 435.900 819.000 ;
        RECT 437.100 815.400 438.900 818.400 ;
        RECT 440.100 815.400 441.900 819.000 ;
        RECT 410.100 811.950 417.900 813.300 ;
        RECT 386.700 808.800 390.000 810.000 ;
        RECT 407.700 809.400 411.300 810.300 ;
        RECT 353.100 805.050 354.900 806.850 ;
        RECT 359.100 805.050 360.900 806.850 ;
        RECT 362.100 805.050 363.000 808.800 ;
        RECT 380.100 805.050 381.900 806.850 ;
        RECT 386.100 805.050 387.900 806.850 ;
        RECT 389.100 805.050 390.000 808.800 ;
        RECT 407.100 805.050 408.900 806.850 ;
        RECT 410.100 805.050 411.300 809.400 ;
        RECT 413.100 805.050 414.900 806.850 ;
        RECT 437.400 805.050 438.300 815.400 ;
        RECT 460.500 810.000 462.300 818.400 ;
        RECT 459.000 808.800 462.300 810.000 ;
        RECT 467.100 809.400 468.900 819.000 ;
        RECT 472.950 816.450 475.050 817.050 ;
        RECT 478.950 816.450 481.050 817.050 ;
        RECT 472.950 815.550 481.050 816.450 ;
        RECT 472.950 814.950 475.050 815.550 ;
        RECT 478.950 814.950 481.050 815.550 ;
        RECT 485.100 815.400 486.900 819.000 ;
        RECT 488.100 815.400 489.900 818.400 ;
        RECT 491.100 815.400 492.900 819.000 ;
        RECT 509.100 815.400 510.900 819.000 ;
        RECT 512.100 815.400 513.900 818.400 ;
        RECT 515.100 815.400 516.900 819.000 ;
        RECT 533.100 815.400 534.900 818.400 ;
        RECT 536.100 815.400 537.900 819.000 ;
        RECT 554.100 815.400 555.900 818.400 ;
        RECT 557.100 815.400 558.900 819.000 ;
        RECT 575.100 815.400 576.900 819.000 ;
        RECT 578.100 815.400 579.900 818.400 ;
        RECT 581.100 815.400 582.900 819.000 ;
        RECT 459.000 805.050 459.900 808.800 ;
        RECT 461.100 805.050 462.900 806.850 ;
        RECT 467.100 805.050 468.900 806.850 ;
        RECT 488.400 805.050 489.300 815.400 ;
        RECT 512.400 805.050 513.300 815.400 ;
        RECT 533.700 805.050 534.900 815.400 ;
        RECT 554.700 805.050 555.900 815.400 ;
        RECT 578.400 805.050 579.300 815.400 ;
        RECT 599.400 812.400 601.200 819.000 ;
        RECT 604.500 811.200 606.300 818.400 ;
        RECT 623.700 815.400 625.500 819.000 ;
        RECT 626.700 813.600 628.500 818.400 ;
        RECT 586.950 810.450 589.050 811.050 ;
        RECT 598.950 810.450 601.050 811.050 ;
        RECT 586.950 809.550 601.050 810.450 ;
        RECT 586.950 808.950 589.050 809.550 ;
        RECT 598.950 808.950 601.050 809.550 ;
        RECT 602.100 810.300 606.300 811.200 ;
        RECT 623.400 812.400 628.500 813.600 ;
        RECT 631.200 812.400 633.000 819.000 ;
        RECT 599.250 805.050 601.050 806.850 ;
        RECT 602.100 805.050 603.300 810.300 ;
        RECT 605.100 805.050 606.900 806.850 ;
        RECT 623.400 805.050 624.300 812.400 ;
        RECT 650.700 811.200 652.500 818.400 ;
        RECT 655.800 812.400 657.600 819.000 ;
        RECT 674.100 812.400 675.900 818.400 ;
        RECT 677.100 813.000 678.900 819.000 ;
        RECT 683.700 818.400 684.900 819.000 ;
        RECT 680.100 815.400 681.900 818.400 ;
        RECT 683.100 815.400 684.900 818.400 ;
        RECT 650.700 810.300 654.900 811.200 ;
        RECT 625.950 805.050 627.750 806.850 ;
        RECT 632.100 805.050 633.900 806.850 ;
        RECT 650.100 805.050 651.900 806.850 ;
        RECT 653.700 805.050 654.900 810.300 ;
        RECT 655.950 805.050 657.750 806.850 ;
        RECT 674.100 805.050 675.000 812.400 ;
        RECT 680.700 811.200 681.600 815.400 ;
        RECT 701.100 812.400 702.900 818.400 ;
        RECT 676.200 810.300 681.600 811.200 ;
        RECT 701.700 810.300 702.900 812.400 ;
        RECT 704.100 813.300 705.900 818.400 ;
        RECT 707.100 814.200 708.900 819.000 ;
        RECT 710.100 813.300 711.900 818.400 ;
        RECT 704.100 811.950 711.900 813.300 ;
        RECT 728.100 810.600 729.900 818.400 ;
        RECT 732.600 812.400 734.400 819.000 ;
        RECT 735.600 814.200 737.400 818.400 ;
        RECT 735.600 812.400 738.300 814.200 ;
        RECT 734.700 810.600 736.500 811.500 ;
        RECT 676.200 809.400 678.300 810.300 ;
        RECT 701.700 809.400 705.300 810.300 ;
        RECT 728.100 809.700 736.500 810.600 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 361.950 802.950 364.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 382.950 802.950 385.050 805.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 674.100 802.950 676.200 805.050 ;
        RECT 208.500 799.950 210.900 802.050 ;
        RECT 202.800 789.600 204.000 790.500 ;
        RECT 208.500 789.600 210.000 799.950 ;
        RECT 231.000 790.800 231.900 802.950 ;
        RECT 236.100 801.150 237.900 802.950 ;
        RECT 247.950 801.450 250.050 802.050 ;
        RECT 253.950 801.450 256.050 802.050 ;
        RECT 247.950 800.550 256.050 801.450 ;
        RECT 247.950 799.950 250.050 800.550 ;
        RECT 253.950 799.950 256.050 800.550 ;
        RECT 231.000 789.900 237.600 790.800 ;
        RECT 231.000 789.600 231.900 789.900 ;
        RECT 178.200 783.000 180.000 789.600 ;
        RECT 181.200 783.600 183.000 789.600 ;
        RECT 184.200 786.600 186.300 788.700 ;
        RECT 187.200 786.600 189.300 788.700 ;
        RECT 190.200 786.600 192.300 788.700 ;
        RECT 184.200 783.600 186.000 786.600 ;
        RECT 187.200 783.600 189.000 786.600 ;
        RECT 190.200 783.600 192.000 786.600 ;
        RECT 193.200 783.000 195.000 789.600 ;
        RECT 196.200 783.600 198.000 789.600 ;
        RECT 199.200 783.000 201.000 789.600 ;
        RECT 202.200 783.600 204.000 789.600 ;
        RECT 205.200 783.000 207.000 789.600 ;
        RECT 208.500 783.600 210.300 789.600 ;
        RECT 211.500 783.000 213.300 789.600 ;
        RECT 230.100 783.600 231.900 789.600 ;
        RECT 236.100 789.600 237.600 789.900 ;
        RECT 257.700 789.600 258.900 802.950 ;
        RECT 260.100 801.150 261.900 802.950 ;
        RECT 281.700 789.600 282.900 802.950 ;
        RECT 302.100 801.150 303.900 802.950 ;
        RECT 308.700 795.600 309.900 802.950 ;
        RECT 329.250 801.150 331.050 802.950 ;
        RECT 310.950 798.450 313.050 799.050 ;
        RECT 316.950 798.450 319.050 799.050 ;
        RECT 310.950 797.550 319.050 798.450 ;
        RECT 310.950 796.950 313.050 797.550 ;
        RECT 316.950 796.950 319.050 797.550 ;
        RECT 332.400 795.600 333.300 802.950 ;
        RECT 335.100 801.150 336.900 802.950 ;
        RECT 356.100 801.150 357.900 802.950 ;
        RECT 233.100 783.000 234.900 789.000 ;
        RECT 236.100 783.600 237.900 789.600 ;
        RECT 239.100 783.000 240.900 789.600 ;
        RECT 257.100 783.600 258.900 789.600 ;
        RECT 260.100 783.000 261.900 789.600 ;
        RECT 278.100 783.000 279.900 789.600 ;
        RECT 281.100 783.600 282.900 789.600 ;
        RECT 284.100 783.000 285.900 789.600 ;
        RECT 302.400 783.000 304.200 795.600 ;
        RECT 307.500 794.100 309.900 795.600 ;
        RECT 307.500 783.600 309.300 794.100 ;
        RECT 310.200 791.100 312.000 792.900 ;
        RECT 310.500 783.000 312.300 789.600 ;
        RECT 329.100 783.000 330.900 795.600 ;
        RECT 332.400 794.400 336.000 795.600 ;
        RECT 334.200 783.600 336.000 794.400 ;
        RECT 352.950 795.450 355.050 796.050 ;
        RECT 358.950 795.450 361.050 796.050 ;
        RECT 352.950 794.550 361.050 795.450 ;
        RECT 352.950 793.950 355.050 794.550 ;
        RECT 358.950 793.950 361.050 794.550 ;
        RECT 362.100 790.800 363.000 802.950 ;
        RECT 383.100 801.150 384.900 802.950 ;
        RECT 389.100 790.800 390.000 802.950 ;
        RECT 410.100 795.600 411.300 802.950 ;
        RECT 416.100 801.150 417.900 802.950 ;
        RECT 434.250 801.150 436.050 802.950 ;
        RECT 437.400 795.600 438.300 802.950 ;
        RECT 440.100 801.150 441.900 802.950 ;
        RECT 410.100 794.100 412.500 795.600 ;
        RECT 408.000 791.100 409.800 792.900 ;
        RECT 356.400 789.900 363.000 790.800 ;
        RECT 356.400 789.600 357.900 789.900 ;
        RECT 353.100 783.000 354.900 789.600 ;
        RECT 356.100 783.600 357.900 789.600 ;
        RECT 362.100 789.600 363.000 789.900 ;
        RECT 383.400 789.900 390.000 790.800 ;
        RECT 383.400 789.600 384.900 789.900 ;
        RECT 359.100 783.000 360.900 789.000 ;
        RECT 362.100 783.600 363.900 789.600 ;
        RECT 380.100 783.000 381.900 789.600 ;
        RECT 383.100 783.600 384.900 789.600 ;
        RECT 389.100 789.600 390.000 789.900 ;
        RECT 386.100 783.000 387.900 789.000 ;
        RECT 389.100 783.600 390.900 789.600 ;
        RECT 407.700 783.000 409.500 789.600 ;
        RECT 410.700 783.600 412.500 794.100 ;
        RECT 415.800 783.000 417.600 795.600 ;
        RECT 434.100 783.000 435.900 795.600 ;
        RECT 437.400 794.400 441.000 795.600 ;
        RECT 439.200 783.600 441.000 794.400 ;
        RECT 459.000 790.800 459.900 802.950 ;
        RECT 464.100 801.150 465.900 802.950 ;
        RECT 485.250 801.150 487.050 802.950 ;
        RECT 488.400 795.600 489.300 802.950 ;
        RECT 491.100 801.150 492.900 802.950 ;
        RECT 509.250 801.150 511.050 802.950 ;
        RECT 512.400 795.600 513.300 802.950 ;
        RECT 515.100 801.150 516.900 802.950 ;
        RECT 459.000 789.900 465.600 790.800 ;
        RECT 459.000 789.600 459.900 789.900 ;
        RECT 458.100 783.600 459.900 789.600 ;
        RECT 464.100 789.600 465.600 789.900 ;
        RECT 461.100 783.000 462.900 789.000 ;
        RECT 464.100 783.600 465.900 789.600 ;
        RECT 467.100 783.000 468.900 789.600 ;
        RECT 485.100 783.000 486.900 795.600 ;
        RECT 488.400 794.400 492.000 795.600 ;
        RECT 490.200 783.600 492.000 794.400 ;
        RECT 509.100 783.000 510.900 795.600 ;
        RECT 512.400 794.400 516.000 795.600 ;
        RECT 514.200 783.600 516.000 794.400 ;
        RECT 533.700 789.600 534.900 802.950 ;
        RECT 536.100 801.150 537.900 802.950 ;
        RECT 554.700 789.600 555.900 802.950 ;
        RECT 557.100 801.150 558.900 802.950 ;
        RECT 575.250 801.150 577.050 802.950 ;
        RECT 578.400 795.600 579.300 802.950 ;
        RECT 581.100 801.150 582.900 802.950 ;
        RECT 533.100 783.600 534.900 789.600 ;
        RECT 536.100 783.000 537.900 789.600 ;
        RECT 554.100 783.600 555.900 789.600 ;
        RECT 557.100 783.000 558.900 789.600 ;
        RECT 575.100 783.000 576.900 795.600 ;
        RECT 578.400 794.400 582.000 795.600 ;
        RECT 580.200 783.600 582.000 794.400 ;
        RECT 602.100 789.600 603.300 802.950 ;
        RECT 623.400 795.600 624.300 802.950 ;
        RECT 628.950 801.150 630.750 802.950 ;
        RECT 599.100 783.000 600.900 789.600 ;
        RECT 602.100 783.600 603.900 789.600 ;
        RECT 605.100 783.000 606.900 789.600 ;
        RECT 623.100 783.600 624.900 795.600 ;
        RECT 626.100 794.700 633.900 795.600 ;
        RECT 626.100 783.600 627.900 794.700 ;
        RECT 629.100 783.000 630.900 793.800 ;
        RECT 632.100 783.600 633.900 794.700 ;
        RECT 653.700 789.600 654.900 802.950 ;
        RECT 675.000 795.600 676.200 802.950 ;
        RECT 677.400 798.900 678.300 809.400 ;
        RECT 682.800 805.050 684.600 806.850 ;
        RECT 701.100 805.050 702.900 806.850 ;
        RECT 704.100 805.050 705.300 809.400 ;
        RECT 707.100 805.050 708.900 806.850 ;
        RECT 728.250 805.050 730.050 806.850 ;
        RECT 679.500 802.950 681.600 805.050 ;
        RECT 682.800 802.950 684.900 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 728.100 802.950 730.200 805.050 ;
        RECT 679.200 801.150 681.000 802.950 ;
        RECT 677.100 798.300 678.900 798.900 ;
        RECT 677.100 797.100 684.900 798.300 ;
        RECT 683.700 795.600 684.900 797.100 ;
        RECT 675.000 794.100 677.400 795.600 ;
        RECT 650.100 783.000 651.900 789.600 ;
        RECT 653.100 783.600 654.900 789.600 ;
        RECT 656.100 783.000 657.900 789.600 ;
        RECT 675.600 783.600 677.400 794.100 ;
        RECT 678.600 783.000 680.400 795.600 ;
        RECT 683.100 783.600 684.900 795.600 ;
        RECT 704.100 795.600 705.300 802.950 ;
        RECT 710.100 801.150 711.900 802.950 ;
        RECT 706.950 798.450 709.050 799.050 ;
        RECT 718.950 798.450 721.050 799.050 ;
        RECT 706.950 797.550 721.050 798.450 ;
        RECT 706.950 796.950 709.050 797.550 ;
        RECT 718.950 796.950 721.050 797.550 ;
        RECT 704.100 794.100 706.500 795.600 ;
        RECT 702.000 791.100 703.800 792.900 ;
        RECT 701.700 783.000 703.500 789.600 ;
        RECT 704.700 783.600 706.500 794.100 ;
        RECT 709.800 783.000 711.600 795.600 ;
        RECT 731.100 789.600 732.000 809.700 ;
        RECT 737.400 805.050 738.300 812.400 ;
        RECT 757.500 810.000 759.300 818.400 ;
        RECT 756.000 808.800 759.300 810.000 ;
        RECT 764.100 809.400 765.900 819.000 ;
        RECT 784.500 810.000 786.300 818.400 ;
        RECT 783.000 808.800 786.300 810.000 ;
        RECT 791.100 809.400 792.900 819.000 ;
        RECT 809.100 809.400 810.900 819.000 ;
        RECT 815.700 810.000 817.500 818.400 ;
        RECT 837.000 812.400 838.800 819.000 ;
        RECT 841.500 813.600 843.300 818.400 ;
        RECT 844.500 815.400 846.300 819.000 ;
        RECT 841.500 812.400 846.600 813.600 ;
        RECT 823.950 810.450 826.050 811.050 ;
        RECT 838.950 810.450 841.050 811.050 ;
        RECT 815.700 808.800 819.000 810.000 ;
        RECT 823.950 809.550 841.050 810.450 ;
        RECT 823.950 808.950 826.050 809.550 ;
        RECT 838.950 808.950 841.050 809.550 ;
        RECT 756.000 805.050 756.900 808.800 ;
        RECT 758.100 805.050 759.900 806.850 ;
        RECT 764.100 805.050 765.900 806.850 ;
        RECT 783.000 805.050 783.900 808.800 ;
        RECT 793.950 807.450 798.000 808.050 ;
        RECT 785.100 805.050 786.900 806.850 ;
        RECT 791.100 805.050 792.900 806.850 ;
        RECT 793.950 805.950 798.450 807.450 ;
        RECT 733.500 802.950 735.600 805.050 ;
        RECT 736.800 802.950 738.900 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 763.950 802.950 766.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 733.200 801.150 735.000 802.950 ;
        RECT 737.400 795.600 738.300 802.950 ;
        RECT 728.100 783.000 729.900 789.600 ;
        RECT 731.100 783.600 732.900 789.600 ;
        RECT 734.100 783.000 735.900 795.000 ;
        RECT 737.100 783.600 738.900 795.600 ;
        RECT 756.000 790.800 756.900 802.950 ;
        RECT 761.100 801.150 762.900 802.950 ;
        RECT 783.000 790.800 783.900 802.950 ;
        RECT 788.100 801.150 789.900 802.950 ;
        RECT 797.550 798.450 798.450 805.950 ;
        RECT 809.100 805.050 810.900 806.850 ;
        RECT 815.100 805.050 816.900 806.850 ;
        RECT 818.100 805.050 819.000 808.800 ;
        RECT 836.100 805.050 837.900 806.850 ;
        RECT 842.250 805.050 844.050 806.850 ;
        RECT 845.700 805.050 846.600 812.400 ;
        RECT 863.100 813.300 864.900 818.400 ;
        RECT 866.100 814.200 867.900 819.000 ;
        RECT 869.100 813.300 870.900 818.400 ;
        RECT 863.100 811.950 870.900 813.300 ;
        RECT 872.100 812.400 873.900 818.400 ;
        RECT 890.100 815.400 891.900 819.000 ;
        RECT 893.100 815.400 894.900 818.400 ;
        RECT 896.100 815.400 897.900 819.000 ;
        RECT 872.100 810.300 873.300 812.400 ;
        RECT 869.700 809.400 873.300 810.300 ;
        RECT 877.950 810.450 880.050 811.050 ;
        RECT 889.950 810.450 892.050 811.050 ;
        RECT 877.950 809.550 892.050 810.450 ;
        RECT 866.100 805.050 867.900 806.850 ;
        RECT 869.700 805.050 870.900 809.400 ;
        RECT 877.950 808.950 880.050 809.550 ;
        RECT 889.950 808.950 892.050 809.550 ;
        RECT 872.100 805.050 873.900 806.850 ;
        RECT 893.700 805.050 894.600 815.400 ;
        RECT 914.700 811.200 916.500 818.400 ;
        RECT 919.800 812.400 921.600 819.000 ;
        RECT 935.100 812.400 936.900 818.400 ;
        RECT 895.950 810.450 898.050 811.050 ;
        RECT 910.950 810.450 913.050 811.050 ;
        RECT 895.950 809.550 913.050 810.450 ;
        RECT 914.700 810.300 918.900 811.200 ;
        RECT 895.950 808.950 898.050 809.550 ;
        RECT 910.950 808.950 913.050 809.550 ;
        RECT 914.100 805.050 915.900 806.850 ;
        RECT 917.700 805.050 918.900 810.300 ;
        RECT 935.700 810.300 936.900 812.400 ;
        RECT 938.100 813.300 939.900 818.400 ;
        RECT 941.100 814.200 942.900 819.000 ;
        RECT 944.100 813.300 945.900 818.400 ;
        RECT 938.100 811.950 945.900 813.300 ;
        RECT 935.700 809.400 939.300 810.300 ;
        RECT 964.500 810.000 966.300 818.400 ;
        RECT 919.950 805.050 921.750 806.850 ;
        RECT 935.100 805.050 936.900 806.850 ;
        RECT 938.100 805.050 939.300 809.400 ;
        RECT 963.000 808.800 966.300 810.000 ;
        RECT 971.100 809.400 972.900 819.000 ;
        RECT 989.700 811.200 991.500 818.400 ;
        RECT 994.800 812.400 996.600 819.000 ;
        RECT 1013.100 812.400 1014.900 818.400 ;
        RECT 989.700 810.300 993.900 811.200 ;
        RECT 957.000 807.450 961.050 808.050 ;
        RECT 941.100 805.050 942.900 806.850 ;
        RECT 956.550 805.950 961.050 807.450 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 841.950 802.950 844.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 865.950 802.950 868.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 895.950 802.950 898.050 805.050 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 919.950 802.950 922.050 805.050 ;
        RECT 934.950 802.950 937.050 805.050 ;
        RECT 937.950 802.950 940.050 805.050 ;
        RECT 940.950 802.950 943.050 805.050 ;
        RECT 943.950 802.950 946.050 805.050 ;
        RECT 812.100 801.150 813.900 802.950 ;
        RECT 808.950 798.450 811.050 799.050 ;
        RECT 797.550 797.550 811.050 798.450 ;
        RECT 808.950 796.950 811.050 797.550 ;
        RECT 796.950 795.450 799.050 796.050 ;
        RECT 814.950 795.450 817.050 799.050 ;
        RECT 796.950 795.000 817.050 795.450 ;
        RECT 796.950 794.550 816.450 795.000 ;
        RECT 796.950 793.950 799.050 794.550 ;
        RECT 818.100 790.800 819.000 802.950 ;
        RECT 839.250 801.150 841.050 802.950 ;
        RECT 820.950 798.450 823.050 799.050 ;
        RECT 835.950 798.450 838.050 799.050 ;
        RECT 820.950 797.550 838.050 798.450 ;
        RECT 820.950 796.950 823.050 797.550 ;
        RECT 835.950 796.950 838.050 797.550 ;
        RECT 845.700 795.600 846.600 802.950 ;
        RECT 863.100 801.150 864.900 802.950 ;
        RECT 847.950 798.450 850.050 799.050 ;
        RECT 865.950 798.450 868.050 799.050 ;
        RECT 847.950 797.550 868.050 798.450 ;
        RECT 847.950 796.950 850.050 797.550 ;
        RECT 865.950 796.950 868.050 797.550 ;
        RECT 869.700 795.600 870.900 802.950 ;
        RECT 890.100 801.150 891.900 802.950 ;
        RECT 880.950 798.450 883.050 799.050 ;
        RECT 889.950 798.450 892.050 799.050 ;
        RECT 880.950 797.550 892.050 798.450 ;
        RECT 880.950 796.950 883.050 797.550 ;
        RECT 889.950 796.950 892.050 797.550 ;
        RECT 893.700 795.600 894.600 802.950 ;
        RECT 895.950 801.150 897.750 802.950 ;
        RECT 756.000 789.900 762.600 790.800 ;
        RECT 756.000 789.600 756.900 789.900 ;
        RECT 755.100 783.600 756.900 789.600 ;
        RECT 761.100 789.600 762.600 789.900 ;
        RECT 783.000 789.900 789.600 790.800 ;
        RECT 783.000 789.600 783.900 789.900 ;
        RECT 758.100 783.000 759.900 789.000 ;
        RECT 761.100 783.600 762.900 789.600 ;
        RECT 764.100 783.000 765.900 789.600 ;
        RECT 782.100 783.600 783.900 789.600 ;
        RECT 788.100 789.600 789.600 789.900 ;
        RECT 812.400 789.900 819.000 790.800 ;
        RECT 812.400 789.600 813.900 789.900 ;
        RECT 785.100 783.000 786.900 789.000 ;
        RECT 788.100 783.600 789.900 789.600 ;
        RECT 791.100 783.000 792.900 789.600 ;
        RECT 809.100 783.000 810.900 789.600 ;
        RECT 812.100 783.600 813.900 789.600 ;
        RECT 818.100 789.600 819.000 789.900 ;
        RECT 836.100 794.700 843.900 795.600 ;
        RECT 815.100 783.000 816.900 789.000 ;
        RECT 818.100 783.600 819.900 789.600 ;
        RECT 836.100 783.600 837.900 794.700 ;
        RECT 839.100 783.000 840.900 793.800 ;
        RECT 842.100 783.600 843.900 794.700 ;
        RECT 845.100 783.600 846.900 795.600 ;
        RECT 863.400 783.000 865.200 795.600 ;
        RECT 868.500 794.100 870.900 795.600 ;
        RECT 891.000 794.400 894.600 795.600 ;
        RECT 868.500 783.600 870.300 794.100 ;
        RECT 871.200 791.100 873.000 792.900 ;
        RECT 871.500 783.000 873.300 789.600 ;
        RECT 891.000 783.600 892.800 794.400 ;
        RECT 896.100 783.000 897.900 795.600 ;
        RECT 917.700 789.600 918.900 802.950 ;
        RECT 938.100 795.600 939.300 802.950 ;
        RECT 944.100 801.150 945.900 802.950 ;
        RECT 956.550 802.050 957.450 805.950 ;
        RECT 963.000 805.050 963.900 808.800 ;
        RECT 965.100 805.050 966.900 806.850 ;
        RECT 971.100 805.050 972.900 806.850 ;
        RECT 989.100 805.050 990.900 806.850 ;
        RECT 992.700 805.050 993.900 810.300 ;
        RECT 1003.950 808.950 1006.050 811.050 ;
        RECT 1013.700 810.300 1014.900 812.400 ;
        RECT 1016.100 813.300 1017.900 818.400 ;
        RECT 1019.100 814.200 1020.900 819.000 ;
        RECT 1022.100 813.300 1023.900 818.400 ;
        RECT 1037.100 815.400 1038.900 818.400 ;
        RECT 1040.100 815.400 1041.900 819.000 ;
        RECT 1016.100 811.950 1023.900 813.300 ;
        RECT 1013.700 809.400 1017.300 810.300 ;
        RECT 997.950 807.450 1002.000 808.050 ;
        RECT 994.950 805.050 996.750 806.850 ;
        RECT 997.950 805.950 1002.450 807.450 ;
        RECT 961.950 802.950 964.050 805.050 ;
        RECT 964.950 802.950 967.050 805.050 ;
        RECT 967.950 802.950 970.050 805.050 ;
        RECT 970.950 802.950 973.050 805.050 ;
        RECT 988.950 802.950 991.050 805.050 ;
        RECT 991.950 802.950 994.050 805.050 ;
        RECT 994.950 802.950 997.050 805.050 ;
        RECT 956.550 800.550 961.050 802.050 ;
        RECT 957.000 799.950 961.050 800.550 ;
        RECT 940.950 798.450 943.050 799.050 ;
        RECT 952.950 798.450 955.050 799.050 ;
        RECT 940.950 797.550 955.050 798.450 ;
        RECT 940.950 796.950 943.050 797.550 ;
        RECT 952.950 796.950 955.050 797.550 ;
        RECT 938.100 794.100 940.500 795.600 ;
        RECT 936.000 791.100 937.800 792.900 ;
        RECT 914.100 783.000 915.900 789.600 ;
        RECT 917.100 783.600 918.900 789.600 ;
        RECT 920.100 783.000 921.900 789.600 ;
        RECT 935.700 783.000 937.500 789.600 ;
        RECT 938.700 783.600 940.500 794.100 ;
        RECT 943.800 783.000 945.600 795.600 ;
        RECT 963.000 790.800 963.900 802.950 ;
        RECT 968.100 801.150 969.900 802.950 ;
        RECT 964.950 795.450 967.050 796.050 ;
        RECT 979.950 795.450 982.050 796.050 ;
        RECT 964.950 794.550 982.050 795.450 ;
        RECT 964.950 793.950 967.050 794.550 ;
        RECT 979.950 793.950 982.050 794.550 ;
        RECT 963.000 789.900 969.600 790.800 ;
        RECT 963.000 789.600 963.900 789.900 ;
        RECT 962.100 783.600 963.900 789.600 ;
        RECT 968.100 789.600 969.600 789.900 ;
        RECT 992.700 789.600 993.900 802.950 ;
        RECT 1001.550 802.050 1002.450 805.950 ;
        RECT 997.950 800.550 1002.450 802.050 ;
        RECT 997.950 799.950 1002.000 800.550 ;
        RECT 1004.550 798.450 1005.450 808.950 ;
        RECT 1008.000 807.450 1012.050 808.050 ;
        RECT 1007.550 805.950 1012.050 807.450 ;
        RECT 1007.550 802.050 1008.450 805.950 ;
        RECT 1013.100 805.050 1014.900 806.850 ;
        RECT 1016.100 805.050 1017.300 809.400 ;
        RECT 1024.950 807.450 1029.000 808.050 ;
        RECT 1019.100 805.050 1020.900 806.850 ;
        RECT 1024.950 805.950 1029.450 807.450 ;
        RECT 1012.950 802.950 1015.050 805.050 ;
        RECT 1015.950 802.950 1018.050 805.050 ;
        RECT 1018.950 802.950 1021.050 805.050 ;
        RECT 1021.950 802.950 1024.050 805.050 ;
        RECT 1007.550 800.550 1012.050 802.050 ;
        RECT 1008.000 799.950 1012.050 800.550 ;
        RECT 1012.950 798.450 1015.050 799.050 ;
        RECT 1004.550 797.550 1015.050 798.450 ;
        RECT 1012.950 796.950 1015.050 797.550 ;
        RECT 1016.100 795.600 1017.300 802.950 ;
        RECT 1022.100 801.150 1023.900 802.950 ;
        RECT 1021.950 798.450 1024.050 799.050 ;
        RECT 1028.550 798.450 1029.450 805.950 ;
        RECT 1037.700 805.050 1038.900 815.400 ;
        RECT 1036.950 802.950 1039.050 805.050 ;
        RECT 1039.950 802.950 1042.050 805.050 ;
        RECT 1021.950 797.550 1029.450 798.450 ;
        RECT 1021.950 796.950 1024.050 797.550 ;
        RECT 1016.100 794.100 1018.500 795.600 ;
        RECT 1014.000 791.100 1015.800 792.900 ;
        RECT 965.100 783.000 966.900 789.000 ;
        RECT 968.100 783.600 969.900 789.600 ;
        RECT 971.100 783.000 972.900 789.600 ;
        RECT 989.100 783.000 990.900 789.600 ;
        RECT 992.100 783.600 993.900 789.600 ;
        RECT 995.100 783.000 996.900 789.600 ;
        RECT 1013.700 783.000 1015.500 789.600 ;
        RECT 1016.700 783.600 1018.500 794.100 ;
        RECT 1021.800 783.000 1023.600 795.600 ;
        RECT 1037.700 789.600 1038.900 802.950 ;
        RECT 1040.100 801.150 1041.900 802.950 ;
        RECT 1037.100 783.600 1038.900 789.600 ;
        RECT 1040.100 783.000 1041.900 789.600 ;
        RECT 17.100 767.400 18.900 779.400 ;
        RECT 20.100 769.200 21.900 780.000 ;
        RECT 23.100 773.400 24.900 779.400 ;
        RECT 17.100 760.050 18.300 767.400 ;
        RECT 23.700 766.500 24.900 773.400 ;
        RECT 41.100 778.500 48.900 779.400 ;
        RECT 41.100 769.200 42.900 778.500 ;
        RECT 44.100 769.800 45.900 777.600 ;
        RECT 19.200 765.600 24.900 766.500 ;
        RECT 19.200 764.700 21.000 765.600 ;
        RECT 17.100 757.950 19.200 760.050 ;
        RECT 17.100 750.600 18.300 757.950 ;
        RECT 20.100 753.300 21.000 764.700 ;
        RECT 22.800 760.050 24.600 761.850 ;
        RECT 44.700 760.050 45.900 769.800 ;
        RECT 47.100 769.800 48.900 778.500 ;
        RECT 50.100 778.500 57.900 779.400 ;
        RECT 50.100 770.700 51.900 778.500 ;
        RECT 53.100 769.800 54.900 777.600 ;
        RECT 47.100 768.900 54.900 769.800 ;
        RECT 56.100 769.500 57.900 778.500 ;
        RECT 59.100 770.400 60.900 780.000 ;
        RECT 62.100 769.500 63.900 779.400 ;
        RECT 56.100 768.600 63.900 769.500 ;
        RECT 80.100 778.500 87.900 779.400 ;
        RECT 80.100 769.200 81.900 778.500 ;
        RECT 83.100 769.800 84.900 777.600 ;
        RECT 49.950 760.050 51.750 761.850 ;
        RECT 59.100 760.050 60.900 761.850 ;
        RECT 83.700 760.050 84.900 769.800 ;
        RECT 86.100 769.800 87.900 778.500 ;
        RECT 89.100 778.500 96.900 779.400 ;
        RECT 89.100 770.700 90.900 778.500 ;
        RECT 92.100 769.800 93.900 777.600 ;
        RECT 86.100 768.900 93.900 769.800 ;
        RECT 95.100 769.500 96.900 778.500 ;
        RECT 98.100 770.400 99.900 780.000 ;
        RECT 101.100 769.500 102.900 779.400 ;
        RECT 95.100 768.600 102.900 769.500 ;
        RECT 120.000 768.600 121.800 779.400 ;
        RECT 120.000 767.400 123.600 768.600 ;
        RECT 125.100 767.400 126.900 780.000 ;
        RECT 143.700 773.400 145.500 780.000 ;
        RECT 144.000 770.100 145.800 771.900 ;
        RECT 146.700 768.900 148.500 779.400 ;
        RECT 146.100 767.400 148.500 768.900 ;
        RECT 151.800 767.400 153.600 780.000 ;
        RECT 170.100 773.400 171.900 780.000 ;
        RECT 173.100 773.400 174.900 779.400 ;
        RECT 88.950 760.050 90.750 761.850 ;
        RECT 98.100 760.050 99.900 761.850 ;
        RECT 119.100 760.050 120.900 761.850 ;
        RECT 122.700 760.050 123.600 767.400 ;
        RECT 124.950 760.050 126.750 761.850 ;
        RECT 146.100 760.050 147.300 767.400 ;
        RECT 152.100 760.050 153.900 761.850 ;
        RECT 170.100 760.050 171.900 761.850 ;
        RECT 173.100 760.050 174.300 773.400 ;
        RECT 191.400 767.400 193.200 780.000 ;
        RECT 196.500 768.900 198.300 779.400 ;
        RECT 199.500 773.400 201.300 780.000 ;
        RECT 218.700 773.400 220.500 780.000 ;
        RECT 199.200 770.100 201.000 771.900 ;
        RECT 219.000 770.100 220.800 771.900 ;
        RECT 221.700 768.900 223.500 779.400 ;
        RECT 196.500 767.400 198.900 768.900 ;
        RECT 191.100 760.050 192.900 761.850 ;
        RECT 197.700 760.050 198.900 767.400 ;
        RECT 221.100 767.400 223.500 768.900 ;
        RECT 226.800 767.400 228.600 780.000 ;
        RECT 246.000 768.600 247.800 779.400 ;
        RECT 246.000 767.400 249.600 768.600 ;
        RECT 251.100 767.400 252.900 780.000 ;
        RECT 269.100 767.400 270.900 779.400 ;
        RECT 272.100 768.300 273.900 779.400 ;
        RECT 275.100 769.200 276.900 780.000 ;
        RECT 278.100 768.300 279.900 779.400 ;
        RECT 272.100 767.400 279.900 768.300 ;
        RECT 296.100 767.400 297.900 780.000 ;
        RECT 202.950 765.450 205.050 766.050 ;
        RECT 208.950 765.450 211.050 766.050 ;
        RECT 202.950 764.550 211.050 765.450 ;
        RECT 202.950 763.950 205.050 764.550 ;
        RECT 208.950 763.950 211.050 764.550 ;
        RECT 221.100 760.050 222.300 767.400 ;
        RECT 227.100 760.050 228.900 761.850 ;
        RECT 245.100 760.050 246.900 761.850 ;
        RECT 248.700 760.050 249.600 767.400 ;
        RECT 250.950 760.050 252.750 761.850 ;
        RECT 269.400 760.050 270.300 767.400 ;
        RECT 299.100 766.500 300.900 779.400 ;
        RECT 302.100 767.400 303.900 780.000 ;
        RECT 305.100 766.500 306.900 779.400 ;
        RECT 308.100 767.400 309.900 780.000 ;
        RECT 311.100 766.500 312.900 779.400 ;
        RECT 314.100 767.400 315.900 780.000 ;
        RECT 317.100 766.500 318.900 779.400 ;
        RECT 320.100 767.400 321.900 780.000 ;
        RECT 339.600 768.900 341.400 779.400 ;
        RECT 339.000 767.400 341.400 768.900 ;
        RECT 342.600 767.400 344.400 780.000 ;
        RECT 347.100 767.400 348.900 779.400 ;
        RECT 365.100 767.400 366.900 780.000 ;
        RECT 370.200 768.600 372.000 779.400 ;
        RECT 368.400 767.400 372.000 768.600 ;
        RECT 389.100 767.400 390.900 779.400 ;
        RECT 393.600 767.400 395.400 780.000 ;
        RECT 396.600 768.900 398.400 779.400 ;
        RECT 396.600 767.400 399.000 768.900 ;
        RECT 416.400 767.400 418.200 780.000 ;
        RECT 421.500 768.900 423.300 779.400 ;
        RECT 424.500 773.400 426.300 780.000 ;
        RECT 424.200 770.100 426.000 771.900 ;
        RECT 421.500 767.400 423.900 768.900 ;
        RECT 443.100 767.400 444.900 779.400 ;
        RECT 446.100 768.300 447.900 779.400 ;
        RECT 449.100 769.200 450.900 780.000 ;
        RECT 452.100 768.300 453.900 779.400 ;
        RECT 470.100 773.400 471.900 779.400 ;
        RECT 473.100 773.400 474.900 780.000 ;
        RECT 446.100 767.400 453.900 768.300 ;
        RECT 298.050 765.300 300.900 766.500 ;
        RECT 303.000 765.300 306.900 766.500 ;
        RECT 309.000 765.300 312.900 766.500 ;
        RECT 315.000 765.300 318.900 766.500 ;
        RECT 274.950 760.050 276.750 761.850 ;
        RECT 298.050 760.050 299.100 765.300 ;
        RECT 22.500 757.950 24.600 760.050 ;
        RECT 44.400 757.950 46.500 760.050 ;
        RECT 49.950 757.950 52.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 59.100 757.950 61.200 760.050 ;
        RECT 83.400 757.950 85.500 760.050 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 91.950 757.950 94.050 760.050 ;
        RECT 98.100 757.950 100.200 760.050 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 172.950 757.950 175.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 199.950 757.950 202.050 760.050 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 220.950 757.950 223.050 760.050 ;
        RECT 223.950 757.950 226.050 760.050 ;
        RECT 226.950 757.950 229.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 247.950 757.950 250.050 760.050 ;
        RECT 250.950 757.950 253.050 760.050 ;
        RECT 268.950 757.950 271.050 760.050 ;
        RECT 271.950 757.950 274.050 760.050 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 298.050 757.950 301.200 760.050 ;
        RECT 19.200 752.400 21.000 753.300 ;
        RECT 19.200 751.500 24.900 752.400 ;
        RECT 17.100 744.600 18.900 750.600 ;
        RECT 20.100 744.000 21.900 750.600 ;
        RECT 23.700 747.600 24.900 751.500 ;
        RECT 44.700 749.400 45.900 757.950 ;
        RECT 53.250 756.150 55.050 757.950 ;
        RECT 52.950 753.450 55.050 754.050 ;
        RECT 76.950 753.450 79.050 754.050 ;
        RECT 52.950 752.550 79.050 753.450 ;
        RECT 52.950 751.950 55.050 752.550 ;
        RECT 76.950 751.950 79.050 752.550 ;
        RECT 83.700 749.400 84.900 757.950 ;
        RECT 92.250 756.150 94.050 757.950 ;
        RECT 91.950 753.450 94.050 754.050 ;
        RECT 118.950 753.450 121.050 754.050 ;
        RECT 91.950 752.550 121.050 753.450 ;
        RECT 91.950 751.950 94.050 752.550 ;
        RECT 118.950 751.950 121.050 752.550 ;
        RECT 97.950 750.450 100.050 751.050 ;
        RECT 115.950 750.450 118.050 751.050 ;
        RECT 97.950 749.550 118.050 750.450 ;
        RECT 44.700 748.500 57.300 749.400 ;
        RECT 83.700 748.500 96.300 749.400 ;
        RECT 97.950 748.950 100.050 749.550 ;
        RECT 115.950 748.950 118.050 749.550 ;
        RECT 23.100 744.600 24.900 747.600 ;
        RECT 49.200 747.600 50.100 748.500 ;
        RECT 56.400 747.600 57.300 748.500 ;
        RECT 88.200 747.600 89.100 748.500 ;
        RECT 95.400 747.600 96.300 748.500 ;
        RECT 122.700 747.600 123.600 757.950 ;
        RECT 143.100 756.150 144.900 757.950 ;
        RECT 146.100 753.600 147.300 757.950 ;
        RECT 149.100 756.150 150.900 757.950 ;
        RECT 143.700 752.700 147.300 753.600 ;
        RECT 143.700 750.600 144.900 752.700 ;
        RECT 49.200 744.600 51.900 747.600 ;
        RECT 53.100 744.000 54.900 747.600 ;
        RECT 56.100 744.600 57.900 747.600 ;
        RECT 59.100 744.000 61.200 747.600 ;
        RECT 88.200 744.600 90.900 747.600 ;
        RECT 92.100 744.000 93.900 747.600 ;
        RECT 95.100 744.600 96.900 747.600 ;
        RECT 98.100 744.000 100.200 747.600 ;
        RECT 119.100 744.000 120.900 747.600 ;
        RECT 122.100 744.600 123.900 747.600 ;
        RECT 125.100 744.000 126.900 747.600 ;
        RECT 143.100 744.600 144.900 750.600 ;
        RECT 146.100 749.700 153.900 751.050 ;
        RECT 146.100 744.600 147.900 749.700 ;
        RECT 149.100 744.000 150.900 748.800 ;
        RECT 152.100 744.600 153.900 749.700 ;
        RECT 173.100 747.600 174.300 757.950 ;
        RECT 194.100 756.150 195.900 757.950 ;
        RECT 197.700 753.600 198.900 757.950 ;
        RECT 200.100 756.150 201.900 757.950 ;
        RECT 218.100 756.150 219.900 757.950 ;
        RECT 221.100 753.600 222.300 757.950 ;
        RECT 224.100 756.150 225.900 757.950 ;
        RECT 197.700 752.700 201.300 753.600 ;
        RECT 191.100 749.700 198.900 751.050 ;
        RECT 170.100 744.000 171.900 747.600 ;
        RECT 173.100 744.600 174.900 747.600 ;
        RECT 191.100 744.600 192.900 749.700 ;
        RECT 194.100 744.000 195.900 748.800 ;
        RECT 197.100 744.600 198.900 749.700 ;
        RECT 200.100 750.600 201.300 752.700 ;
        RECT 218.700 752.700 222.300 753.600 ;
        RECT 218.700 750.600 219.900 752.700 ;
        RECT 200.100 744.600 201.900 750.600 ;
        RECT 218.100 744.600 219.900 750.600 ;
        RECT 221.100 749.700 228.900 751.050 ;
        RECT 221.100 744.600 222.900 749.700 ;
        RECT 224.100 744.000 225.900 748.800 ;
        RECT 227.100 744.600 228.900 749.700 ;
        RECT 248.700 747.600 249.600 757.950 ;
        RECT 269.400 750.600 270.300 757.950 ;
        RECT 271.950 756.150 273.750 757.950 ;
        RECT 278.100 756.150 279.900 757.950 ;
        RECT 298.050 752.700 299.100 757.950 ;
        RECT 300.000 754.800 301.800 755.400 ;
        RECT 303.000 754.800 304.200 765.300 ;
        RECT 300.000 753.600 304.200 754.800 ;
        RECT 306.000 754.800 307.800 755.400 ;
        RECT 309.000 754.800 310.200 765.300 ;
        RECT 306.000 753.600 310.200 754.800 ;
        RECT 312.000 754.800 313.800 755.400 ;
        RECT 315.000 754.800 316.200 765.300 ;
        RECT 339.000 760.050 340.200 767.400 ;
        RECT 347.700 765.900 348.900 767.400 ;
        RECT 341.100 764.700 348.900 765.900 ;
        RECT 341.100 764.100 342.900 764.700 ;
        RECT 317.100 757.950 319.200 760.050 ;
        RECT 317.400 756.150 319.200 757.950 ;
        RECT 338.100 757.950 340.200 760.050 ;
        RECT 312.000 753.600 316.200 754.800 ;
        RECT 303.000 752.700 304.200 753.600 ;
        RECT 309.000 752.700 310.200 753.600 ;
        RECT 315.000 752.700 316.200 753.600 ;
        RECT 298.050 751.500 300.900 752.700 ;
        RECT 303.000 751.500 306.900 752.700 ;
        RECT 309.000 751.500 312.900 752.700 ;
        RECT 315.000 751.500 318.900 752.700 ;
        RECT 269.400 749.400 274.500 750.600 ;
        RECT 245.100 744.000 246.900 747.600 ;
        RECT 248.100 744.600 249.900 747.600 ;
        RECT 251.100 744.000 252.900 747.600 ;
        RECT 269.700 744.000 271.500 747.600 ;
        RECT 272.700 744.600 274.500 749.400 ;
        RECT 277.200 744.000 279.000 750.600 ;
        RECT 296.100 744.000 297.900 750.600 ;
        RECT 299.100 744.600 300.900 751.500 ;
        RECT 302.100 744.000 303.900 750.600 ;
        RECT 305.100 744.600 306.900 751.500 ;
        RECT 308.100 744.000 309.900 750.600 ;
        RECT 311.100 744.600 312.900 751.500 ;
        RECT 314.100 744.000 315.900 750.600 ;
        RECT 317.100 744.600 318.900 751.500 ;
        RECT 338.100 750.600 339.000 757.950 ;
        RECT 341.400 753.600 342.300 764.100 ;
        RECT 343.200 760.050 345.000 761.850 ;
        RECT 365.250 760.050 367.050 761.850 ;
        RECT 368.400 760.050 369.300 767.400 ;
        RECT 389.100 765.900 390.300 767.400 ;
        RECT 389.100 764.700 396.900 765.900 ;
        RECT 395.100 764.100 396.900 764.700 ;
        RECT 371.100 760.050 372.900 761.850 ;
        RECT 393.000 760.050 394.800 761.850 ;
        RECT 343.500 757.950 345.600 760.050 ;
        RECT 346.800 757.950 348.900 760.050 ;
        RECT 364.950 757.950 367.050 760.050 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 389.100 757.950 391.200 760.050 ;
        RECT 392.400 757.950 394.500 760.050 ;
        RECT 346.800 756.150 348.600 757.950 ;
        RECT 340.200 752.700 342.300 753.600 ;
        RECT 340.200 751.800 345.600 752.700 ;
        RECT 320.100 744.000 321.900 750.600 ;
        RECT 338.100 744.600 339.900 750.600 ;
        RECT 341.100 744.000 342.900 750.000 ;
        RECT 344.700 747.600 345.600 751.800 ;
        RECT 368.400 747.600 369.300 757.950 ;
        RECT 389.400 756.150 391.200 757.950 ;
        RECT 395.700 753.600 396.600 764.100 ;
        RECT 397.800 760.050 399.000 767.400 ;
        RECT 416.100 760.050 417.900 761.850 ;
        RECT 422.700 760.050 423.900 767.400 ;
        RECT 439.950 762.450 442.050 763.050 ;
        RECT 431.550 761.550 442.050 762.450 ;
        RECT 397.800 757.950 399.900 760.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 418.950 757.950 421.050 760.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 395.700 752.700 397.800 753.600 ;
        RECT 392.400 751.800 397.800 752.700 ;
        RECT 392.400 747.600 393.300 751.800 ;
        RECT 399.000 750.600 399.900 757.950 ;
        RECT 419.100 756.150 420.900 757.950 ;
        RECT 422.700 753.600 423.900 757.950 ;
        RECT 425.100 756.150 426.900 757.950 ;
        RECT 431.550 753.900 432.450 761.550 ;
        RECT 439.950 760.950 442.050 761.550 ;
        RECT 443.400 760.050 444.300 767.400 ;
        RECT 448.950 765.450 451.050 766.050 ;
        RECT 460.950 765.450 463.050 766.050 ;
        RECT 448.950 764.550 463.050 765.450 ;
        RECT 448.950 763.950 451.050 764.550 ;
        RECT 460.950 763.950 463.050 764.550 ;
        RECT 448.950 760.050 450.750 761.850 ;
        RECT 470.700 760.050 471.900 773.400 ;
        RECT 492.600 768.900 494.400 779.400 ;
        RECT 492.000 767.400 494.400 768.900 ;
        RECT 495.600 767.400 497.400 780.000 ;
        RECT 500.100 767.400 501.900 779.400 ;
        RECT 518.100 767.400 519.900 780.000 ;
        RECT 523.200 768.600 525.000 779.400 ;
        RECT 521.400 767.400 525.000 768.600 ;
        RECT 542.100 767.400 543.900 780.000 ;
        RECT 547.200 768.600 549.000 779.400 ;
        RECT 545.400 767.400 549.000 768.600 ;
        RECT 566.400 767.400 568.200 780.000 ;
        RECT 571.500 768.900 573.300 779.400 ;
        RECT 574.500 773.400 576.300 780.000 ;
        RECT 574.200 770.100 576.000 771.900 ;
        RECT 571.500 767.400 573.900 768.900 ;
        RECT 593.100 767.400 594.900 779.400 ;
        RECT 596.100 768.300 597.900 779.400 ;
        RECT 599.100 769.200 600.900 780.000 ;
        RECT 602.100 768.300 603.900 779.400 ;
        RECT 596.100 767.400 603.900 768.300 ;
        RECT 620.100 767.400 621.900 780.000 ;
        RECT 625.200 768.600 627.000 779.400 ;
        RECT 644.100 773.400 645.900 779.400 ;
        RECT 647.100 774.000 648.900 780.000 ;
        RECT 623.400 767.400 627.000 768.600 ;
        RECT 645.000 773.100 645.900 773.400 ;
        RECT 650.100 773.400 651.900 779.400 ;
        RECT 653.100 773.400 654.900 780.000 ;
        RECT 671.100 773.400 672.900 780.000 ;
        RECT 674.100 773.400 675.900 779.400 ;
        RECT 677.100 773.400 678.900 780.000 ;
        RECT 650.100 773.100 651.600 773.400 ;
        RECT 645.000 772.200 651.600 773.100 ;
        RECT 473.100 760.050 474.900 761.850 ;
        RECT 492.000 760.050 493.200 767.400 ;
        RECT 500.700 765.900 501.900 767.400 ;
        RECT 494.100 764.700 501.900 765.900 ;
        RECT 494.100 764.100 495.900 764.700 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 491.100 757.950 493.200 760.050 ;
        RECT 422.700 752.700 426.300 753.600 ;
        RECT 344.100 744.600 345.900 747.600 ;
        RECT 347.100 744.600 348.900 747.600 ;
        RECT 347.700 744.000 348.900 744.600 ;
        RECT 365.100 744.000 366.900 747.600 ;
        RECT 368.100 744.600 369.900 747.600 ;
        RECT 371.100 744.000 372.900 747.600 ;
        RECT 389.100 744.600 390.900 747.600 ;
        RECT 392.100 744.600 393.900 747.600 ;
        RECT 389.100 744.000 390.300 744.600 ;
        RECT 395.100 744.000 396.900 750.000 ;
        RECT 398.100 744.600 399.900 750.600 ;
        RECT 416.100 749.700 423.900 751.050 ;
        RECT 416.100 744.600 417.900 749.700 ;
        RECT 419.100 744.000 420.900 748.800 ;
        RECT 422.100 744.600 423.900 749.700 ;
        RECT 425.100 750.600 426.300 752.700 ;
        RECT 430.950 751.800 433.050 753.900 ;
        RECT 443.400 750.600 444.300 757.950 ;
        RECT 445.950 756.150 447.750 757.950 ;
        RECT 452.100 756.150 453.900 757.950 ;
        RECT 425.100 744.600 426.900 750.600 ;
        RECT 443.400 749.400 448.500 750.600 ;
        RECT 443.700 744.000 445.500 747.600 ;
        RECT 446.700 744.600 448.500 749.400 ;
        RECT 451.200 744.000 453.000 750.600 ;
        RECT 470.700 747.600 471.900 757.950 ;
        RECT 472.950 753.450 475.050 753.750 ;
        RECT 478.950 753.450 481.050 754.050 ;
        RECT 472.950 752.550 481.050 753.450 ;
        RECT 472.950 751.650 475.050 752.550 ;
        RECT 478.950 751.950 481.050 752.550 ;
        RECT 491.100 750.600 492.000 757.950 ;
        RECT 494.400 753.600 495.300 764.100 ;
        RECT 496.200 760.050 498.000 761.850 ;
        RECT 518.250 760.050 520.050 761.850 ;
        RECT 521.400 760.050 522.300 767.400 ;
        RECT 524.100 760.050 525.900 761.850 ;
        RECT 542.250 760.050 544.050 761.850 ;
        RECT 545.400 760.050 546.300 767.400 ;
        RECT 548.100 760.050 549.900 761.850 ;
        RECT 566.100 760.050 567.900 761.850 ;
        RECT 572.700 760.050 573.900 767.400 ;
        RECT 583.950 765.450 586.050 766.050 ;
        RECT 589.950 765.450 592.050 766.050 ;
        RECT 583.950 764.550 592.050 765.450 ;
        RECT 583.950 763.950 586.050 764.550 ;
        RECT 589.950 763.950 592.050 764.550 ;
        RECT 593.400 760.050 594.300 767.400 ;
        RECT 598.950 760.050 600.750 761.850 ;
        RECT 620.250 760.050 622.050 761.850 ;
        RECT 623.400 760.050 624.300 767.400 ;
        RECT 626.100 760.050 627.900 761.850 ;
        RECT 645.000 760.050 645.900 772.200 ;
        RECT 650.100 760.050 651.900 761.850 ;
        RECT 674.700 760.050 675.900 773.400 ;
        RECT 695.100 767.400 696.900 780.000 ;
        RECT 700.200 768.600 702.000 779.400 ;
        RECT 698.400 767.400 702.000 768.600 ;
        RECT 719.100 767.400 720.900 780.000 ;
        RECT 722.100 767.400 723.900 779.400 ;
        RECT 740.100 767.400 741.900 780.000 ;
        RECT 745.200 768.600 747.000 779.400 ;
        RECT 743.400 767.400 747.000 768.600 ;
        RECT 764.100 767.400 765.900 779.400 ;
        RECT 767.100 767.400 768.900 780.000 ;
        RECT 786.000 768.600 787.800 779.400 ;
        RECT 786.000 767.400 789.600 768.600 ;
        RECT 791.100 767.400 792.900 780.000 ;
        RECT 809.100 773.400 810.900 780.000 ;
        RECT 812.100 773.400 813.900 779.400 ;
        RECT 815.100 773.400 816.900 780.000 ;
        RECT 695.250 760.050 697.050 761.850 ;
        RECT 698.400 760.050 699.300 767.400 ;
        RECT 703.950 762.450 708.000 763.050 ;
        RECT 701.100 760.050 702.900 761.850 ;
        RECT 703.950 760.950 708.450 762.450 ;
        RECT 496.500 757.950 498.600 760.050 ;
        RECT 499.800 757.950 501.900 760.050 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 652.950 757.950 655.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 499.800 756.150 501.600 757.950 ;
        RECT 493.200 752.700 495.300 753.600 ;
        RECT 493.200 751.800 498.600 752.700 ;
        RECT 470.100 744.600 471.900 747.600 ;
        RECT 473.100 744.000 474.900 747.600 ;
        RECT 491.100 744.600 492.900 750.600 ;
        RECT 494.100 744.000 495.900 750.000 ;
        RECT 497.700 747.600 498.600 751.800 ;
        RECT 521.400 747.600 522.300 757.950 ;
        RECT 529.950 753.450 532.050 754.050 ;
        RECT 541.950 753.450 544.050 754.050 ;
        RECT 529.950 752.550 544.050 753.450 ;
        RECT 529.950 751.950 532.050 752.550 ;
        RECT 541.950 751.950 544.050 752.550 ;
        RECT 545.400 747.600 546.300 757.950 ;
        RECT 569.100 756.150 570.900 757.950 ;
        RECT 572.700 753.600 573.900 757.950 ;
        RECT 575.100 756.150 576.900 757.950 ;
        RECT 572.700 752.700 576.300 753.600 ;
        RECT 566.100 749.700 573.900 751.050 ;
        RECT 497.100 744.600 498.900 747.600 ;
        RECT 500.100 744.600 501.900 747.600 ;
        RECT 500.700 744.000 501.900 744.600 ;
        RECT 518.100 744.000 519.900 747.600 ;
        RECT 521.100 744.600 522.900 747.600 ;
        RECT 524.100 744.000 525.900 747.600 ;
        RECT 542.100 744.000 543.900 747.600 ;
        RECT 545.100 744.600 546.900 747.600 ;
        RECT 548.100 744.000 549.900 747.600 ;
        RECT 566.100 744.600 567.900 749.700 ;
        RECT 569.100 744.000 570.900 748.800 ;
        RECT 572.100 744.600 573.900 749.700 ;
        RECT 575.100 750.600 576.300 752.700 ;
        RECT 593.400 750.600 594.300 757.950 ;
        RECT 595.950 756.150 597.750 757.950 ;
        RECT 602.100 756.150 603.900 757.950 ;
        RECT 575.100 744.600 576.900 750.600 ;
        RECT 593.400 749.400 598.500 750.600 ;
        RECT 593.700 744.000 595.500 747.600 ;
        RECT 596.700 744.600 598.500 749.400 ;
        RECT 601.200 744.000 603.000 750.600 ;
        RECT 623.400 747.600 624.300 757.950 ;
        RECT 645.000 754.200 645.900 757.950 ;
        RECT 647.100 756.150 648.900 757.950 ;
        RECT 653.100 756.150 654.900 757.950 ;
        RECT 671.100 756.150 672.900 757.950 ;
        RECT 645.000 753.000 648.300 754.200 ;
        RECT 620.100 744.000 621.900 747.600 ;
        RECT 623.100 744.600 624.900 747.600 ;
        RECT 626.100 744.000 627.900 747.600 ;
        RECT 646.500 744.600 648.300 753.000 ;
        RECT 653.100 744.000 654.900 753.600 ;
        RECT 674.700 752.700 675.900 757.950 ;
        RECT 676.950 756.150 678.750 757.950 ;
        RECT 671.700 751.800 675.900 752.700 ;
        RECT 671.700 744.600 673.500 751.800 ;
        RECT 676.800 744.000 678.600 750.600 ;
        RECT 698.400 747.600 699.300 757.950 ;
        RECT 707.550 757.050 708.450 760.950 ;
        RECT 722.100 760.050 723.300 767.400 ;
        RECT 740.250 760.050 742.050 761.850 ;
        RECT 743.400 760.050 744.300 767.400 ;
        RECT 748.950 762.450 753.000 763.050 ;
        RECT 746.100 760.050 747.900 761.850 ;
        RECT 748.950 760.950 753.450 762.450 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 703.950 755.550 708.450 757.050 ;
        RECT 719.100 756.150 720.900 757.950 ;
        RECT 703.950 754.950 708.000 755.550 ;
        RECT 722.100 750.600 723.300 757.950 ;
        RECT 695.100 744.000 696.900 747.600 ;
        RECT 698.100 744.600 699.900 747.600 ;
        RECT 701.100 744.000 702.900 747.600 ;
        RECT 719.100 744.000 720.900 750.600 ;
        RECT 722.100 744.600 723.900 750.600 ;
        RECT 743.400 747.600 744.300 757.950 ;
        RECT 752.550 756.450 753.450 760.950 ;
        RECT 764.700 760.050 765.900 767.400 ;
        RECT 785.100 760.050 786.900 761.850 ;
        RECT 788.700 760.050 789.600 767.400 ;
        RECT 790.950 760.050 792.750 761.850 ;
        RECT 812.100 760.050 813.300 773.400 ;
        RECT 833.100 767.400 834.900 779.400 ;
        RECT 836.100 768.300 837.900 779.400 ;
        RECT 839.100 769.200 840.900 780.000 ;
        RECT 842.100 768.300 843.900 779.400 ;
        RECT 836.100 767.400 843.900 768.300 ;
        RECT 860.100 767.400 861.900 780.000 ;
        RECT 863.100 767.400 864.900 779.400 ;
        RECT 881.100 773.400 882.900 780.000 ;
        RECT 884.100 773.400 885.900 779.400 ;
        RECT 865.950 768.450 868.050 769.050 ;
        RECT 874.950 768.450 877.050 769.050 ;
        RECT 865.950 767.550 877.050 768.450 ;
        RECT 833.400 760.050 834.300 767.400 ;
        RECT 847.950 762.450 850.050 763.050 ;
        RECT 856.950 762.450 859.050 763.050 ;
        RECT 838.950 760.050 840.750 761.850 ;
        RECT 847.950 761.550 859.050 762.450 ;
        RECT 847.950 760.950 850.050 761.550 ;
        RECT 856.950 760.950 859.050 761.550 ;
        RECT 863.100 760.050 864.300 767.400 ;
        RECT 865.950 766.950 868.050 767.550 ;
        RECT 874.950 766.950 877.050 767.550 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 881.100 757.950 883.200 760.050 ;
        RECT 760.950 756.450 763.050 757.050 ;
        RECT 752.550 755.550 763.050 756.450 ;
        RECT 760.950 754.950 763.050 755.550 ;
        RECT 764.700 750.600 765.900 757.950 ;
        RECT 767.100 756.150 768.900 757.950 ;
        RECT 740.100 744.000 741.900 747.600 ;
        RECT 743.100 744.600 744.900 747.600 ;
        RECT 746.100 744.000 747.900 747.600 ;
        RECT 764.100 744.600 765.900 750.600 ;
        RECT 767.100 744.000 768.900 750.600 ;
        RECT 788.700 747.600 789.600 757.950 ;
        RECT 809.250 756.150 811.050 757.950 ;
        RECT 812.100 752.700 813.300 757.950 ;
        RECT 815.100 756.150 816.900 757.950 ;
        RECT 817.950 756.450 820.050 757.050 ;
        RECT 826.950 756.450 829.050 757.050 ;
        RECT 817.950 755.550 829.050 756.450 ;
        RECT 817.950 754.950 820.050 755.550 ;
        RECT 826.950 754.950 829.050 755.550 ;
        RECT 812.100 751.800 816.300 752.700 ;
        RECT 785.100 744.000 786.900 747.600 ;
        RECT 788.100 744.600 789.900 747.600 ;
        RECT 791.100 744.000 792.900 747.600 ;
        RECT 809.400 744.000 811.200 750.600 ;
        RECT 814.500 744.600 816.300 751.800 ;
        RECT 833.400 750.600 834.300 757.950 ;
        RECT 835.950 756.150 837.750 757.950 ;
        RECT 842.100 756.150 843.900 757.950 ;
        RECT 860.100 756.150 861.900 757.950 ;
        RECT 863.100 750.600 864.300 757.950 ;
        RECT 881.250 756.150 883.050 757.950 ;
        RECT 884.100 753.300 885.000 773.400 ;
        RECT 887.100 768.000 888.900 780.000 ;
        RECT 890.100 767.400 891.900 779.400 ;
        RECT 908.100 767.400 909.900 780.000 ;
        RECT 911.100 767.400 912.900 779.400 ;
        RECT 886.200 760.050 888.000 761.850 ;
        RECT 890.400 760.050 891.300 767.400 ;
        RECT 911.100 760.050 912.300 767.400 ;
        RECT 919.950 766.950 922.050 769.050 ;
        RECT 929.100 767.400 930.900 779.400 ;
        RECT 932.100 768.300 933.900 779.400 ;
        RECT 935.100 769.200 936.900 780.000 ;
        RECT 938.100 768.300 939.900 779.400 ;
        RECT 932.100 767.400 939.900 768.300 ;
        RECT 953.100 767.400 954.900 780.000 ;
        RECT 958.200 768.600 960.000 779.400 ;
        RECT 977.100 773.400 978.900 780.000 ;
        RECT 980.100 773.400 981.900 779.400 ;
        RECT 983.100 773.400 984.900 780.000 ;
        RECT 956.400 767.400 960.000 768.600 ;
        RECT 886.500 757.950 888.600 760.050 ;
        RECT 889.800 757.950 891.900 760.050 ;
        RECT 907.950 757.950 910.050 760.050 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 881.100 752.400 889.500 753.300 ;
        RECT 833.400 749.400 838.500 750.600 ;
        RECT 833.700 744.000 835.500 747.600 ;
        RECT 836.700 744.600 838.500 749.400 ;
        RECT 841.200 744.000 843.000 750.600 ;
        RECT 860.100 744.000 861.900 750.600 ;
        RECT 863.100 744.600 864.900 750.600 ;
        RECT 881.100 744.600 882.900 752.400 ;
        RECT 887.700 751.500 889.500 752.400 ;
        RECT 890.400 750.600 891.300 757.950 ;
        RECT 908.100 756.150 909.900 757.950 ;
        RECT 911.100 750.600 912.300 757.950 ;
        RECT 920.550 751.050 921.450 766.950 ;
        RECT 929.400 760.050 930.300 767.400 ;
        RECT 934.950 760.050 936.750 761.850 ;
        RECT 953.250 760.050 955.050 761.850 ;
        RECT 956.400 760.050 957.300 767.400 ;
        RECT 967.950 765.450 970.050 766.050 ;
        RECT 976.950 765.450 979.050 766.050 ;
        RECT 967.950 764.550 979.050 765.450 ;
        RECT 967.950 763.950 970.050 764.550 ;
        RECT 976.950 763.950 979.050 764.550 ;
        RECT 961.950 762.450 964.050 763.050 ;
        RECT 959.100 760.050 960.900 761.850 ;
        RECT 961.950 761.550 972.450 762.450 ;
        RECT 961.950 760.950 964.050 761.550 ;
        RECT 928.950 757.950 931.050 760.050 ;
        RECT 931.950 757.950 934.050 760.050 ;
        RECT 934.950 757.950 937.050 760.050 ;
        RECT 937.950 757.950 940.050 760.050 ;
        RECT 952.950 757.950 955.050 760.050 ;
        RECT 955.950 757.950 958.050 760.050 ;
        RECT 958.950 757.950 961.050 760.050 ;
        RECT 885.600 744.000 887.400 750.600 ;
        RECT 888.600 748.800 891.300 750.600 ;
        RECT 888.600 744.600 890.400 748.800 ;
        RECT 908.100 744.000 909.900 750.600 ;
        RECT 911.100 744.600 912.900 750.600 ;
        RECT 919.950 748.950 922.050 751.050 ;
        RECT 929.400 750.600 930.300 757.950 ;
        RECT 931.950 756.150 933.750 757.950 ;
        RECT 938.100 756.150 939.900 757.950 ;
        RECT 929.400 749.400 934.500 750.600 ;
        RECT 929.700 744.000 931.500 747.600 ;
        RECT 932.700 744.600 934.500 749.400 ;
        RECT 937.200 744.000 939.000 750.600 ;
        RECT 956.400 747.600 957.300 757.950 ;
        RECT 961.950 756.450 964.050 757.050 ;
        RECT 967.950 756.450 970.050 760.050 ;
        RECT 961.950 756.000 970.050 756.450 ;
        RECT 971.550 757.050 972.450 761.550 ;
        RECT 980.100 760.050 981.300 773.400 ;
        RECT 1001.400 767.400 1003.200 780.000 ;
        RECT 1006.500 768.900 1008.300 779.400 ;
        RECT 1009.500 773.400 1011.300 780.000 ;
        RECT 1009.200 770.100 1011.000 771.900 ;
        RECT 1029.600 768.900 1031.400 779.400 ;
        RECT 1006.500 767.400 1008.900 768.900 ;
        RECT 997.950 762.450 1000.050 763.050 ;
        RECT 989.550 761.550 1000.050 762.450 ;
        RECT 976.950 757.950 979.050 760.050 ;
        RECT 979.950 757.950 982.050 760.050 ;
        RECT 982.950 757.950 985.050 760.050 ;
        RECT 961.950 755.550 969.450 756.000 ;
        RECT 971.550 755.550 976.050 757.050 ;
        RECT 977.250 756.150 979.050 757.950 ;
        RECT 961.950 754.950 964.050 755.550 ;
        RECT 972.000 754.950 976.050 755.550 ;
        RECT 980.100 752.700 981.300 757.950 ;
        RECT 983.100 756.150 984.900 757.950 ;
        RECT 989.550 757.050 990.450 761.550 ;
        RECT 997.950 760.950 1000.050 761.550 ;
        RECT 1001.100 760.050 1002.900 761.850 ;
        RECT 1007.700 760.050 1008.900 767.400 ;
        RECT 1029.000 767.400 1031.400 768.900 ;
        RECT 1032.600 767.400 1034.400 780.000 ;
        RECT 1037.100 767.400 1038.900 779.400 ;
        RECT 1018.950 763.950 1021.050 766.050 ;
        RECT 1000.950 757.950 1003.050 760.050 ;
        RECT 1003.950 757.950 1006.050 760.050 ;
        RECT 1006.950 757.950 1009.050 760.050 ;
        RECT 1009.950 757.950 1012.050 760.050 ;
        RECT 985.950 755.550 990.450 757.050 ;
        RECT 1004.100 756.150 1005.900 757.950 ;
        RECT 985.950 754.950 990.000 755.550 ;
        RECT 1007.700 753.600 1008.900 757.950 ;
        RECT 1010.100 756.150 1011.900 757.950 ;
        RECT 1007.700 752.700 1011.300 753.600 ;
        RECT 980.100 751.800 984.300 752.700 ;
        RECT 953.100 744.000 954.900 747.600 ;
        RECT 956.100 744.600 957.900 747.600 ;
        RECT 959.100 744.000 960.900 747.600 ;
        RECT 977.400 744.000 979.200 750.600 ;
        RECT 982.500 744.600 984.300 751.800 ;
        RECT 1001.100 749.700 1008.900 751.050 ;
        RECT 1001.100 744.600 1002.900 749.700 ;
        RECT 1004.100 744.000 1005.900 748.800 ;
        RECT 1007.100 744.600 1008.900 749.700 ;
        RECT 1010.100 750.600 1011.300 752.700 ;
        RECT 1019.550 751.050 1020.450 763.950 ;
        RECT 1029.000 760.050 1030.200 767.400 ;
        RECT 1037.700 765.900 1038.900 767.400 ;
        RECT 1031.100 764.700 1038.900 765.900 ;
        RECT 1031.100 764.100 1032.900 764.700 ;
        RECT 1028.100 757.950 1030.200 760.050 ;
        RECT 1019.550 750.900 1023.000 751.050 ;
        RECT 1010.100 744.600 1011.900 750.600 ;
        RECT 1019.550 749.550 1024.050 750.900 ;
        RECT 1020.000 748.950 1024.050 749.550 ;
        RECT 1021.950 748.800 1024.050 748.950 ;
        RECT 1028.100 750.600 1029.000 757.950 ;
        RECT 1031.400 753.600 1032.300 764.100 ;
        RECT 1033.200 760.050 1035.000 761.850 ;
        RECT 1033.500 757.950 1035.600 760.050 ;
        RECT 1036.800 757.950 1038.900 760.050 ;
        RECT 1036.800 756.150 1038.600 757.950 ;
        RECT 1030.200 752.700 1032.300 753.600 ;
        RECT 1030.200 751.800 1035.600 752.700 ;
        RECT 1028.100 744.600 1029.900 750.600 ;
        RECT 1031.100 744.000 1032.900 750.000 ;
        RECT 1034.700 747.600 1035.600 751.800 ;
        RECT 1034.100 744.600 1035.900 747.600 ;
        RECT 1037.100 744.600 1038.900 747.600 ;
        RECT 1037.700 744.000 1038.900 744.600 ;
        RECT 17.100 734.400 18.900 740.400 ;
        RECT 20.100 734.400 21.900 741.000 ;
        RECT 23.100 737.400 24.900 740.400 ;
        RECT 17.100 727.050 18.300 734.400 ;
        RECT 23.700 733.500 24.900 737.400 ;
        RECT 19.200 732.600 24.900 733.500 ;
        RECT 41.100 737.400 42.900 740.400 ;
        RECT 41.100 733.500 42.300 737.400 ;
        RECT 44.100 734.400 45.900 741.000 ;
        RECT 47.100 734.400 48.900 740.400 ;
        RECT 41.100 732.600 46.800 733.500 ;
        RECT 19.200 731.700 21.000 732.600 ;
        RECT 17.100 724.950 19.200 727.050 ;
        RECT 17.100 717.600 18.300 724.950 ;
        RECT 20.100 720.300 21.000 731.700 ;
        RECT 45.000 731.700 46.800 732.600 ;
        RECT 22.500 724.950 24.600 727.050 ;
        RECT 22.800 723.150 24.600 724.950 ;
        RECT 41.400 724.950 43.500 727.050 ;
        RECT 41.400 723.150 43.200 724.950 ;
        RECT 19.200 719.400 21.000 720.300 ;
        RECT 45.000 720.300 45.900 731.700 ;
        RECT 47.700 727.050 48.900 734.400 ;
        RECT 65.100 737.400 66.900 740.400 ;
        RECT 65.100 733.500 66.300 737.400 ;
        RECT 68.100 734.400 69.900 741.000 ;
        RECT 71.100 734.400 72.900 740.400 ;
        RECT 65.100 732.600 70.800 733.500 ;
        RECT 69.000 731.700 70.800 732.600 ;
        RECT 46.800 724.950 48.900 727.050 ;
        RECT 45.000 719.400 46.800 720.300 ;
        RECT 19.200 718.500 24.900 719.400 ;
        RECT 17.100 705.600 18.900 717.600 ;
        RECT 20.100 705.000 21.900 715.800 ;
        RECT 23.700 711.600 24.900 718.500 ;
        RECT 23.100 705.600 24.900 711.600 ;
        RECT 41.100 718.500 46.800 719.400 ;
        RECT 41.100 711.600 42.300 718.500 ;
        RECT 47.700 717.600 48.900 724.950 ;
        RECT 65.400 724.950 67.500 727.050 ;
        RECT 65.400 723.150 67.200 724.950 ;
        RECT 69.000 720.300 69.900 731.700 ;
        RECT 71.700 727.050 72.900 734.400 ;
        RECT 89.700 733.200 91.500 740.400 ;
        RECT 94.800 734.400 96.600 741.000 ;
        RECT 113.100 737.400 114.900 740.400 ;
        RECT 116.100 737.400 117.900 741.000 ;
        RECT 134.100 737.400 135.900 741.000 ;
        RECT 137.100 737.400 138.900 740.400 ;
        RECT 140.100 737.400 141.900 741.000 ;
        RECT 89.700 732.300 93.900 733.200 ;
        RECT 89.100 727.050 90.900 728.850 ;
        RECT 92.700 727.050 93.900 732.300 ;
        RECT 94.950 727.050 96.750 728.850 ;
        RECT 113.700 727.050 114.900 737.400 ;
        RECT 115.950 732.450 118.050 733.050 ;
        RECT 133.950 732.450 136.050 733.050 ;
        RECT 115.950 731.550 136.050 732.450 ;
        RECT 115.950 730.950 118.050 731.550 ;
        RECT 133.950 730.950 136.050 731.550 ;
        RECT 137.400 727.050 138.300 737.400 ;
        RECT 158.100 735.300 159.900 740.400 ;
        RECT 161.100 736.200 162.900 741.000 ;
        RECT 164.100 735.300 165.900 740.400 ;
        RECT 158.100 733.950 165.900 735.300 ;
        RECT 167.100 734.400 168.900 740.400 ;
        RECT 170.700 734.400 172.500 740.400 ;
        RECT 176.100 734.400 177.900 741.000 ;
        RECT 181.500 734.400 183.300 740.400 ;
        RECT 185.700 737.400 187.500 740.400 ;
        RECT 188.700 737.400 190.500 740.400 ;
        RECT 191.700 737.400 193.500 740.400 ;
        RECT 194.700 737.400 196.500 741.000 ;
        RECT 185.700 735.300 187.800 737.400 ;
        RECT 188.700 735.300 190.800 737.400 ;
        RECT 191.700 735.300 193.800 737.400 ;
        RECT 199.200 736.500 201.000 740.400 ;
        RECT 202.200 737.400 204.000 741.000 ;
        RECT 205.200 737.400 207.000 740.400 ;
        RECT 208.200 737.400 210.000 740.400 ;
        RECT 211.200 737.400 213.000 740.400 ;
        RECT 214.200 737.400 216.000 740.400 ;
        RECT 195.600 735.600 197.400 736.500 ;
        RECT 194.700 734.400 197.400 735.600 ;
        RECT 199.200 734.400 201.900 736.500 ;
        RECT 205.200 735.300 207.300 737.400 ;
        RECT 208.200 735.300 210.300 737.400 ;
        RECT 211.200 735.300 213.300 737.400 ;
        RECT 214.200 735.300 216.300 737.400 ;
        RECT 218.400 735.600 220.200 740.400 ;
        RECT 218.400 734.400 222.600 735.600 ;
        RECT 223.500 734.400 225.300 741.000 ;
        RECT 228.900 734.400 230.700 740.400 ;
        RECT 167.100 732.300 168.300 734.400 ;
        RECT 164.700 731.400 168.300 732.300 ;
        RECT 161.100 727.050 162.900 728.850 ;
        RECT 164.700 727.050 165.900 731.400 ;
        RECT 170.700 730.800 171.900 734.400 ;
        RECT 181.800 733.500 183.300 734.400 ;
        RECT 190.800 733.800 192.600 734.400 ;
        RECT 194.700 733.800 195.600 734.400 ;
        RECT 174.900 732.300 183.300 733.500 ;
        RECT 188.400 732.600 195.600 733.800 ;
        RECT 210.300 732.600 216.900 734.400 ;
        RECT 174.900 731.700 176.700 732.300 ;
        RECT 185.400 730.800 187.500 731.700 ;
        RECT 170.700 729.600 187.500 730.800 ;
        RECT 188.400 729.600 189.300 732.600 ;
        RECT 193.800 729.900 195.600 730.800 ;
        RECT 203.100 730.500 204.900 732.300 ;
        RECT 221.100 731.100 222.600 734.400 ;
        RECT 196.800 729.900 198.900 730.050 ;
        RECT 167.100 727.050 168.900 728.850 ;
        RECT 70.800 724.950 72.900 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 91.950 724.950 94.050 727.050 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 115.950 724.950 118.050 727.050 ;
        RECT 133.950 724.950 136.050 727.050 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 157.950 724.950 160.050 727.050 ;
        RECT 160.950 724.950 163.050 727.050 ;
        RECT 163.950 724.950 166.050 727.050 ;
        RECT 166.950 724.950 169.050 727.050 ;
        RECT 69.000 719.400 70.800 720.300 ;
        RECT 41.100 705.600 42.900 711.600 ;
        RECT 44.100 705.000 45.900 715.800 ;
        RECT 47.100 705.600 48.900 717.600 ;
        RECT 65.100 718.500 70.800 719.400 ;
        RECT 65.100 711.600 66.300 718.500 ;
        RECT 71.700 717.600 72.900 724.950 ;
        RECT 65.100 705.600 66.900 711.600 ;
        RECT 68.100 705.000 69.900 715.800 ;
        RECT 71.100 705.600 72.900 717.600 ;
        RECT 92.700 711.600 93.900 724.950 ;
        RECT 113.700 711.600 114.900 724.950 ;
        RECT 116.100 723.150 117.900 724.950 ;
        RECT 134.250 723.150 136.050 724.950 ;
        RECT 137.400 717.600 138.300 724.950 ;
        RECT 140.100 723.150 141.900 724.950 ;
        RECT 158.100 723.150 159.900 724.950 ;
        RECT 164.700 717.600 165.900 724.950 ;
        RECT 89.100 705.000 90.900 711.600 ;
        RECT 92.100 705.600 93.900 711.600 ;
        RECT 95.100 705.000 96.900 711.600 ;
        RECT 113.100 705.600 114.900 711.600 ;
        RECT 116.100 705.000 117.900 711.600 ;
        RECT 134.100 705.000 135.900 717.600 ;
        RECT 137.400 716.400 141.000 717.600 ;
        RECT 139.200 705.600 141.000 716.400 ;
        RECT 158.400 705.000 160.200 717.600 ;
        RECT 163.500 716.100 165.900 717.600 ;
        RECT 163.500 705.600 165.300 716.100 ;
        RECT 166.200 713.100 168.000 714.900 ;
        RECT 170.700 713.400 171.900 729.600 ;
        RECT 188.400 727.800 190.200 729.600 ;
        RECT 193.800 729.000 198.900 729.900 ;
        RECT 196.800 727.950 198.900 729.000 ;
        RECT 203.100 729.900 205.200 730.500 ;
        RECT 203.100 728.400 220.200 729.900 ;
        RECT 221.100 729.300 228.900 731.100 ;
        RECT 218.700 726.900 225.300 728.400 ;
        RECT 173.100 725.700 217.500 726.900 ;
        RECT 173.100 724.050 174.900 725.700 ;
        RECT 172.800 721.950 174.900 724.050 ;
        RECT 178.800 723.750 180.900 724.050 ;
        RECT 191.400 723.900 193.200 724.500 ;
        RECT 200.400 723.900 213.900 724.800 ;
        RECT 178.800 721.950 182.700 723.750 ;
        RECT 191.400 722.700 202.500 723.900 ;
        RECT 180.900 721.200 182.700 721.950 ;
        RECT 200.400 721.800 202.500 722.700 ;
        RECT 204.000 721.200 207.900 723.000 ;
        RECT 213.000 722.700 213.900 723.900 ;
        RECT 180.900 720.300 194.400 721.200 ;
        RECT 205.800 720.900 207.900 721.200 ;
        RECT 212.100 720.900 213.900 722.700 ;
        RECT 216.600 724.200 217.500 725.700 ;
        RECT 216.600 722.400 221.700 724.200 ;
        RECT 223.800 724.050 225.300 726.900 ;
        RECT 223.800 721.950 225.900 724.050 ;
        RECT 193.200 719.700 194.400 720.300 ;
        RECT 227.100 719.700 228.900 720.300 ;
        RECT 188.400 718.500 190.500 718.800 ;
        RECT 193.200 718.500 228.900 719.700 ;
        RECT 178.500 717.300 190.500 718.500 ;
        RECT 229.800 717.600 230.700 734.400 ;
        RECT 178.500 716.700 180.300 717.300 ;
        RECT 188.400 716.700 190.500 717.300 ;
        RECT 193.200 716.400 210.900 717.600 ;
        RECT 175.200 715.800 177.000 716.100 ;
        RECT 193.200 715.800 194.400 716.400 ;
        RECT 175.200 714.600 194.400 715.800 ;
        RECT 208.800 715.500 210.900 716.400 ;
        RECT 214.200 716.700 230.700 717.600 ;
        RECT 214.200 715.500 216.300 716.700 ;
        RECT 175.200 714.300 177.000 714.600 ;
        RECT 170.700 712.500 174.300 713.400 ;
        RECT 173.400 711.600 174.300 712.500 ;
        RECT 166.500 705.000 168.300 711.600 ;
        RECT 170.700 705.000 172.500 711.600 ;
        RECT 173.400 710.700 175.500 711.600 ;
        RECT 173.700 705.600 175.500 710.700 ;
        RECT 176.700 705.000 178.500 711.600 ;
        RECT 179.700 705.600 181.500 714.600 ;
        RECT 191.700 711.600 193.800 713.700 ;
        RECT 199.200 713.100 202.500 715.200 ;
        RECT 182.700 705.000 184.500 711.600 ;
        RECT 186.300 708.600 188.400 710.700 ;
        RECT 189.300 708.600 191.400 710.700 ;
        RECT 186.300 705.600 188.100 708.600 ;
        RECT 189.300 705.600 191.100 708.600 ;
        RECT 192.300 705.600 194.100 711.600 ;
        RECT 195.300 705.000 197.100 711.600 ;
        RECT 199.200 705.600 201.000 713.100 ;
        RECT 205.200 711.600 207.900 715.500 ;
        RECT 220.200 714.600 225.900 715.800 ;
        RECT 217.500 713.700 219.300 714.300 ;
        RECT 211.200 712.500 219.300 713.700 ;
        RECT 211.200 711.600 213.300 712.500 ;
        RECT 220.200 711.600 221.400 714.600 ;
        RECT 224.100 714.000 225.900 714.600 ;
        RECT 229.800 713.400 230.700 716.700 ;
        RECT 226.800 712.500 230.700 713.400 ;
        RECT 232.500 737.400 234.300 740.400 ;
        RECT 235.500 737.400 237.300 741.000 ;
        RECT 232.500 724.050 234.000 737.400 ;
        RECT 255.000 734.400 256.800 741.000 ;
        RECT 259.500 735.600 261.300 740.400 ;
        RECT 262.500 737.400 264.300 741.000 ;
        RECT 281.100 737.400 282.900 741.000 ;
        RECT 284.100 737.400 285.900 740.400 ;
        RECT 259.500 734.400 264.600 735.600 ;
        RECT 241.950 732.450 244.050 733.050 ;
        RECT 259.950 732.450 262.050 733.050 ;
        RECT 241.950 731.550 262.050 732.450 ;
        RECT 241.950 730.950 244.050 731.550 ;
        RECT 259.950 730.950 262.050 731.550 ;
        RECT 254.100 727.050 255.900 728.850 ;
        RECT 260.250 727.050 262.050 728.850 ;
        RECT 263.700 727.050 264.600 734.400 ;
        RECT 284.100 727.050 285.300 737.400 ;
        RECT 302.400 734.400 304.200 741.000 ;
        RECT 307.500 733.200 309.300 740.400 ;
        RECT 326.100 737.400 327.900 741.000 ;
        RECT 329.100 737.400 330.900 740.400 ;
        RECT 305.100 732.300 309.300 733.200 ;
        RECT 316.950 732.450 319.050 733.050 ;
        RECT 325.950 732.450 328.050 733.050 ;
        RECT 302.250 727.050 304.050 728.850 ;
        RECT 305.100 727.050 306.300 732.300 ;
        RECT 316.950 731.550 328.050 732.450 ;
        RECT 316.950 730.950 319.050 731.550 ;
        RECT 325.950 730.950 328.050 731.550 ;
        RECT 308.100 727.050 309.900 728.850 ;
        RECT 329.100 727.050 330.300 737.400 ;
        RECT 347.100 735.300 348.900 740.400 ;
        RECT 350.100 736.200 351.900 741.000 ;
        RECT 353.100 735.300 354.900 740.400 ;
        RECT 347.100 733.950 354.900 735.300 ;
        RECT 356.100 734.400 357.900 740.400 ;
        RECT 374.400 734.400 376.200 741.000 ;
        RECT 356.100 732.300 357.300 734.400 ;
        RECT 379.500 733.200 381.300 740.400 ;
        RECT 398.100 737.400 399.900 740.400 ;
        RECT 401.100 737.400 402.900 741.000 ;
        RECT 353.700 731.400 357.300 732.300 ;
        RECT 377.100 732.300 381.300 733.200 ;
        RECT 350.100 727.050 351.900 728.850 ;
        RECT 353.700 727.050 354.900 731.400 ;
        RECT 356.100 727.050 357.900 728.850 ;
        RECT 374.250 727.050 376.050 728.850 ;
        RECT 377.100 727.050 378.300 732.300 ;
        RECT 382.950 729.450 385.050 730.050 ;
        RECT 391.950 729.450 394.050 730.050 ;
        RECT 380.100 727.050 381.900 728.850 ;
        RECT 382.950 728.550 394.050 729.450 ;
        RECT 382.950 727.950 385.050 728.550 ;
        RECT 391.950 727.950 394.050 728.550 ;
        RECT 398.700 727.050 399.900 737.400 ;
        RECT 419.400 734.400 421.200 741.000 ;
        RECT 424.500 733.200 426.300 740.400 ;
        RECT 443.100 734.400 444.900 741.000 ;
        RECT 446.100 734.400 447.900 740.400 ;
        RECT 422.100 732.300 426.300 733.200 ;
        RECT 419.250 727.050 421.050 728.850 ;
        RECT 422.100 727.050 423.300 732.300 ;
        RECT 425.100 727.050 426.900 728.850 ;
        RECT 443.100 727.050 444.900 728.850 ;
        RECT 446.100 727.050 447.300 734.400 ;
        RECT 464.100 731.400 465.900 741.000 ;
        RECT 470.700 732.000 472.500 740.400 ;
        RECT 491.400 734.400 493.200 741.000 ;
        RECT 496.500 733.200 498.300 740.400 ;
        RECT 515.100 737.400 516.900 741.000 ;
        RECT 518.100 737.400 519.900 740.400 ;
        RECT 521.100 737.400 522.900 741.000 ;
        RECT 494.100 732.300 498.300 733.200 ;
        RECT 470.700 730.800 474.000 732.000 ;
        RECT 464.100 727.050 465.900 728.850 ;
        RECT 470.100 727.050 471.900 728.850 ;
        RECT 473.100 727.050 474.000 730.800 ;
        RECT 491.250 727.050 493.050 728.850 ;
        RECT 494.100 727.050 495.300 732.300 ;
        RECT 497.100 727.050 498.900 728.850 ;
        RECT 518.400 727.050 519.300 737.400 ;
        RECT 539.100 735.300 540.900 740.400 ;
        RECT 542.100 736.200 543.900 741.000 ;
        RECT 545.100 735.300 546.900 740.400 ;
        RECT 539.100 733.950 546.900 735.300 ;
        RECT 548.100 734.400 549.900 740.400 ;
        RECT 566.100 737.400 567.900 741.000 ;
        RECT 569.100 737.400 570.900 740.400 ;
        RECT 572.100 737.400 573.900 741.000 ;
        RECT 548.100 732.300 549.300 734.400 ;
        RECT 545.700 731.400 549.300 732.300 ;
        RECT 529.950 729.450 532.050 730.050 ;
        RECT 535.950 729.450 538.050 730.050 ;
        RECT 529.950 728.550 538.050 729.450 ;
        RECT 529.950 727.950 532.050 728.550 ;
        RECT 535.950 727.950 538.050 728.550 ;
        RECT 542.100 727.050 543.900 728.850 ;
        RECT 545.700 727.050 546.900 731.400 ;
        RECT 548.100 727.050 549.900 728.850 ;
        RECT 569.400 727.050 570.300 737.400 ;
        RECT 590.400 734.400 592.200 741.000 ;
        RECT 595.500 733.200 597.300 740.400 ;
        RECT 593.100 732.300 597.300 733.200 ;
        RECT 614.100 734.400 615.900 740.400 ;
        RECT 617.100 735.000 618.900 741.000 ;
        RECT 623.700 740.400 624.900 741.000 ;
        RECT 620.100 737.400 621.900 740.400 ;
        RECT 623.100 737.400 624.900 740.400 ;
        RECT 590.250 727.050 592.050 728.850 ;
        RECT 593.100 727.050 594.300 732.300 ;
        RECT 596.100 727.050 597.900 728.850 ;
        RECT 614.100 727.050 615.000 734.400 ;
        RECT 620.700 733.200 621.600 737.400 ;
        RECT 641.100 735.000 642.900 740.400 ;
        RECT 644.100 735.900 645.900 741.000 ;
        RECT 647.100 739.500 654.900 740.400 ;
        RECT 647.100 735.000 648.900 739.500 ;
        RECT 641.100 734.100 648.900 735.000 ;
        RECT 650.100 734.400 651.900 738.600 ;
        RECT 653.100 734.400 654.900 739.500 ;
        RECT 616.200 732.300 621.600 733.200 ;
        RECT 622.950 732.450 625.050 733.050 ;
        RECT 640.950 732.450 643.050 733.200 ;
        RECT 650.400 732.900 651.300 734.400 ;
        RECT 616.200 731.400 618.300 732.300 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 262.950 724.950 265.050 727.050 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 541.950 724.950 544.050 727.050 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 571.950 724.950 574.050 727.050 ;
        RECT 589.950 724.950 592.050 727.050 ;
        RECT 592.950 724.950 595.050 727.050 ;
        RECT 595.950 724.950 598.050 727.050 ;
        RECT 614.100 724.950 616.200 727.050 ;
        RECT 232.500 721.950 234.900 724.050 ;
        RECT 257.250 723.150 259.050 724.950 ;
        RECT 226.800 711.600 228.000 712.500 ;
        RECT 232.500 711.600 234.000 721.950 ;
        RECT 263.700 717.600 264.600 724.950 ;
        RECT 281.100 723.150 282.900 724.950 ;
        RECT 254.100 716.700 261.900 717.600 ;
        RECT 202.200 705.000 204.000 711.600 ;
        RECT 205.200 705.600 207.000 711.600 ;
        RECT 208.200 708.600 210.300 710.700 ;
        RECT 211.200 708.600 213.300 710.700 ;
        RECT 214.200 708.600 216.300 710.700 ;
        RECT 208.200 705.600 210.000 708.600 ;
        RECT 211.200 705.600 213.000 708.600 ;
        RECT 214.200 705.600 216.000 708.600 ;
        RECT 217.200 705.000 219.000 711.600 ;
        RECT 220.200 705.600 222.000 711.600 ;
        RECT 223.200 705.000 225.000 711.600 ;
        RECT 226.200 705.600 228.000 711.600 ;
        RECT 229.200 705.000 231.000 711.600 ;
        RECT 232.500 705.600 234.300 711.600 ;
        RECT 235.500 705.000 237.300 711.600 ;
        RECT 254.100 705.600 255.900 716.700 ;
        RECT 257.100 705.000 258.900 715.800 ;
        RECT 260.100 705.600 261.900 716.700 ;
        RECT 263.100 705.600 264.900 717.600 ;
        RECT 284.100 711.600 285.300 724.950 ;
        RECT 305.100 711.600 306.300 724.950 ;
        RECT 326.100 723.150 327.900 724.950 ;
        RECT 329.100 711.600 330.300 724.950 ;
        RECT 347.100 723.150 348.900 724.950 ;
        RECT 353.700 717.600 354.900 724.950 ;
        RECT 281.100 705.000 282.900 711.600 ;
        RECT 284.100 705.600 285.900 711.600 ;
        RECT 302.100 705.000 303.900 711.600 ;
        RECT 305.100 705.600 306.900 711.600 ;
        RECT 308.100 705.000 309.900 711.600 ;
        RECT 326.100 705.000 327.900 711.600 ;
        RECT 329.100 705.600 330.900 711.600 ;
        RECT 347.400 705.000 349.200 717.600 ;
        RECT 352.500 716.100 354.900 717.600 ;
        RECT 352.500 705.600 354.300 716.100 ;
        RECT 355.200 713.100 357.000 714.900 ;
        RECT 377.100 711.600 378.300 724.950 ;
        RECT 379.950 714.450 382.050 715.050 ;
        RECT 391.950 714.450 394.050 715.050 ;
        RECT 379.950 713.550 394.050 714.450 ;
        RECT 379.950 712.950 382.050 713.550 ;
        RECT 391.950 712.950 394.050 713.550 ;
        RECT 398.700 711.600 399.900 724.950 ;
        RECT 401.100 723.150 402.900 724.950 ;
        RECT 422.100 711.600 423.300 724.950 ;
        RECT 433.950 720.450 436.050 721.050 ;
        RECT 442.950 720.450 445.050 721.050 ;
        RECT 433.950 719.550 445.050 720.450 ;
        RECT 433.950 718.950 436.050 719.550 ;
        RECT 442.950 718.950 445.050 719.550 ;
        RECT 446.100 717.600 447.300 724.950 ;
        RECT 467.100 723.150 468.900 724.950 ;
        RECT 355.500 705.000 357.300 711.600 ;
        RECT 374.100 705.000 375.900 711.600 ;
        RECT 377.100 705.600 378.900 711.600 ;
        RECT 380.100 705.000 381.900 711.600 ;
        RECT 398.100 705.600 399.900 711.600 ;
        RECT 401.100 705.000 402.900 711.600 ;
        RECT 419.100 705.000 420.900 711.600 ;
        RECT 422.100 705.600 423.900 711.600 ;
        RECT 425.100 705.000 426.900 711.600 ;
        RECT 443.100 705.000 444.900 717.600 ;
        RECT 446.100 705.600 447.900 717.600 ;
        RECT 473.100 712.800 474.000 724.950 ;
        RECT 467.400 711.900 474.000 712.800 ;
        RECT 467.400 711.600 468.900 711.900 ;
        RECT 448.950 708.450 451.050 709.050 ;
        RECT 460.950 708.450 463.050 709.050 ;
        RECT 448.950 707.550 463.050 708.450 ;
        RECT 448.950 706.950 451.050 707.550 ;
        RECT 460.950 706.950 463.050 707.550 ;
        RECT 464.100 705.000 465.900 711.600 ;
        RECT 467.100 705.600 468.900 711.600 ;
        RECT 473.100 711.600 474.000 711.900 ;
        RECT 494.100 711.600 495.300 724.950 ;
        RECT 515.250 723.150 517.050 724.950 ;
        RECT 518.400 717.600 519.300 724.950 ;
        RECT 521.100 723.150 522.900 724.950 ;
        RECT 539.100 723.150 540.900 724.950 ;
        RECT 545.700 717.600 546.900 724.950 ;
        RECT 566.250 723.150 568.050 724.950 ;
        RECT 569.400 717.600 570.300 724.950 ;
        RECT 572.100 723.150 573.900 724.950 ;
        RECT 577.950 723.450 580.050 724.050 ;
        RECT 586.950 723.450 589.050 724.050 ;
        RECT 577.950 722.550 589.050 723.450 ;
        RECT 577.950 721.950 580.050 722.550 ;
        RECT 586.950 721.950 589.050 722.550 ;
        RECT 470.100 705.000 471.900 711.000 ;
        RECT 473.100 705.600 474.900 711.600 ;
        RECT 491.100 705.000 492.900 711.600 ;
        RECT 494.100 705.600 495.900 711.600 ;
        RECT 497.100 705.000 498.900 711.600 ;
        RECT 515.100 705.000 516.900 717.600 ;
        RECT 518.400 716.400 522.000 717.600 ;
        RECT 520.200 705.600 522.000 716.400 ;
        RECT 539.400 705.000 541.200 717.600 ;
        RECT 544.500 716.100 546.900 717.600 ;
        RECT 544.500 705.600 546.300 716.100 ;
        RECT 547.200 713.100 549.000 714.900 ;
        RECT 547.500 705.000 549.300 711.600 ;
        RECT 566.100 705.000 567.900 717.600 ;
        RECT 569.400 716.400 573.000 717.600 ;
        RECT 571.200 705.600 573.000 716.400 ;
        RECT 593.100 711.600 594.300 724.950 ;
        RECT 615.000 717.600 616.200 724.950 ;
        RECT 617.400 720.900 618.300 731.400 ;
        RECT 622.950 731.550 643.050 732.450 ;
        RECT 622.950 730.950 625.050 731.550 ;
        RECT 640.950 731.100 643.050 731.550 ;
        RECT 646.950 731.700 651.300 732.900 ;
        RECT 671.700 733.200 673.500 740.400 ;
        RECT 676.800 734.400 678.600 741.000 ;
        RECT 695.100 737.400 696.900 741.000 ;
        RECT 698.100 737.400 699.900 740.400 ;
        RECT 701.100 737.400 702.900 741.000 ;
        RECT 671.700 732.300 675.900 733.200 ;
        RECT 622.800 727.050 624.600 728.850 ;
        RECT 644.250 727.050 646.050 728.850 ;
        RECT 619.500 724.950 621.600 727.050 ;
        RECT 622.800 724.950 624.900 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 727.050 648.000 731.700 ;
        RECT 667.950 729.450 670.050 730.050 ;
        RECT 649.950 727.050 651.750 728.850 ;
        RECT 659.550 728.550 670.050 729.450 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 649.950 724.950 652.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 619.200 723.150 621.000 724.950 ;
        RECT 641.100 723.150 642.900 724.950 ;
        RECT 617.100 720.300 618.900 720.900 ;
        RECT 617.100 719.100 624.900 720.300 ;
        RECT 623.700 717.600 624.900 719.100 ;
        RECT 646.950 717.600 648.000 724.950 ;
        RECT 652.950 723.150 654.750 724.950 ;
        RECT 659.550 724.050 660.450 728.550 ;
        RECT 667.950 727.950 670.050 728.550 ;
        RECT 671.100 727.050 672.900 728.850 ;
        RECT 674.700 727.050 675.900 732.300 ;
        RECT 676.950 727.050 678.750 728.850 ;
        RECT 698.400 727.050 699.300 737.400 ;
        RECT 719.400 734.400 721.200 741.000 ;
        RECT 724.500 733.200 726.300 740.400 ;
        RECT 722.100 732.300 726.300 733.200 ;
        RECT 719.250 727.050 721.050 728.850 ;
        RECT 722.100 727.050 723.300 732.300 ;
        RECT 745.500 732.000 747.300 740.400 ;
        RECT 744.000 730.800 747.300 732.000 ;
        RECT 752.100 731.400 753.900 741.000 ;
        RECT 757.950 738.450 760.050 739.050 ;
        RECT 766.950 738.450 769.050 739.050 ;
        RECT 757.950 737.550 769.050 738.450 ;
        RECT 757.950 736.950 760.050 737.550 ;
        RECT 766.950 736.950 769.050 737.550 ;
        RECT 770.100 731.400 771.900 741.000 ;
        RECT 776.700 732.000 778.500 740.400 ;
        RECT 797.400 734.400 799.200 741.000 ;
        RECT 802.500 733.200 804.300 740.400 ;
        RECT 800.100 732.300 804.300 733.200 ;
        RECT 776.700 730.800 780.000 732.000 ;
        RECT 725.100 727.050 726.900 728.850 ;
        RECT 744.000 727.050 744.900 730.800 ;
        RECT 754.950 729.450 759.000 730.050 ;
        RECT 746.100 727.050 747.900 728.850 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 754.950 727.950 759.450 729.450 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 736.950 726.450 739.050 727.050 ;
        RECT 731.550 725.550 739.050 726.450 ;
        RECT 655.950 722.550 660.450 724.050 ;
        RECT 655.950 721.950 660.000 722.550 ;
        RECT 649.950 720.450 652.050 720.750 ;
        RECT 670.950 720.450 673.050 721.050 ;
        RECT 649.950 719.550 673.050 720.450 ;
        RECT 649.950 718.650 652.050 719.550 ;
        RECT 670.950 718.950 673.050 719.550 ;
        RECT 615.000 716.100 617.400 717.600 ;
        RECT 590.100 705.000 591.900 711.600 ;
        RECT 593.100 705.600 594.900 711.600 ;
        RECT 596.100 705.000 597.900 711.600 ;
        RECT 615.600 705.600 617.400 716.100 ;
        RECT 618.600 705.000 620.400 717.600 ;
        RECT 623.100 705.600 624.900 717.600 ;
        RECT 641.100 705.000 642.900 717.600 ;
        RECT 645.600 705.600 648.900 717.600 ;
        RECT 651.600 705.000 653.400 717.600 ;
        RECT 661.950 714.450 664.050 714.900 ;
        RECT 670.950 714.450 673.050 715.050 ;
        RECT 661.950 713.550 673.050 714.450 ;
        RECT 661.950 712.800 664.050 713.550 ;
        RECT 670.950 712.950 673.050 713.550 ;
        RECT 674.700 711.600 675.900 724.950 ;
        RECT 695.250 723.150 697.050 724.950 ;
        RECT 698.400 717.600 699.300 724.950 ;
        RECT 701.100 723.150 702.900 724.950 ;
        RECT 655.950 708.450 658.050 709.050 ;
        RECT 667.950 708.450 670.050 709.050 ;
        RECT 655.950 707.550 670.050 708.450 ;
        RECT 655.950 706.950 658.050 707.550 ;
        RECT 667.950 706.950 670.050 707.550 ;
        RECT 671.100 705.000 672.900 711.600 ;
        RECT 674.100 705.600 675.900 711.600 ;
        RECT 677.100 705.000 678.900 711.600 ;
        RECT 695.100 705.000 696.900 717.600 ;
        RECT 698.400 716.400 702.000 717.600 ;
        RECT 700.200 705.600 702.000 716.400 ;
        RECT 722.100 711.600 723.300 724.950 ;
        RECT 731.550 724.050 732.450 725.550 ;
        RECT 736.950 724.950 739.050 725.550 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 727.950 722.550 732.450 724.050 ;
        RECT 727.950 721.950 732.000 722.550 ;
        RECT 727.950 720.450 730.050 720.900 ;
        RECT 739.950 720.450 742.050 721.050 ;
        RECT 727.950 719.550 742.050 720.450 ;
        RECT 727.950 718.800 730.050 719.550 ;
        RECT 739.950 718.950 742.050 719.550 ;
        RECT 744.000 712.800 744.900 724.950 ;
        RECT 749.100 723.150 750.900 724.950 ;
        RECT 758.550 724.050 759.450 727.950 ;
        RECT 770.100 727.050 771.900 728.850 ;
        RECT 776.100 727.050 777.900 728.850 ;
        RECT 779.100 727.050 780.000 730.800 ;
        RECT 792.000 729.450 796.050 730.050 ;
        RECT 791.550 727.950 796.050 729.450 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 754.950 722.550 759.450 724.050 ;
        RECT 760.950 723.450 763.050 724.050 ;
        RECT 766.950 723.450 769.050 724.050 ;
        RECT 760.950 722.550 769.050 723.450 ;
        RECT 773.100 723.150 774.900 724.950 ;
        RECT 754.950 721.950 759.000 722.550 ;
        RECT 760.950 721.950 763.050 722.550 ;
        RECT 766.950 721.950 769.050 722.550 ;
        RECT 757.950 717.450 760.050 718.050 ;
        RECT 769.950 717.450 772.050 718.050 ;
        RECT 775.950 717.450 778.050 717.900 ;
        RECT 757.950 716.550 778.050 717.450 ;
        RECT 757.950 715.950 760.050 716.550 ;
        RECT 769.950 715.950 772.050 716.550 ;
        RECT 775.950 715.800 778.050 716.550 ;
        RECT 779.100 712.800 780.000 724.950 ;
        RECT 791.550 724.050 792.450 727.950 ;
        RECT 797.250 727.050 799.050 728.850 ;
        RECT 800.100 727.050 801.300 732.300 ;
        RECT 821.100 731.400 822.900 741.000 ;
        RECT 827.700 732.000 829.500 740.400 ;
        RECT 848.100 737.400 849.900 741.000 ;
        RECT 851.100 737.400 852.900 740.400 ;
        RECT 854.100 737.400 855.900 741.000 ;
        RECT 827.700 730.800 831.000 732.000 ;
        RECT 803.100 727.050 804.900 728.850 ;
        RECT 821.100 727.050 822.900 728.850 ;
        RECT 827.100 727.050 828.900 728.850 ;
        RECT 830.100 727.050 831.000 730.800 ;
        RECT 851.400 727.050 852.300 737.400 ;
        RECT 872.700 733.200 874.500 740.400 ;
        RECT 877.800 734.400 879.600 741.000 ;
        RECT 896.100 737.400 897.900 741.000 ;
        RECT 899.100 737.400 900.900 740.400 ;
        RECT 902.100 737.400 903.900 741.000 ;
        RECT 920.100 737.400 921.900 741.000 ;
        RECT 923.100 737.400 924.900 740.400 ;
        RECT 926.100 737.400 927.900 741.000 ;
        RECT 883.950 735.450 886.050 736.050 ;
        RECT 895.950 735.450 898.050 736.050 ;
        RECT 883.950 734.550 898.050 735.450 ;
        RECT 883.950 733.950 886.050 734.550 ;
        RECT 895.950 733.950 898.050 734.550 ;
        RECT 872.700 732.300 876.900 733.200 ;
        RECT 872.100 727.050 873.900 728.850 ;
        RECT 875.700 727.050 876.900 732.300 ;
        RECT 883.950 732.450 886.050 732.900 ;
        RECT 895.950 732.450 898.050 732.900 ;
        RECT 883.950 731.550 898.050 732.450 ;
        RECT 883.950 730.800 886.050 731.550 ;
        RECT 895.950 730.800 898.050 731.550 ;
        RECT 877.950 727.050 879.750 728.850 ;
        RECT 899.400 727.050 900.300 737.400 ;
        RECT 904.950 732.450 907.050 733.050 ;
        RECT 919.950 732.450 922.050 733.050 ;
        RECT 904.950 731.550 922.050 732.450 ;
        RECT 904.950 730.950 907.050 731.550 ;
        RECT 919.950 730.950 922.050 731.550 ;
        RECT 923.400 727.050 924.300 737.400 ;
        RECT 946.500 732.000 948.300 740.400 ;
        RECT 945.000 730.800 948.300 732.000 ;
        RECT 953.100 731.400 954.900 741.000 ;
        RECT 971.100 737.400 972.900 741.000 ;
        RECT 974.100 737.400 975.900 740.400 ;
        RECT 992.100 737.400 993.900 741.000 ;
        RECT 995.100 737.400 996.900 740.400 ;
        RECT 998.100 737.400 999.900 741.000 ;
        RECT 958.950 732.450 961.050 733.050 ;
        RECT 970.950 732.450 973.050 733.200 ;
        RECT 958.950 731.550 973.050 732.450 ;
        RECT 958.950 730.950 961.050 731.550 ;
        RECT 970.950 731.100 973.050 731.550 ;
        RECT 940.950 729.450 943.050 730.050 ;
        RECT 932.550 728.550 943.050 729.450 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 877.950 724.950 880.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 898.950 724.950 901.050 727.050 ;
        RECT 901.950 724.950 904.050 727.050 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 922.950 724.950 925.050 727.050 ;
        RECT 925.950 724.950 928.050 727.050 ;
        RECT 791.550 722.550 796.050 724.050 ;
        RECT 792.000 721.950 796.050 722.550 ;
        RECT 781.950 717.450 784.050 718.050 ;
        RECT 793.950 717.450 796.050 718.050 ;
        RECT 781.950 716.550 796.050 717.450 ;
        RECT 781.950 715.950 784.050 716.550 ;
        RECT 793.950 715.950 796.050 716.550 ;
        RECT 744.000 711.900 750.600 712.800 ;
        RECT 744.000 711.600 744.900 711.900 ;
        RECT 719.100 705.000 720.900 711.600 ;
        RECT 722.100 705.600 723.900 711.600 ;
        RECT 725.100 705.000 726.900 711.600 ;
        RECT 743.100 705.600 744.900 711.600 ;
        RECT 749.100 711.600 750.600 711.900 ;
        RECT 773.400 711.900 780.000 712.800 ;
        RECT 773.400 711.600 774.900 711.900 ;
        RECT 746.100 705.000 747.900 711.000 ;
        RECT 749.100 705.600 750.900 711.600 ;
        RECT 752.100 705.000 753.900 711.600 ;
        RECT 770.100 705.000 771.900 711.600 ;
        RECT 773.100 705.600 774.900 711.600 ;
        RECT 779.100 711.600 780.000 711.900 ;
        RECT 776.100 705.000 777.900 711.000 ;
        RECT 779.100 705.600 780.900 711.600 ;
        RECT 781.950 711.450 784.050 712.050 ;
        RECT 790.950 711.450 793.050 712.050 ;
        RECT 800.100 711.600 801.300 724.950 ;
        RECT 824.100 723.150 825.900 724.950 ;
        RECT 802.950 720.450 805.050 721.050 ;
        RECT 826.950 720.450 829.050 721.050 ;
        RECT 802.950 719.550 829.050 720.450 ;
        RECT 802.950 718.950 805.050 719.550 ;
        RECT 826.950 718.950 829.050 719.550 ;
        RECT 830.100 712.800 831.000 724.950 ;
        RECT 848.250 723.150 850.050 724.950 ;
        RECT 851.400 717.600 852.300 724.950 ;
        RECT 854.100 723.150 855.900 724.950 ;
        RECT 824.400 711.900 831.000 712.800 ;
        RECT 824.400 711.600 825.900 711.900 ;
        RECT 781.950 710.550 793.050 711.450 ;
        RECT 781.950 709.950 784.050 710.550 ;
        RECT 790.950 709.950 793.050 710.550 ;
        RECT 797.100 705.000 798.900 711.600 ;
        RECT 800.100 705.600 801.900 711.600 ;
        RECT 803.100 705.000 804.900 711.600 ;
        RECT 821.100 705.000 822.900 711.600 ;
        RECT 824.100 705.600 825.900 711.600 ;
        RECT 830.100 711.600 831.000 711.900 ;
        RECT 827.100 705.000 828.900 711.000 ;
        RECT 830.100 705.600 831.900 711.600 ;
        RECT 848.100 705.000 849.900 717.600 ;
        RECT 851.400 716.400 855.000 717.600 ;
        RECT 853.200 705.600 855.000 716.400 ;
        RECT 875.700 711.600 876.900 724.950 ;
        RECT 896.250 723.150 898.050 724.950 ;
        RECT 877.950 720.450 880.050 721.050 ;
        RECT 889.950 720.450 892.050 721.050 ;
        RECT 877.950 719.550 892.050 720.450 ;
        RECT 877.950 718.950 880.050 719.550 ;
        RECT 889.950 718.950 892.050 719.550 ;
        RECT 899.400 717.600 900.300 724.950 ;
        RECT 902.100 723.150 903.900 724.950 ;
        RECT 920.250 723.150 922.050 724.950 ;
        RECT 901.950 720.450 904.050 721.050 ;
        RECT 919.950 720.450 922.050 721.050 ;
        RECT 901.950 719.550 922.050 720.450 ;
        RECT 901.950 718.950 904.050 719.550 ;
        RECT 919.950 718.950 922.050 719.550 ;
        RECT 923.400 717.600 924.300 724.950 ;
        RECT 926.100 723.150 927.900 724.950 ;
        RECT 932.550 724.050 933.450 728.550 ;
        RECT 940.950 727.950 943.050 728.550 ;
        RECT 945.000 727.050 945.900 730.800 ;
        RECT 947.100 727.050 948.900 728.850 ;
        RECT 953.100 727.050 954.900 728.850 ;
        RECT 974.100 727.050 975.300 737.400 ;
        RECT 982.950 732.450 985.050 733.050 ;
        RECT 991.950 732.450 994.050 733.050 ;
        RECT 982.950 731.550 994.050 732.450 ;
        RECT 982.950 730.950 985.050 731.550 ;
        RECT 991.950 730.950 994.050 731.550 ;
        RECT 976.950 729.450 979.050 730.050 ;
        RECT 976.950 728.550 987.450 729.450 ;
        RECT 976.950 727.950 979.050 728.550 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 946.950 724.950 949.050 727.050 ;
        RECT 949.950 724.950 952.050 727.050 ;
        RECT 952.950 724.950 955.050 727.050 ;
        RECT 970.950 724.950 973.050 727.050 ;
        RECT 973.950 724.950 976.050 727.050 ;
        RECT 928.950 722.550 933.450 724.050 ;
        RECT 928.950 721.950 933.000 722.550 ;
        RECT 925.950 720.450 928.050 721.050 ;
        RECT 940.950 720.450 943.050 721.050 ;
        RECT 925.950 719.550 943.050 720.450 ;
        RECT 925.950 718.950 928.050 719.550 ;
        RECT 940.950 718.950 943.050 719.550 ;
        RECT 872.100 705.000 873.900 711.600 ;
        RECT 875.100 705.600 876.900 711.600 ;
        RECT 878.100 705.000 879.900 711.600 ;
        RECT 896.100 705.000 897.900 717.600 ;
        RECT 899.400 716.400 903.000 717.600 ;
        RECT 901.200 705.600 903.000 716.400 ;
        RECT 920.100 705.000 921.900 717.600 ;
        RECT 923.400 716.400 927.000 717.600 ;
        RECT 925.200 705.600 927.000 716.400 ;
        RECT 928.950 717.450 931.050 717.900 ;
        RECT 937.950 717.450 940.050 718.050 ;
        RECT 928.950 716.550 940.050 717.450 ;
        RECT 928.950 715.800 931.050 716.550 ;
        RECT 937.950 715.950 940.050 716.550 ;
        RECT 945.000 712.800 945.900 724.950 ;
        RECT 950.100 723.150 951.900 724.950 ;
        RECT 971.100 723.150 972.900 724.950 ;
        RECT 945.000 711.900 951.600 712.800 ;
        RECT 945.000 711.600 945.900 711.900 ;
        RECT 944.100 705.600 945.900 711.600 ;
        RECT 950.100 711.600 951.600 711.900 ;
        RECT 974.100 711.600 975.300 724.950 ;
        RECT 986.550 724.050 987.450 728.550 ;
        RECT 995.400 727.050 996.300 737.400 ;
        RECT 1016.700 733.200 1018.500 740.400 ;
        RECT 1021.800 734.400 1023.600 741.000 ;
        RECT 1016.700 732.300 1020.900 733.200 ;
        RECT 1016.100 727.050 1017.900 728.850 ;
        RECT 1019.700 727.050 1020.900 732.300 ;
        RECT 1024.950 729.450 1029.000 730.050 ;
        RECT 1021.950 727.050 1023.750 728.850 ;
        RECT 1024.950 727.950 1029.450 729.450 ;
        RECT 991.950 724.950 994.050 727.050 ;
        RECT 994.950 724.950 997.050 727.050 ;
        RECT 997.950 724.950 1000.050 727.050 ;
        RECT 1015.950 724.950 1018.050 727.050 ;
        RECT 1018.950 724.950 1021.050 727.050 ;
        RECT 1021.950 724.950 1024.050 727.050 ;
        RECT 1028.550 726.450 1029.450 727.950 ;
        RECT 1033.950 726.450 1036.050 726.900 ;
        RECT 1028.550 725.550 1036.050 726.450 ;
        RECT 986.550 722.550 991.050 724.050 ;
        RECT 992.250 723.150 994.050 724.950 ;
        RECT 987.000 721.950 991.050 722.550 ;
        RECT 995.400 717.600 996.300 724.950 ;
        RECT 998.100 723.150 999.900 724.950 ;
        RECT 947.100 705.000 948.900 711.000 ;
        RECT 950.100 705.600 951.900 711.600 ;
        RECT 953.100 705.000 954.900 711.600 ;
        RECT 971.100 705.000 972.900 711.600 ;
        RECT 974.100 705.600 975.900 711.600 ;
        RECT 992.100 705.000 993.900 717.600 ;
        RECT 995.400 716.400 999.000 717.600 ;
        RECT 997.200 705.600 999.000 716.400 ;
        RECT 1019.700 711.600 1020.900 724.950 ;
        RECT 1033.950 724.800 1036.050 725.550 ;
        RECT 1016.100 705.000 1017.900 711.600 ;
        RECT 1019.100 705.600 1020.900 711.600 ;
        RECT 1022.100 705.000 1023.900 711.600 ;
        RECT 17.100 689.400 18.900 701.400 ;
        RECT 20.100 691.200 21.900 702.000 ;
        RECT 23.100 695.400 24.900 701.400 ;
        RECT 26.700 695.400 28.500 702.000 ;
        RECT 29.700 696.300 31.500 701.400 ;
        RECT 29.400 695.400 31.500 696.300 ;
        RECT 32.700 695.400 34.500 702.000 ;
        RECT 17.100 682.050 18.300 689.400 ;
        RECT 23.700 688.500 24.900 695.400 ;
        RECT 29.400 694.500 30.300 695.400 ;
        RECT 19.200 687.600 24.900 688.500 ;
        RECT 26.700 693.600 30.300 694.500 ;
        RECT 19.200 686.700 21.000 687.600 ;
        RECT 17.100 679.950 19.200 682.050 ;
        RECT 17.100 672.600 18.300 679.950 ;
        RECT 20.100 675.300 21.000 686.700 ;
        RECT 22.800 682.050 24.600 683.850 ;
        RECT 22.500 679.950 24.600 682.050 ;
        RECT 19.200 674.400 21.000 675.300 ;
        RECT 26.700 677.400 27.900 693.600 ;
        RECT 31.200 692.400 33.000 692.700 ;
        RECT 35.700 692.400 37.500 701.400 ;
        RECT 38.700 695.400 40.500 702.000 ;
        RECT 42.300 698.400 44.100 701.400 ;
        RECT 45.300 698.400 47.100 701.400 ;
        RECT 42.300 696.300 44.400 698.400 ;
        RECT 45.300 696.300 47.400 698.400 ;
        RECT 48.300 695.400 50.100 701.400 ;
        RECT 51.300 695.400 53.100 702.000 ;
        RECT 47.700 693.300 49.800 695.400 ;
        RECT 55.200 693.900 57.000 701.400 ;
        RECT 58.200 695.400 60.000 702.000 ;
        RECT 61.200 695.400 63.000 701.400 ;
        RECT 64.200 698.400 66.000 701.400 ;
        RECT 67.200 698.400 69.000 701.400 ;
        RECT 70.200 698.400 72.000 701.400 ;
        RECT 64.200 696.300 66.300 698.400 ;
        RECT 67.200 696.300 69.300 698.400 ;
        RECT 70.200 696.300 72.300 698.400 ;
        RECT 73.200 695.400 75.000 702.000 ;
        RECT 76.200 695.400 78.000 701.400 ;
        RECT 79.200 695.400 81.000 702.000 ;
        RECT 82.200 695.400 84.000 701.400 ;
        RECT 85.200 695.400 87.000 702.000 ;
        RECT 88.500 695.400 90.300 701.400 ;
        RECT 91.500 695.400 93.300 702.000 ;
        RECT 31.200 691.200 50.400 692.400 ;
        RECT 55.200 691.800 58.500 693.900 ;
        RECT 61.200 691.500 63.900 695.400 ;
        RECT 67.200 694.500 69.300 695.400 ;
        RECT 67.200 693.300 75.300 694.500 ;
        RECT 73.500 692.700 75.300 693.300 ;
        RECT 76.200 692.400 77.400 695.400 ;
        RECT 82.800 694.500 84.000 695.400 ;
        RECT 82.800 693.600 86.700 694.500 ;
        RECT 80.100 692.400 81.900 693.000 ;
        RECT 31.200 690.900 33.000 691.200 ;
        RECT 49.200 690.600 50.400 691.200 ;
        RECT 64.800 690.600 66.900 691.500 ;
        RECT 34.500 689.700 36.300 690.300 ;
        RECT 44.400 689.700 46.500 690.300 ;
        RECT 34.500 688.500 46.500 689.700 ;
        RECT 49.200 689.400 66.900 690.600 ;
        RECT 70.200 690.300 72.300 691.500 ;
        RECT 76.200 691.200 81.900 692.400 ;
        RECT 85.800 690.300 86.700 693.600 ;
        RECT 70.200 689.400 86.700 690.300 ;
        RECT 44.400 688.200 46.500 688.500 ;
        RECT 49.200 687.300 84.900 688.500 ;
        RECT 49.200 686.700 50.400 687.300 ;
        RECT 83.100 686.700 84.900 687.300 ;
        RECT 36.900 685.800 50.400 686.700 ;
        RECT 61.800 685.800 63.900 686.100 ;
        RECT 36.900 685.050 38.700 685.800 ;
        RECT 28.800 682.950 30.900 685.050 ;
        RECT 34.800 683.250 38.700 685.050 ;
        RECT 56.400 684.300 58.500 685.200 ;
        RECT 34.800 682.950 36.900 683.250 ;
        RECT 47.400 683.100 58.500 684.300 ;
        RECT 60.000 684.000 63.900 685.800 ;
        RECT 68.100 684.300 69.900 686.100 ;
        RECT 69.000 683.100 69.900 684.300 ;
        RECT 29.100 681.300 30.900 682.950 ;
        RECT 47.400 682.500 49.200 683.100 ;
        RECT 56.400 682.200 69.900 683.100 ;
        RECT 72.600 682.800 77.700 684.600 ;
        RECT 79.800 682.950 81.900 685.050 ;
        RECT 72.600 681.300 73.500 682.800 ;
        RECT 29.100 680.100 73.500 681.300 ;
        RECT 79.800 680.100 81.300 682.950 ;
        RECT 44.400 677.400 46.200 679.200 ;
        RECT 52.800 678.000 54.900 679.050 ;
        RECT 74.700 678.600 81.300 680.100 ;
        RECT 26.700 676.200 43.500 677.400 ;
        RECT 19.200 673.500 24.900 674.400 ;
        RECT 17.100 666.600 18.900 672.600 ;
        RECT 20.100 666.000 21.900 672.600 ;
        RECT 23.700 669.600 24.900 673.500 ;
        RECT 23.100 666.600 24.900 669.600 ;
        RECT 26.700 672.600 27.900 676.200 ;
        RECT 41.400 675.300 43.500 676.200 ;
        RECT 30.900 674.700 32.700 675.300 ;
        RECT 30.900 673.500 39.300 674.700 ;
        RECT 37.800 672.600 39.300 673.500 ;
        RECT 44.400 674.400 45.300 677.400 ;
        RECT 49.800 677.100 54.900 678.000 ;
        RECT 49.800 676.200 51.600 677.100 ;
        RECT 52.800 676.950 54.900 677.100 ;
        RECT 59.100 677.100 76.200 678.600 ;
        RECT 59.100 676.500 61.200 677.100 ;
        RECT 59.100 674.700 60.900 676.500 ;
        RECT 77.100 675.900 84.900 677.700 ;
        RECT 44.400 673.200 51.600 674.400 ;
        RECT 46.800 672.600 48.600 673.200 ;
        RECT 50.700 672.600 51.600 673.200 ;
        RECT 66.300 672.600 72.900 674.400 ;
        RECT 77.100 672.600 78.600 675.900 ;
        RECT 85.800 672.600 86.700 689.400 ;
        RECT 26.700 666.600 28.500 672.600 ;
        RECT 32.100 666.000 33.900 672.600 ;
        RECT 37.500 666.600 39.300 672.600 ;
        RECT 41.700 669.600 43.800 671.700 ;
        RECT 44.700 669.600 46.800 671.700 ;
        RECT 47.700 669.600 49.800 671.700 ;
        RECT 50.700 671.400 53.400 672.600 ;
        RECT 51.600 670.500 53.400 671.400 ;
        RECT 55.200 670.500 57.900 672.600 ;
        RECT 41.700 666.600 43.500 669.600 ;
        RECT 44.700 666.600 46.500 669.600 ;
        RECT 47.700 666.600 49.500 669.600 ;
        RECT 50.700 666.000 52.500 669.600 ;
        RECT 55.200 666.600 57.000 670.500 ;
        RECT 61.200 669.600 63.300 671.700 ;
        RECT 64.200 669.600 66.300 671.700 ;
        RECT 67.200 669.600 69.300 671.700 ;
        RECT 70.200 669.600 72.300 671.700 ;
        RECT 74.400 671.400 78.600 672.600 ;
        RECT 58.200 666.000 60.000 669.600 ;
        RECT 61.200 666.600 63.000 669.600 ;
        RECT 64.200 666.600 66.000 669.600 ;
        RECT 67.200 666.600 69.000 669.600 ;
        RECT 70.200 666.600 72.000 669.600 ;
        RECT 74.400 666.600 76.200 671.400 ;
        RECT 79.500 666.000 81.300 672.600 ;
        RECT 84.900 666.600 86.700 672.600 ;
        RECT 88.500 685.050 90.000 695.400 ;
        RECT 111.000 690.600 112.800 701.400 ;
        RECT 111.000 689.400 114.600 690.600 ;
        RECT 116.100 689.400 117.900 702.000 ;
        RECT 134.400 689.400 136.200 702.000 ;
        RECT 139.500 690.900 141.300 701.400 ;
        RECT 142.500 695.400 144.300 702.000 ;
        RECT 161.100 695.400 162.900 702.000 ;
        RECT 164.100 695.400 165.900 701.400 ;
        RECT 167.100 696.000 168.900 702.000 ;
        RECT 164.400 695.100 165.900 695.400 ;
        RECT 170.100 695.400 171.900 701.400 ;
        RECT 188.100 695.400 189.900 702.000 ;
        RECT 191.100 695.400 192.900 701.400 ;
        RECT 194.100 695.400 195.900 702.000 ;
        RECT 212.100 695.400 213.900 701.400 ;
        RECT 215.100 695.400 216.900 702.000 ;
        RECT 233.100 695.400 234.900 701.400 ;
        RECT 236.100 695.400 237.900 702.000 ;
        RECT 170.100 695.100 171.000 695.400 ;
        RECT 164.400 694.200 171.000 695.100 ;
        RECT 142.200 692.100 144.000 693.900 ;
        RECT 139.500 689.400 141.900 690.900 ;
        RECT 88.500 682.950 90.900 685.050 ;
        RECT 88.500 669.600 90.000 682.950 ;
        RECT 110.100 682.050 111.900 683.850 ;
        RECT 113.700 682.050 114.600 689.400 ;
        RECT 115.950 682.050 117.750 683.850 ;
        RECT 134.100 682.050 135.900 683.850 ;
        RECT 140.700 682.050 141.900 689.400 ;
        RECT 142.950 687.450 145.050 688.050 ;
        RECT 166.950 687.450 169.050 688.050 ;
        RECT 142.950 686.550 169.050 687.450 ;
        RECT 142.950 685.950 145.050 686.550 ;
        RECT 166.950 685.950 169.050 686.550 ;
        RECT 164.100 682.050 165.900 683.850 ;
        RECT 170.100 682.050 171.000 694.200 ;
        RECT 191.700 682.050 192.900 695.400 ;
        RECT 212.700 682.050 213.900 695.400 ;
        RECT 215.100 682.050 216.900 683.850 ;
        RECT 233.700 682.050 234.900 695.400 ;
        RECT 254.100 690.600 255.900 701.400 ;
        RECT 257.100 691.500 258.900 702.000 ;
        RECT 254.100 689.400 258.900 690.600 ;
        RECT 256.800 688.500 258.900 689.400 ;
        RECT 261.600 689.400 263.400 701.400 ;
        RECT 266.100 691.500 267.900 702.000 ;
        RECT 269.100 690.300 270.900 701.400 ;
        RECT 266.400 689.400 270.900 690.300 ;
        RECT 288.000 690.600 289.800 701.400 ;
        RECT 288.000 689.400 291.600 690.600 ;
        RECT 293.100 689.400 294.900 702.000 ;
        RECT 311.100 689.400 312.900 701.400 ;
        RECT 314.100 690.300 315.900 701.400 ;
        RECT 317.100 691.200 318.900 702.000 ;
        RECT 320.100 690.300 321.900 701.400 ;
        RECT 314.100 689.400 321.900 690.300 ;
        RECT 338.100 689.400 339.900 701.400 ;
        RECT 341.100 690.000 342.900 702.000 ;
        RECT 344.100 695.400 345.900 701.400 ;
        RECT 347.100 695.400 348.900 702.000 ;
        RECT 261.600 688.050 262.800 689.400 ;
        RECT 261.300 687.000 262.800 688.050 ;
        RECT 266.400 687.300 268.500 689.400 ;
        RECT 261.300 685.050 262.200 687.000 ;
        RECT 236.100 682.050 237.900 683.850 ;
        RECT 254.400 682.050 256.200 683.850 ;
        RECT 260.100 682.950 262.200 685.050 ;
        RECT 263.100 685.500 265.200 685.800 ;
        RECT 263.100 683.700 267.000 685.500 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 112.950 679.950 115.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 679.950 169.050 682.050 ;
        RECT 169.950 679.950 172.050 682.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 190.950 679.950 193.050 682.050 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 254.100 679.950 256.200 682.050 ;
        RECT 260.700 682.800 262.200 682.950 ;
        RECT 260.700 681.900 263.100 682.800 ;
        RECT 113.700 669.600 114.600 679.950 ;
        RECT 137.100 678.150 138.900 679.950 ;
        RECT 140.700 675.600 141.900 679.950 ;
        RECT 143.100 678.150 144.900 679.950 ;
        RECT 161.100 678.150 162.900 679.950 ;
        RECT 167.100 678.150 168.900 679.950 ;
        RECT 170.100 676.200 171.000 679.950 ;
        RECT 188.100 678.150 189.900 679.950 ;
        RECT 140.700 674.700 144.300 675.600 ;
        RECT 134.100 671.700 141.900 673.050 ;
        RECT 88.500 666.600 90.300 669.600 ;
        RECT 91.500 666.000 93.300 669.600 ;
        RECT 110.100 666.000 111.900 669.600 ;
        RECT 113.100 666.600 114.900 669.600 ;
        RECT 116.100 666.000 117.900 669.600 ;
        RECT 134.100 666.600 135.900 671.700 ;
        RECT 137.100 666.000 138.900 670.800 ;
        RECT 140.100 666.600 141.900 671.700 ;
        RECT 143.100 672.600 144.300 674.700 ;
        RECT 143.100 666.600 144.900 672.600 ;
        RECT 151.950 669.450 154.050 670.050 ;
        RECT 157.950 669.450 160.050 670.050 ;
        RECT 151.950 668.550 160.050 669.450 ;
        RECT 151.950 667.950 154.050 668.550 ;
        RECT 157.950 667.950 160.050 668.550 ;
        RECT 161.100 666.000 162.900 675.600 ;
        RECT 167.700 675.000 171.000 676.200 ;
        RECT 167.700 666.600 169.500 675.000 ;
        RECT 191.700 674.700 192.900 679.950 ;
        RECT 193.950 678.150 195.750 679.950 ;
        RECT 188.700 673.800 192.900 674.700 ;
        RECT 188.700 666.600 190.500 673.800 ;
        RECT 193.800 666.000 195.600 672.600 ;
        RECT 212.700 669.600 213.900 679.950 ;
        RECT 233.700 669.600 234.900 679.950 ;
        RECT 258.900 679.200 260.700 681.000 ;
        RECT 258.900 677.100 261.000 679.200 ;
        RECT 261.900 676.200 263.100 681.900 ;
        RECT 264.000 682.050 265.800 682.500 ;
        RECT 287.100 682.050 288.900 683.850 ;
        RECT 290.700 682.050 291.600 689.400 ;
        RECT 292.950 682.050 294.750 683.850 ;
        RECT 311.400 682.050 312.300 689.400 ;
        RECT 316.950 682.050 318.750 683.850 ;
        RECT 338.700 682.050 339.600 689.400 ;
        RECT 342.000 682.050 343.800 683.850 ;
        RECT 264.000 680.700 270.900 682.050 ;
        RECT 268.800 679.950 270.900 680.700 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 338.100 679.950 340.200 682.050 ;
        RECT 341.400 679.950 343.500 682.050 ;
        RECT 256.800 673.500 258.900 674.700 ;
        RECT 260.100 674.100 263.100 676.200 ;
        RECT 264.000 677.400 265.800 679.200 ;
        RECT 268.800 678.150 270.600 679.950 ;
        RECT 264.000 675.300 266.100 677.400 ;
        RECT 264.000 674.400 270.300 675.300 ;
        RECT 254.100 672.600 258.900 673.500 ;
        RECT 261.900 672.600 263.100 674.100 ;
        RECT 269.100 672.600 270.300 674.400 ;
        RECT 212.100 666.600 213.900 669.600 ;
        RECT 215.100 666.000 216.900 669.600 ;
        RECT 233.100 666.600 234.900 669.600 ;
        RECT 236.100 666.000 237.900 669.600 ;
        RECT 254.100 666.600 255.900 672.600 ;
        RECT 257.100 666.000 258.900 671.700 ;
        RECT 261.600 666.600 263.400 672.600 ;
        RECT 266.100 666.000 267.900 671.700 ;
        RECT 269.100 666.600 270.900 672.600 ;
        RECT 290.700 669.600 291.600 679.950 ;
        RECT 311.400 672.600 312.300 679.950 ;
        RECT 313.950 678.150 315.750 679.950 ;
        RECT 320.100 678.150 321.900 679.950 ;
        RECT 338.700 672.600 339.600 679.950 ;
        RECT 345.000 675.300 345.900 695.400 ;
        RECT 366.000 690.600 367.800 701.400 ;
        RECT 366.000 689.400 369.600 690.600 ;
        RECT 371.100 689.400 372.900 702.000 ;
        RECT 389.400 689.400 391.200 702.000 ;
        RECT 394.500 690.900 396.300 701.400 ;
        RECT 397.500 695.400 399.300 702.000 ;
        RECT 416.700 695.400 418.500 702.000 ;
        RECT 397.200 692.100 399.000 693.900 ;
        RECT 417.000 692.100 418.800 693.900 ;
        RECT 419.700 690.900 421.500 701.400 ;
        RECT 394.500 689.400 396.900 690.900 ;
        RECT 365.100 682.050 366.900 683.850 ;
        RECT 368.700 682.050 369.600 689.400 ;
        RECT 370.950 682.050 372.750 683.850 ;
        RECT 389.100 682.050 390.900 683.850 ;
        RECT 395.700 682.050 396.900 689.400 ;
        RECT 419.100 689.400 421.500 690.900 ;
        RECT 424.800 689.400 426.600 702.000 ;
        RECT 443.100 689.400 444.900 702.000 ;
        RECT 448.200 690.600 450.000 701.400 ;
        RECT 467.700 695.400 469.500 702.000 ;
        RECT 468.000 692.100 469.800 693.900 ;
        RECT 470.700 690.900 472.500 701.400 ;
        RECT 446.400 689.400 450.000 690.600 ;
        RECT 470.100 689.400 472.500 690.900 ;
        RECT 475.800 689.400 477.600 702.000 ;
        RECT 494.100 695.400 495.900 701.400 ;
        RECT 497.100 695.400 498.900 702.000 ;
        RECT 419.100 682.050 420.300 689.400 ;
        RECT 425.100 682.050 426.900 683.850 ;
        RECT 443.250 682.050 445.050 683.850 ;
        RECT 446.400 682.050 447.300 689.400 ;
        RECT 451.950 684.450 456.000 685.050 ;
        RECT 449.100 682.050 450.900 683.850 ;
        RECT 451.950 682.950 456.450 684.450 ;
        RECT 346.800 679.950 348.900 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 370.950 679.950 373.050 682.050 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 394.950 679.950 397.050 682.050 ;
        RECT 397.950 679.950 400.050 682.050 ;
        RECT 415.950 679.950 418.050 682.050 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 442.950 679.950 445.050 682.050 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 448.950 679.950 451.050 682.050 ;
        RECT 346.950 678.150 348.750 679.950 ;
        RECT 340.500 674.400 348.900 675.300 ;
        RECT 340.500 673.500 342.300 674.400 ;
        RECT 311.400 671.400 316.500 672.600 ;
        RECT 287.100 666.000 288.900 669.600 ;
        RECT 290.100 666.600 291.900 669.600 ;
        RECT 293.100 666.000 294.900 669.600 ;
        RECT 311.700 666.000 313.500 669.600 ;
        RECT 314.700 666.600 316.500 671.400 ;
        RECT 319.200 666.000 321.000 672.600 ;
        RECT 338.700 670.800 341.400 672.600 ;
        RECT 339.600 666.600 341.400 670.800 ;
        RECT 342.600 666.000 344.400 672.600 ;
        RECT 347.100 666.600 348.900 674.400 ;
        RECT 368.700 669.600 369.600 679.950 ;
        RECT 392.100 678.150 393.900 679.950 ;
        RECT 395.700 675.600 396.900 679.950 ;
        RECT 398.100 678.150 399.900 679.950 ;
        RECT 416.100 678.150 417.900 679.950 ;
        RECT 419.100 675.600 420.300 679.950 ;
        RECT 422.100 678.150 423.900 679.950 ;
        RECT 395.700 674.700 399.300 675.600 ;
        RECT 389.100 671.700 396.900 673.050 ;
        RECT 365.100 666.000 366.900 669.600 ;
        RECT 368.100 666.600 369.900 669.600 ;
        RECT 371.100 666.000 372.900 669.600 ;
        RECT 389.100 666.600 390.900 671.700 ;
        RECT 392.100 666.000 393.900 670.800 ;
        RECT 395.100 666.600 396.900 671.700 ;
        RECT 398.100 672.600 399.300 674.700 ;
        RECT 416.700 674.700 420.300 675.600 ;
        RECT 416.700 672.600 417.900 674.700 ;
        RECT 398.100 666.600 399.900 672.600 ;
        RECT 416.100 666.600 417.900 672.600 ;
        RECT 419.100 671.700 426.900 673.050 ;
        RECT 419.100 666.600 420.900 671.700 ;
        RECT 422.100 666.000 423.900 670.800 ;
        RECT 425.100 666.600 426.900 671.700 ;
        RECT 446.400 669.600 447.300 679.950 ;
        RECT 455.550 679.050 456.450 682.950 ;
        RECT 470.100 682.050 471.300 689.400 ;
        RECT 481.950 687.450 484.050 688.050 ;
        RECT 487.950 687.450 490.050 688.050 ;
        RECT 481.950 686.550 490.050 687.450 ;
        RECT 481.950 685.950 484.050 686.550 ;
        RECT 487.950 685.950 490.050 686.550 ;
        RECT 476.100 682.050 477.900 683.850 ;
        RECT 494.700 682.050 495.900 695.400 ;
        RECT 516.000 690.600 517.800 701.400 ;
        RECT 516.000 689.400 519.600 690.600 ;
        RECT 521.100 689.400 522.900 702.000 ;
        RECT 539.100 689.400 540.900 701.400 ;
        RECT 542.100 690.300 543.900 701.400 ;
        RECT 545.100 691.200 546.900 702.000 ;
        RECT 548.100 690.300 549.900 701.400 ;
        RECT 542.100 689.400 549.900 690.300 ;
        RECT 566.400 689.400 568.200 702.000 ;
        RECT 571.500 690.900 573.300 701.400 ;
        RECT 574.500 695.400 576.300 702.000 ;
        RECT 593.100 695.400 594.900 702.000 ;
        RECT 596.100 695.400 597.900 701.400 ;
        RECT 599.100 695.400 600.900 702.000 ;
        RECT 574.200 692.100 576.000 693.900 ;
        RECT 571.500 689.400 573.900 690.900 ;
        RECT 497.100 682.050 498.900 683.850 ;
        RECT 515.100 682.050 516.900 683.850 ;
        RECT 518.700 682.050 519.600 689.400 ;
        RECT 520.950 682.050 522.750 683.850 ;
        RECT 539.400 682.050 540.300 689.400 ;
        RECT 544.950 682.050 546.750 683.850 ;
        RECT 566.100 682.050 567.900 683.850 ;
        RECT 572.700 682.050 573.900 689.400 ;
        RECT 596.100 682.050 597.300 695.400 ;
        RECT 617.100 689.400 618.900 701.400 ;
        RECT 620.100 690.300 621.900 701.400 ;
        RECT 623.100 691.200 624.900 702.000 ;
        RECT 626.100 690.300 627.900 701.400 ;
        RECT 628.950 699.450 631.050 700.050 ;
        RECT 640.950 699.450 643.050 700.050 ;
        RECT 628.950 698.550 643.050 699.450 ;
        RECT 628.950 697.950 631.050 698.550 ;
        RECT 640.950 697.950 643.050 698.550 ;
        RECT 644.100 695.400 645.900 702.000 ;
        RECT 647.100 695.400 648.900 701.400 ;
        RECT 650.100 695.400 651.900 702.000 ;
        RECT 658.950 699.450 661.050 700.050 ;
        RECT 664.950 699.450 667.050 700.050 ;
        RECT 658.950 698.550 667.050 699.450 ;
        RECT 658.950 697.950 661.050 698.550 ;
        RECT 664.950 697.950 667.050 698.550 ;
        RECT 668.700 695.400 670.500 702.000 ;
        RECT 620.100 689.400 627.900 690.300 ;
        RECT 612.000 684.450 616.050 685.050 ;
        RECT 611.550 682.950 616.050 684.450 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 472.950 679.950 475.050 682.050 ;
        RECT 475.950 679.950 478.050 682.050 ;
        RECT 493.950 679.950 496.050 682.050 ;
        RECT 496.950 679.950 499.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 517.950 679.950 520.050 682.050 ;
        RECT 520.950 679.950 523.050 682.050 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 544.950 679.950 547.050 682.050 ;
        RECT 547.950 679.950 550.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 571.950 679.950 574.050 682.050 ;
        RECT 574.950 679.950 577.050 682.050 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 451.950 677.550 456.450 679.050 ;
        RECT 467.100 678.150 468.900 679.950 ;
        RECT 451.950 676.950 456.000 677.550 ;
        RECT 470.100 675.600 471.300 679.950 ;
        RECT 473.100 678.150 474.900 679.950 ;
        RECT 467.700 674.700 471.300 675.600 ;
        RECT 467.700 672.600 468.900 674.700 ;
        RECT 443.100 666.000 444.900 669.600 ;
        RECT 446.100 666.600 447.900 669.600 ;
        RECT 449.100 666.000 450.900 669.600 ;
        RECT 467.100 666.600 468.900 672.600 ;
        RECT 470.100 671.700 477.900 673.050 ;
        RECT 470.100 666.600 471.900 671.700 ;
        RECT 473.100 666.000 474.900 670.800 ;
        RECT 476.100 666.600 477.900 671.700 ;
        RECT 494.700 669.600 495.900 679.950 ;
        RECT 518.700 669.600 519.600 679.950 ;
        RECT 539.400 672.600 540.300 679.950 ;
        RECT 541.950 678.150 543.750 679.950 ;
        RECT 548.100 678.150 549.900 679.950 ;
        RECT 569.100 678.150 570.900 679.950 ;
        RECT 544.950 675.450 547.050 676.050 ;
        RECT 550.950 675.450 553.050 676.050 ;
        RECT 556.950 675.450 559.050 676.050 ;
        RECT 544.950 674.550 559.050 675.450 ;
        RECT 572.700 675.600 573.900 679.950 ;
        RECT 575.100 678.150 576.900 679.950 ;
        RECT 593.250 678.150 595.050 679.950 ;
        RECT 572.700 674.700 576.300 675.600 ;
        RECT 544.950 673.950 547.050 674.550 ;
        RECT 550.950 673.950 553.050 674.550 ;
        RECT 556.950 673.950 559.050 674.550 ;
        RECT 539.400 671.400 544.500 672.600 ;
        RECT 494.100 666.600 495.900 669.600 ;
        RECT 497.100 666.000 498.900 669.600 ;
        RECT 515.100 666.000 516.900 669.600 ;
        RECT 518.100 666.600 519.900 669.600 ;
        RECT 521.100 666.000 522.900 669.600 ;
        RECT 539.700 666.000 541.500 669.600 ;
        RECT 542.700 666.600 544.500 671.400 ;
        RECT 547.200 666.000 549.000 672.600 ;
        RECT 566.100 671.700 573.900 673.050 ;
        RECT 566.100 666.600 567.900 671.700 ;
        RECT 569.100 666.000 570.900 670.800 ;
        RECT 572.100 666.600 573.900 671.700 ;
        RECT 575.100 672.600 576.300 674.700 ;
        RECT 596.100 674.700 597.300 679.950 ;
        RECT 599.100 678.150 600.900 679.950 ;
        RECT 601.950 678.450 604.050 679.050 ;
        RECT 611.550 678.450 612.450 682.950 ;
        RECT 617.400 682.050 618.300 689.400 ;
        RECT 622.950 682.050 624.750 683.850 ;
        RECT 647.700 682.050 648.900 695.400 ;
        RECT 669.000 692.100 670.800 693.900 ;
        RECT 671.700 690.900 673.500 701.400 ;
        RECT 671.100 689.400 673.500 690.900 ;
        RECT 676.800 689.400 678.600 702.000 ;
        RECT 695.100 689.400 696.900 701.400 ;
        RECT 698.100 690.300 699.900 701.400 ;
        RECT 701.100 691.200 702.900 702.000 ;
        RECT 704.100 690.300 705.900 701.400 ;
        RECT 722.700 695.400 724.500 702.000 ;
        RECT 706.950 693.450 709.050 694.050 ;
        RECT 718.950 693.450 721.050 694.050 ;
        RECT 706.950 692.550 721.050 693.450 ;
        RECT 706.950 691.950 709.050 692.550 ;
        RECT 718.950 691.950 721.050 692.550 ;
        RECT 723.000 692.100 724.800 693.900 ;
        RECT 698.100 689.400 705.900 690.300 ;
        RECT 709.950 690.450 712.050 691.050 ;
        RECT 721.950 690.450 724.050 691.050 ;
        RECT 725.700 690.900 727.500 701.400 ;
        RECT 709.950 689.550 724.050 690.450 ;
        RECT 649.950 687.450 652.050 688.050 ;
        RECT 664.950 687.450 667.050 688.050 ;
        RECT 649.950 686.550 667.050 687.450 ;
        RECT 649.950 685.950 652.050 686.550 ;
        RECT 664.950 685.950 667.050 686.550 ;
        RECT 671.100 682.050 672.300 689.400 ;
        RECT 673.950 687.450 676.050 688.050 ;
        RECT 685.950 687.450 688.050 688.050 ;
        RECT 673.950 686.550 688.050 687.450 ;
        RECT 673.950 685.950 676.050 686.550 ;
        RECT 685.950 685.950 688.050 686.550 ;
        RECT 679.950 684.450 684.000 685.050 ;
        RECT 690.000 684.450 694.050 685.050 ;
        RECT 677.100 682.050 678.900 683.850 ;
        RECT 679.950 682.950 684.450 684.450 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 619.950 679.950 622.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 601.950 677.550 612.450 678.450 ;
        RECT 601.950 676.950 604.050 677.550 ;
        RECT 596.100 673.800 600.300 674.700 ;
        RECT 575.100 666.600 576.900 672.600 ;
        RECT 593.400 666.000 595.200 672.600 ;
        RECT 598.500 666.600 600.300 673.800 ;
        RECT 617.400 672.600 618.300 679.950 ;
        RECT 619.950 678.150 621.750 679.950 ;
        RECT 626.100 678.150 627.900 679.950 ;
        RECT 644.100 678.150 645.900 679.950 ;
        RECT 647.700 674.700 648.900 679.950 ;
        RECT 649.950 678.150 651.750 679.950 ;
        RECT 668.100 678.150 669.900 679.950 ;
        RECT 671.100 675.600 672.300 679.950 ;
        RECT 674.100 678.150 675.900 679.950 ;
        RECT 683.550 679.050 684.450 682.950 ;
        RECT 679.950 677.550 684.450 679.050 ;
        RECT 689.550 682.950 694.050 684.450 ;
        RECT 689.550 679.050 690.450 682.950 ;
        RECT 695.400 682.050 696.300 689.400 ;
        RECT 709.950 688.950 712.050 689.550 ;
        RECT 721.950 688.950 724.050 689.550 ;
        RECT 725.100 689.400 727.500 690.900 ;
        RECT 730.800 689.400 732.600 702.000 ;
        RECT 736.950 699.450 739.050 700.050 ;
        RECT 745.950 699.450 748.050 700.050 ;
        RECT 736.950 698.550 748.050 699.450 ;
        RECT 736.950 697.950 739.050 698.550 ;
        RECT 745.950 697.950 748.050 698.550 ;
        RECT 749.400 689.400 751.200 702.000 ;
        RECT 754.500 690.900 756.300 701.400 ;
        RECT 757.500 695.400 759.300 702.000 ;
        RECT 776.100 700.500 783.900 701.400 ;
        RECT 757.200 692.100 759.000 693.900 ;
        RECT 754.500 689.400 756.900 690.900 ;
        RECT 776.100 689.400 777.900 700.500 ;
        RECT 697.950 687.450 700.050 688.050 ;
        RECT 721.950 687.450 724.050 687.900 ;
        RECT 697.950 686.550 724.050 687.450 ;
        RECT 697.950 685.950 700.050 686.550 ;
        RECT 721.950 685.800 724.050 686.550 ;
        RECT 717.000 684.450 721.050 685.050 ;
        RECT 700.950 682.050 702.750 683.850 ;
        RECT 716.550 682.950 721.050 684.450 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 689.550 677.550 694.050 679.050 ;
        RECT 679.950 676.950 684.000 677.550 ;
        RECT 690.000 676.950 694.050 677.550 ;
        RECT 644.700 673.800 648.900 674.700 ;
        RECT 668.700 674.700 672.300 675.600 ;
        RECT 617.400 671.400 622.500 672.600 ;
        RECT 617.700 666.000 619.500 669.600 ;
        RECT 620.700 666.600 622.500 671.400 ;
        RECT 625.200 666.000 627.000 672.600 ;
        RECT 644.700 666.600 646.500 673.800 ;
        RECT 668.700 672.600 669.900 674.700 ;
        RECT 649.800 666.000 651.600 672.600 ;
        RECT 668.100 666.600 669.900 672.600 ;
        RECT 671.100 671.700 678.900 673.050 ;
        RECT 671.100 666.600 672.900 671.700 ;
        RECT 674.100 666.000 675.900 670.800 ;
        RECT 677.100 666.600 678.900 671.700 ;
        RECT 695.400 672.600 696.300 679.950 ;
        RECT 697.950 678.150 699.750 679.950 ;
        RECT 704.100 678.150 705.900 679.950 ;
        RECT 716.550 679.050 717.450 682.950 ;
        RECT 725.100 682.050 726.300 689.400 ;
        RECT 727.950 687.450 730.050 688.050 ;
        RECT 745.950 687.450 748.050 688.050 ;
        RECT 727.950 686.550 748.050 687.450 ;
        RECT 727.950 685.950 730.050 686.550 ;
        RECT 745.950 685.950 748.050 686.550 ;
        RECT 731.100 682.050 732.900 683.850 ;
        RECT 749.100 682.050 750.900 683.850 ;
        RECT 755.700 682.050 756.900 689.400 ;
        RECT 779.100 688.500 780.900 699.600 ;
        RECT 782.100 690.600 783.900 700.500 ;
        RECT 785.100 691.500 786.900 702.000 ;
        RECT 788.100 690.600 789.900 701.400 ;
        RECT 806.100 695.400 807.900 701.400 ;
        RECT 809.100 695.400 810.900 702.000 ;
        RECT 827.100 695.400 828.900 701.400 ;
        RECT 830.100 695.400 831.900 702.000 ;
        RECT 848.100 695.400 849.900 702.000 ;
        RECT 851.100 695.400 852.900 701.400 ;
        RECT 854.100 695.400 855.900 702.000 ;
        RECT 872.100 695.400 873.900 701.400 ;
        RECT 875.100 696.000 876.900 702.000 ;
        RECT 782.100 689.700 789.900 690.600 ;
        RECT 779.100 687.600 783.900 688.500 ;
        RECT 779.100 682.050 780.900 683.850 ;
        RECT 783.000 682.050 783.900 687.600 ;
        RECT 784.950 687.450 787.050 688.050 ;
        RECT 784.950 686.550 792.450 687.450 ;
        RECT 784.950 685.950 787.050 686.550 ;
        RECT 791.550 684.450 792.450 686.550 ;
        RECT 796.950 684.450 799.050 685.050 ;
        RECT 784.950 682.050 786.750 683.850 ;
        RECT 791.550 683.550 799.050 684.450 ;
        RECT 796.950 682.950 799.050 683.550 ;
        RECT 806.700 682.050 807.900 695.400 ;
        RECT 809.100 682.050 810.900 683.850 ;
        RECT 827.700 682.050 828.900 695.400 ;
        RECT 843.000 684.450 847.050 685.050 ;
        RECT 830.100 682.050 831.900 683.850 ;
        RECT 842.550 682.950 847.050 684.450 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 751.950 679.950 754.050 682.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 835.950 681.450 838.050 682.050 ;
        RECT 842.550 681.450 843.450 682.950 ;
        RECT 851.700 682.050 852.900 695.400 ;
        RECT 873.000 695.100 873.900 695.400 ;
        RECT 878.100 695.400 879.900 701.400 ;
        RECT 881.100 695.400 882.900 702.000 ;
        RECT 899.700 695.400 901.500 702.000 ;
        RECT 878.100 695.100 879.600 695.400 ;
        RECT 873.000 694.200 879.600 695.100 ;
        RECT 856.950 684.450 861.000 685.050 ;
        RECT 868.950 684.450 871.050 685.050 ;
        RECT 856.950 682.950 861.450 684.450 ;
        RECT 835.950 680.550 843.450 681.450 ;
        RECT 835.950 679.950 838.050 680.550 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 716.550 677.550 721.050 679.050 ;
        RECT 722.100 678.150 723.900 679.950 ;
        RECT 717.000 676.950 721.050 677.550 ;
        RECT 725.100 675.600 726.300 679.950 ;
        RECT 728.100 678.150 729.900 679.950 ;
        RECT 752.100 678.150 753.900 679.950 ;
        RECT 722.700 674.700 726.300 675.600 ;
        RECT 733.950 675.450 736.050 676.050 ;
        RECT 742.950 675.450 745.050 676.050 ;
        RECT 722.700 672.600 723.900 674.700 ;
        RECT 733.950 674.550 745.050 675.450 ;
        RECT 755.700 675.600 756.900 679.950 ;
        RECT 758.100 678.150 759.900 679.950 ;
        RECT 776.100 678.150 777.900 679.950 ;
        RECT 755.700 674.700 759.300 675.600 ;
        RECT 733.950 673.950 736.050 674.550 ;
        RECT 742.950 673.950 745.050 674.550 ;
        RECT 695.400 671.400 700.500 672.600 ;
        RECT 695.700 666.000 697.500 669.600 ;
        RECT 698.700 666.600 700.500 671.400 ;
        RECT 703.200 666.000 705.000 672.600 ;
        RECT 722.100 666.600 723.900 672.600 ;
        RECT 725.100 671.700 732.900 673.050 ;
        RECT 725.100 666.600 726.900 671.700 ;
        RECT 728.100 666.000 729.900 670.800 ;
        RECT 731.100 666.600 732.900 671.700 ;
        RECT 733.950 672.450 736.050 672.900 ;
        RECT 745.950 672.450 748.050 673.050 ;
        RECT 733.950 671.550 748.050 672.450 ;
        RECT 733.950 670.800 736.050 671.550 ;
        RECT 745.950 670.950 748.050 671.550 ;
        RECT 749.100 671.700 756.900 673.050 ;
        RECT 749.100 666.600 750.900 671.700 ;
        RECT 752.100 666.000 753.900 670.800 ;
        RECT 755.100 666.600 756.900 671.700 ;
        RECT 758.100 672.600 759.300 674.700 ;
        RECT 782.700 672.600 783.900 679.950 ;
        RECT 787.950 678.150 789.750 679.950 ;
        RECT 784.950 675.450 787.050 676.050 ;
        RECT 802.950 675.450 805.050 676.050 ;
        RECT 784.950 674.550 805.050 675.450 ;
        RECT 784.950 673.950 787.050 674.550 ;
        RECT 802.950 673.950 805.050 674.550 ;
        RECT 758.100 666.600 759.900 672.600 ;
        RECT 778.500 666.000 780.300 672.600 ;
        RECT 783.000 666.600 784.800 672.600 ;
        RECT 787.500 666.000 789.300 672.600 ;
        RECT 806.700 669.600 807.900 679.950 ;
        RECT 808.950 675.450 811.050 676.050 ;
        RECT 823.950 675.450 826.050 676.050 ;
        RECT 808.950 674.550 826.050 675.450 ;
        RECT 808.950 673.950 811.050 674.550 ;
        RECT 823.950 673.950 826.050 674.550 ;
        RECT 808.950 672.450 811.050 672.900 ;
        RECT 817.950 672.450 820.050 673.050 ;
        RECT 808.950 671.550 820.050 672.450 ;
        RECT 808.950 670.800 811.050 671.550 ;
        RECT 817.950 670.950 820.050 671.550 ;
        RECT 827.700 669.600 828.900 679.950 ;
        RECT 848.100 678.150 849.900 679.950 ;
        RECT 851.700 674.700 852.900 679.950 ;
        RECT 853.950 678.150 855.750 679.950 ;
        RECT 860.550 679.050 861.450 682.950 ;
        RECT 856.950 677.550 861.450 679.050 ;
        RECT 863.550 683.550 871.050 684.450 ;
        RECT 856.950 676.950 861.000 677.550 ;
        RECT 848.700 673.800 852.900 674.700 ;
        RECT 853.950 675.450 856.050 676.050 ;
        RECT 863.550 675.450 864.450 683.550 ;
        RECT 868.950 682.950 871.050 683.550 ;
        RECT 873.000 682.050 873.900 694.200 ;
        RECT 900.000 692.100 901.800 693.900 ;
        RECT 874.950 690.450 877.050 691.050 ;
        RECT 895.950 690.450 898.050 691.050 ;
        RECT 902.700 690.900 904.500 701.400 ;
        RECT 874.950 689.550 898.050 690.450 ;
        RECT 874.950 688.950 877.050 689.550 ;
        RECT 895.950 688.950 898.050 689.550 ;
        RECT 902.100 689.400 904.500 690.900 ;
        RECT 907.800 689.400 909.600 702.000 ;
        RECT 926.100 700.500 933.900 701.400 ;
        RECT 926.100 691.200 927.900 700.500 ;
        RECT 929.100 691.800 930.900 699.600 ;
        RECT 878.100 682.050 879.900 683.850 ;
        RECT 902.100 682.050 903.300 689.400 ;
        RECT 907.950 687.450 910.050 688.050 ;
        RECT 913.950 687.450 916.050 688.050 ;
        RECT 907.950 686.550 916.050 687.450 ;
        RECT 907.950 685.950 910.050 686.550 ;
        RECT 913.950 685.950 916.050 686.550 ;
        RECT 908.100 682.050 909.900 683.850 ;
        RECT 929.700 682.050 930.900 691.800 ;
        RECT 932.100 691.800 933.900 700.500 ;
        RECT 935.100 700.500 942.900 701.400 ;
        RECT 935.100 692.700 936.900 700.500 ;
        RECT 938.100 691.800 939.900 699.600 ;
        RECT 932.100 690.900 939.900 691.800 ;
        RECT 941.100 691.500 942.900 700.500 ;
        RECT 944.100 692.400 945.900 702.000 ;
        RECT 947.100 691.500 948.900 701.400 ;
        RECT 941.100 690.600 948.900 691.500 ;
        RECT 966.000 690.600 967.800 701.400 ;
        RECT 966.000 689.400 969.600 690.600 ;
        RECT 971.100 689.400 972.900 702.000 ;
        RECT 989.100 689.400 990.900 702.000 ;
        RECT 994.200 690.600 996.000 701.400 ;
        RECT 1013.100 695.400 1014.900 701.400 ;
        RECT 1016.100 696.000 1017.900 702.000 ;
        RECT 992.400 689.400 996.000 690.600 ;
        RECT 1014.000 695.100 1014.900 695.400 ;
        RECT 1019.100 695.400 1020.900 701.400 ;
        RECT 1022.100 695.400 1023.900 702.000 ;
        RECT 1019.100 695.100 1020.600 695.400 ;
        RECT 1014.000 694.200 1020.600 695.100 ;
        RECT 934.950 687.450 937.050 688.050 ;
        RECT 934.950 686.550 954.450 687.450 ;
        RECT 934.950 685.950 937.050 686.550 ;
        RECT 946.950 684.450 951.000 685.050 ;
        RECT 934.950 682.050 936.750 683.850 ;
        RECT 944.100 682.050 945.900 683.850 ;
        RECT 946.950 682.950 951.450 684.450 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 929.400 679.950 931.500 682.050 ;
        RECT 934.950 679.950 937.050 682.050 ;
        RECT 937.950 679.950 940.050 682.050 ;
        RECT 944.100 679.950 946.200 682.050 ;
        RECT 853.950 674.550 864.450 675.450 ;
        RECT 873.000 676.200 873.900 679.950 ;
        RECT 875.100 678.150 876.900 679.950 ;
        RECT 881.100 678.150 882.900 679.950 ;
        RECT 899.100 678.150 900.900 679.950 ;
        RECT 873.000 675.000 876.300 676.200 ;
        RECT 902.100 675.600 903.300 679.950 ;
        RECT 905.100 678.150 906.900 679.950 ;
        RECT 910.950 678.450 913.050 679.050 ;
        RECT 925.950 678.450 928.050 679.050 ;
        RECT 910.950 677.550 928.050 678.450 ;
        RECT 910.950 676.950 913.050 677.550 ;
        RECT 925.950 676.950 928.050 677.550 ;
        RECT 853.950 673.950 856.050 674.550 ;
        RECT 806.100 666.600 807.900 669.600 ;
        RECT 809.100 666.000 810.900 669.600 ;
        RECT 827.100 666.600 828.900 669.600 ;
        RECT 830.100 666.000 831.900 669.600 ;
        RECT 848.700 666.600 850.500 673.800 ;
        RECT 853.800 666.000 855.600 672.600 ;
        RECT 856.950 672.450 859.050 673.050 ;
        RECT 868.950 672.450 871.050 673.050 ;
        RECT 856.950 671.550 871.050 672.450 ;
        RECT 856.950 670.950 859.050 671.550 ;
        RECT 868.950 670.950 871.050 671.550 ;
        RECT 874.500 666.600 876.300 675.000 ;
        RECT 881.100 666.000 882.900 675.600 ;
        RECT 899.700 674.700 903.300 675.600 ;
        RECT 899.700 672.600 900.900 674.700 ;
        RECT 899.100 666.600 900.900 672.600 ;
        RECT 902.100 671.700 909.900 673.050 ;
        RECT 902.100 666.600 903.900 671.700 ;
        RECT 905.100 666.000 906.900 670.800 ;
        RECT 908.100 666.600 909.900 671.700 ;
        RECT 929.700 671.400 930.900 679.950 ;
        RECT 938.250 678.150 940.050 679.950 ;
        RECT 950.550 679.050 951.450 682.950 ;
        RECT 946.950 677.550 951.450 679.050 ;
        RECT 953.550 678.450 954.450 686.550 ;
        RECT 965.100 682.050 966.900 683.850 ;
        RECT 968.700 682.050 969.600 689.400 ;
        RECT 970.950 682.050 972.750 683.850 ;
        RECT 989.250 682.050 991.050 683.850 ;
        RECT 992.400 682.050 993.300 689.400 ;
        RECT 995.100 682.050 996.900 683.850 ;
        RECT 1014.000 682.050 1014.900 694.200 ;
        RECT 1024.950 684.450 1029.000 685.050 ;
        RECT 1019.100 682.050 1020.900 683.850 ;
        RECT 1024.950 682.950 1029.450 684.450 ;
        RECT 964.950 679.950 967.050 682.050 ;
        RECT 967.950 679.950 970.050 682.050 ;
        RECT 970.950 679.950 973.050 682.050 ;
        RECT 988.950 679.950 991.050 682.050 ;
        RECT 991.950 679.950 994.050 682.050 ;
        RECT 994.950 679.950 997.050 682.050 ;
        RECT 1012.950 679.950 1015.050 682.050 ;
        RECT 1015.950 679.950 1018.050 682.050 ;
        RECT 1018.950 679.950 1021.050 682.050 ;
        RECT 1021.950 679.950 1024.050 682.050 ;
        RECT 961.950 678.450 964.050 679.050 ;
        RECT 953.550 677.550 964.050 678.450 ;
        RECT 946.950 676.950 951.000 677.550 ;
        RECT 961.950 676.950 964.050 677.550 ;
        RECT 931.950 675.450 934.050 676.050 ;
        RECT 952.950 675.450 955.050 676.050 ;
        RECT 931.950 674.550 955.050 675.450 ;
        RECT 931.950 673.950 934.050 674.550 ;
        RECT 952.950 673.950 955.050 674.550 ;
        RECT 929.700 670.500 942.300 671.400 ;
        RECT 934.200 669.600 935.100 670.500 ;
        RECT 941.400 669.600 942.300 670.500 ;
        RECT 968.700 669.600 969.600 679.950 ;
        RECT 970.950 675.450 973.050 676.050 ;
        RECT 976.950 675.450 979.050 676.050 ;
        RECT 970.950 674.550 979.050 675.450 ;
        RECT 970.950 673.950 973.050 674.550 ;
        RECT 976.950 673.950 979.050 674.550 ;
        RECT 976.950 672.450 979.050 672.900 ;
        RECT 988.950 672.450 991.050 673.050 ;
        RECT 976.950 671.550 991.050 672.450 ;
        RECT 976.950 670.800 979.050 671.550 ;
        RECT 988.950 670.950 991.050 671.550 ;
        RECT 992.400 669.600 993.300 679.950 ;
        RECT 1014.000 676.200 1014.900 679.950 ;
        RECT 1016.100 678.150 1017.900 679.950 ;
        RECT 1022.100 678.150 1023.900 679.950 ;
        RECT 1028.550 679.050 1029.450 682.950 ;
        RECT 1024.950 677.550 1029.450 679.050 ;
        RECT 1024.950 676.950 1029.000 677.550 ;
        RECT 1014.000 675.000 1017.300 676.200 ;
        RECT 934.200 666.600 936.900 669.600 ;
        RECT 938.100 666.000 939.900 669.600 ;
        RECT 941.100 666.600 942.900 669.600 ;
        RECT 944.100 666.000 946.200 669.600 ;
        RECT 965.100 666.000 966.900 669.600 ;
        RECT 968.100 666.600 969.900 669.600 ;
        RECT 971.100 666.000 972.900 669.600 ;
        RECT 989.100 666.000 990.900 669.600 ;
        RECT 992.100 666.600 993.900 669.600 ;
        RECT 995.100 666.000 996.900 669.600 ;
        RECT 1015.500 666.600 1017.300 675.000 ;
        RECT 1022.100 666.000 1023.900 675.600 ;
        RECT 17.100 659.400 18.900 663.000 ;
        RECT 20.100 659.400 21.900 662.400 ;
        RECT 23.100 659.400 24.900 663.000 ;
        RECT 20.700 649.050 21.600 659.400 ;
        RECT 41.100 657.300 42.900 662.400 ;
        RECT 44.100 658.200 45.900 663.000 ;
        RECT 47.100 657.300 48.900 662.400 ;
        RECT 41.100 655.950 48.900 657.300 ;
        RECT 50.100 656.400 51.900 662.400 ;
        RECT 68.100 656.400 69.900 663.000 ;
        RECT 50.100 654.300 51.300 656.400 ;
        RECT 71.100 655.500 72.900 662.400 ;
        RECT 74.100 656.400 75.900 663.000 ;
        RECT 77.100 655.500 78.900 662.400 ;
        RECT 80.100 656.400 81.900 663.000 ;
        RECT 83.100 655.500 84.900 662.400 ;
        RECT 86.100 656.400 87.900 663.000 ;
        RECT 89.100 655.500 90.900 662.400 ;
        RECT 92.100 656.400 93.900 663.000 ;
        RECT 95.700 656.400 97.500 662.400 ;
        RECT 101.100 656.400 102.900 663.000 ;
        RECT 106.500 656.400 108.300 662.400 ;
        RECT 110.700 659.400 112.500 662.400 ;
        RECT 113.700 659.400 115.500 662.400 ;
        RECT 116.700 659.400 118.500 662.400 ;
        RECT 119.700 659.400 121.500 663.000 ;
        RECT 110.700 657.300 112.800 659.400 ;
        RECT 113.700 657.300 115.800 659.400 ;
        RECT 116.700 657.300 118.800 659.400 ;
        RECT 124.200 658.500 126.000 662.400 ;
        RECT 127.200 659.400 129.000 663.000 ;
        RECT 130.200 659.400 132.000 662.400 ;
        RECT 133.200 659.400 135.000 662.400 ;
        RECT 136.200 659.400 138.000 662.400 ;
        RECT 139.200 659.400 141.000 662.400 ;
        RECT 120.600 657.600 122.400 658.500 ;
        RECT 119.700 656.400 122.400 657.600 ;
        RECT 124.200 656.400 126.900 658.500 ;
        RECT 130.200 657.300 132.300 659.400 ;
        RECT 133.200 657.300 135.300 659.400 ;
        RECT 136.200 657.300 138.300 659.400 ;
        RECT 139.200 657.300 141.300 659.400 ;
        RECT 143.400 657.600 145.200 662.400 ;
        RECT 143.400 656.400 147.600 657.600 ;
        RECT 148.500 656.400 150.300 663.000 ;
        RECT 153.900 656.400 155.700 662.400 ;
        RECT 47.700 653.400 51.300 654.300 ;
        RECT 70.050 654.300 72.900 655.500 ;
        RECT 75.000 654.300 78.900 655.500 ;
        RECT 81.000 654.300 84.900 655.500 ;
        RECT 87.000 654.300 90.900 655.500 ;
        RECT 44.100 649.050 45.900 650.850 ;
        RECT 47.700 649.050 48.900 653.400 ;
        RECT 50.100 649.050 51.900 650.850 ;
        RECT 70.050 649.050 71.100 654.300 ;
        RECT 75.000 653.400 76.200 654.300 ;
        RECT 81.000 653.400 82.200 654.300 ;
        RECT 87.000 653.400 88.200 654.300 ;
        RECT 72.000 652.200 76.200 653.400 ;
        RECT 72.000 651.600 73.800 652.200 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 22.950 646.950 25.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 70.050 646.950 73.200 649.050 ;
        RECT 17.100 645.150 18.900 646.950 ;
        RECT 20.700 639.600 21.600 646.950 ;
        RECT 22.950 645.150 24.750 646.950 ;
        RECT 41.100 645.150 42.900 646.950 ;
        RECT 47.700 639.600 48.900 646.950 ;
        RECT 70.050 641.700 71.100 646.950 ;
        RECT 75.000 641.700 76.200 652.200 ;
        RECT 78.000 652.200 82.200 653.400 ;
        RECT 78.000 651.600 79.800 652.200 ;
        RECT 81.000 641.700 82.200 652.200 ;
        RECT 84.000 652.200 88.200 653.400 ;
        RECT 84.000 651.600 85.800 652.200 ;
        RECT 87.000 641.700 88.200 652.200 ;
        RECT 95.700 652.800 96.900 656.400 ;
        RECT 106.800 655.500 108.300 656.400 ;
        RECT 115.800 655.800 117.600 656.400 ;
        RECT 119.700 655.800 120.600 656.400 ;
        RECT 99.900 654.300 108.300 655.500 ;
        RECT 113.400 654.600 120.600 655.800 ;
        RECT 135.300 654.600 141.900 656.400 ;
        RECT 99.900 653.700 101.700 654.300 ;
        RECT 110.400 652.800 112.500 653.700 ;
        RECT 95.700 651.600 112.500 652.800 ;
        RECT 113.400 651.600 114.300 654.600 ;
        RECT 118.800 651.900 120.600 652.800 ;
        RECT 128.100 652.500 129.900 654.300 ;
        RECT 146.100 653.100 147.600 656.400 ;
        RECT 121.800 651.900 123.900 652.050 ;
        RECT 89.400 649.050 91.200 650.850 ;
        RECT 89.100 646.950 91.200 649.050 ;
        RECT 70.050 640.500 72.900 641.700 ;
        RECT 75.000 640.500 78.900 641.700 ;
        RECT 81.000 640.500 84.900 641.700 ;
        RECT 87.000 640.500 90.900 641.700 ;
        RECT 18.000 638.400 21.600 639.600 ;
        RECT 18.000 627.600 19.800 638.400 ;
        RECT 23.100 627.000 24.900 639.600 ;
        RECT 41.400 627.000 43.200 639.600 ;
        RECT 46.500 638.100 48.900 639.600 ;
        RECT 46.500 627.600 48.300 638.100 ;
        RECT 49.200 635.100 51.000 636.900 ;
        RECT 49.500 627.000 51.300 633.600 ;
        RECT 68.100 627.000 69.900 639.600 ;
        RECT 71.100 627.600 72.900 640.500 ;
        RECT 74.100 627.000 75.900 639.600 ;
        RECT 77.100 627.600 78.900 640.500 ;
        RECT 80.100 627.000 81.900 639.600 ;
        RECT 83.100 627.600 84.900 640.500 ;
        RECT 86.100 627.000 87.900 639.600 ;
        RECT 89.100 627.600 90.900 640.500 ;
        RECT 92.100 627.000 93.900 639.600 ;
        RECT 95.700 635.400 96.900 651.600 ;
        RECT 113.400 649.800 115.200 651.600 ;
        RECT 118.800 651.000 123.900 651.900 ;
        RECT 121.800 649.950 123.900 651.000 ;
        RECT 128.100 651.900 130.200 652.500 ;
        RECT 128.100 650.400 145.200 651.900 ;
        RECT 146.100 651.300 153.900 653.100 ;
        RECT 143.700 648.900 150.300 650.400 ;
        RECT 98.100 647.700 142.500 648.900 ;
        RECT 98.100 646.050 99.900 647.700 ;
        RECT 97.800 643.950 99.900 646.050 ;
        RECT 103.800 645.750 105.900 646.050 ;
        RECT 116.400 645.900 118.200 646.500 ;
        RECT 125.400 645.900 138.900 646.800 ;
        RECT 103.800 643.950 107.700 645.750 ;
        RECT 116.400 644.700 127.500 645.900 ;
        RECT 105.900 643.200 107.700 643.950 ;
        RECT 125.400 643.800 127.500 644.700 ;
        RECT 129.000 643.200 132.900 645.000 ;
        RECT 138.000 644.700 138.900 645.900 ;
        RECT 105.900 642.300 119.400 643.200 ;
        RECT 130.800 642.900 132.900 643.200 ;
        RECT 137.100 642.900 138.900 644.700 ;
        RECT 141.600 646.200 142.500 647.700 ;
        RECT 141.600 644.400 146.700 646.200 ;
        RECT 148.800 646.050 150.300 648.900 ;
        RECT 148.800 643.950 150.900 646.050 ;
        RECT 118.200 641.700 119.400 642.300 ;
        RECT 152.100 641.700 153.900 642.300 ;
        RECT 113.400 640.500 115.500 640.800 ;
        RECT 118.200 640.500 153.900 641.700 ;
        RECT 103.500 639.300 115.500 640.500 ;
        RECT 154.800 639.600 155.700 656.400 ;
        RECT 103.500 638.700 105.300 639.300 ;
        RECT 113.400 638.700 115.500 639.300 ;
        RECT 118.200 638.400 135.900 639.600 ;
        RECT 100.200 637.800 102.000 638.100 ;
        RECT 118.200 637.800 119.400 638.400 ;
        RECT 100.200 636.600 119.400 637.800 ;
        RECT 133.800 637.500 135.900 638.400 ;
        RECT 139.200 638.700 155.700 639.600 ;
        RECT 139.200 637.500 141.300 638.700 ;
        RECT 100.200 636.300 102.000 636.600 ;
        RECT 95.700 634.500 99.300 635.400 ;
        RECT 98.400 633.600 99.300 634.500 ;
        RECT 95.700 627.000 97.500 633.600 ;
        RECT 98.400 632.700 100.500 633.600 ;
        RECT 98.700 627.600 100.500 632.700 ;
        RECT 101.700 627.000 103.500 633.600 ;
        RECT 104.700 627.600 106.500 636.600 ;
        RECT 116.700 633.600 118.800 635.700 ;
        RECT 124.200 635.100 127.500 637.200 ;
        RECT 107.700 627.000 109.500 633.600 ;
        RECT 111.300 630.600 113.400 632.700 ;
        RECT 114.300 630.600 116.400 632.700 ;
        RECT 111.300 627.600 113.100 630.600 ;
        RECT 114.300 627.600 116.100 630.600 ;
        RECT 117.300 627.600 119.100 633.600 ;
        RECT 120.300 627.000 122.100 633.600 ;
        RECT 124.200 627.600 126.000 635.100 ;
        RECT 130.200 633.600 132.900 637.500 ;
        RECT 145.200 636.600 150.900 637.800 ;
        RECT 142.500 635.700 144.300 636.300 ;
        RECT 136.200 634.500 144.300 635.700 ;
        RECT 136.200 633.600 138.300 634.500 ;
        RECT 145.200 633.600 146.400 636.600 ;
        RECT 149.100 636.000 150.900 636.600 ;
        RECT 154.800 635.400 155.700 638.700 ;
        RECT 151.800 634.500 155.700 635.400 ;
        RECT 157.500 659.400 159.300 662.400 ;
        RECT 160.500 659.400 162.300 663.000 ;
        RECT 179.100 659.400 180.900 663.000 ;
        RECT 182.100 659.400 183.900 662.400 ;
        RECT 185.100 659.400 186.900 663.000 ;
        RECT 203.100 659.400 204.900 663.000 ;
        RECT 206.100 659.400 207.900 662.400 ;
        RECT 157.500 646.050 159.000 659.400 ;
        RECT 182.400 649.050 183.300 659.400 ;
        RECT 206.100 649.050 207.300 659.400 ;
        RECT 226.500 654.000 228.300 662.400 ;
        RECT 225.000 652.800 228.300 654.000 ;
        RECT 233.100 653.400 234.900 663.000 ;
        RECT 251.100 657.300 252.900 662.400 ;
        RECT 254.100 658.200 255.900 663.000 ;
        RECT 257.100 657.300 258.900 662.400 ;
        RECT 251.100 655.950 258.900 657.300 ;
        RECT 260.100 656.400 261.900 662.400 ;
        RECT 278.100 657.300 279.900 662.400 ;
        RECT 281.100 658.200 282.900 663.000 ;
        RECT 284.100 657.300 285.900 662.400 ;
        RECT 260.100 654.300 261.300 656.400 ;
        RECT 278.100 655.950 285.900 657.300 ;
        RECT 287.100 656.400 288.900 662.400 ;
        RECT 305.700 659.400 307.500 663.000 ;
        RECT 308.700 657.600 310.500 662.400 ;
        RECT 305.400 656.400 310.500 657.600 ;
        RECT 313.200 656.400 315.000 663.000 ;
        RECT 287.100 654.300 288.300 656.400 ;
        RECT 257.700 653.400 261.300 654.300 ;
        RECT 284.700 653.400 288.300 654.300 ;
        RECT 225.000 649.050 225.900 652.800 ;
        RECT 227.100 649.050 228.900 650.850 ;
        RECT 233.100 649.050 234.900 650.850 ;
        RECT 254.100 649.050 255.900 650.850 ;
        RECT 257.700 649.050 258.900 653.400 ;
        RECT 260.100 649.050 261.900 650.850 ;
        RECT 281.100 649.050 282.900 650.850 ;
        RECT 284.700 649.050 285.900 653.400 ;
        RECT 289.950 651.450 292.050 652.050 ;
        RECT 295.950 651.450 298.050 652.050 ;
        RECT 287.100 649.050 288.900 650.850 ;
        RECT 289.950 650.550 298.050 651.450 ;
        RECT 289.950 649.950 292.050 650.550 ;
        RECT 295.950 649.950 298.050 650.550 ;
        RECT 305.400 649.050 306.300 656.400 ;
        RECT 310.950 654.450 313.050 655.050 ;
        RECT 325.950 654.450 328.050 655.050 ;
        RECT 310.950 653.550 328.050 654.450 ;
        RECT 310.950 652.950 313.050 653.550 ;
        RECT 325.950 652.950 328.050 653.550 ;
        RECT 332.100 653.400 333.900 663.000 ;
        RECT 338.700 654.000 340.500 662.400 ;
        RECT 359.100 659.400 360.900 663.000 ;
        RECT 362.100 659.400 363.900 662.400 ;
        RECT 365.100 659.400 366.900 663.000 ;
        RECT 338.700 652.800 342.000 654.000 ;
        RECT 307.950 649.050 309.750 650.850 ;
        RECT 314.100 649.050 315.900 650.850 ;
        RECT 332.100 649.050 333.900 650.850 ;
        RECT 338.100 649.050 339.900 650.850 ;
        RECT 341.100 649.050 342.000 652.800 ;
        RECT 346.950 651.450 349.050 652.050 ;
        RECT 355.950 651.450 358.050 652.050 ;
        RECT 346.950 650.550 358.050 651.450 ;
        RECT 346.950 649.950 349.050 650.550 ;
        RECT 355.950 649.950 358.050 650.550 ;
        RECT 362.400 649.050 363.300 659.400 ;
        RECT 383.400 656.400 385.200 663.000 ;
        RECT 388.500 655.200 390.300 662.400 ;
        RECT 407.400 656.400 409.200 663.000 ;
        RECT 412.500 655.200 414.300 662.400 ;
        RECT 431.100 659.400 432.900 663.000 ;
        RECT 434.100 659.400 435.900 662.400 ;
        RECT 437.100 659.400 438.900 663.000 ;
        RECT 386.100 654.300 390.300 655.200 ;
        RECT 410.100 654.300 414.300 655.200 ;
        RECT 421.950 654.450 424.050 655.050 ;
        RECT 430.950 654.450 433.050 655.200 ;
        RECT 383.250 649.050 385.050 650.850 ;
        RECT 386.100 649.050 387.300 654.300 ;
        RECT 389.100 649.050 390.900 650.850 ;
        RECT 407.250 649.050 409.050 650.850 ;
        RECT 410.100 649.050 411.300 654.300 ;
        RECT 421.950 653.550 433.050 654.450 ;
        RECT 421.950 652.950 424.050 653.550 ;
        RECT 430.950 653.100 433.050 653.550 ;
        RECT 413.100 649.050 414.900 650.850 ;
        RECT 434.700 649.050 435.600 659.400 ;
        RECT 455.400 656.400 457.200 663.000 ;
        RECT 460.500 655.200 462.300 662.400 ;
        RECT 479.400 656.400 481.200 663.000 ;
        RECT 484.500 655.200 486.300 662.400 ;
        RECT 504.000 656.400 505.800 663.000 ;
        RECT 508.500 657.600 510.300 662.400 ;
        RECT 511.500 659.400 513.300 663.000 ;
        RECT 530.100 659.400 531.900 663.000 ;
        RECT 533.100 659.400 534.900 662.400 ;
        RECT 536.100 659.400 537.900 663.000 ;
        RECT 554.100 659.400 555.900 663.000 ;
        RECT 557.100 659.400 558.900 662.400 ;
        RECT 508.500 656.400 513.600 657.600 ;
        RECT 458.100 654.300 462.300 655.200 ;
        RECT 482.100 654.300 486.300 655.200 ;
        RECT 455.250 649.050 457.050 650.850 ;
        RECT 458.100 649.050 459.300 654.300 ;
        RECT 461.100 649.050 462.900 650.850 ;
        RECT 479.250 649.050 481.050 650.850 ;
        RECT 482.100 649.050 483.300 654.300 ;
        RECT 485.100 649.050 486.900 650.850 ;
        RECT 503.100 649.050 504.900 650.850 ;
        RECT 509.250 649.050 511.050 650.850 ;
        RECT 512.700 649.050 513.600 656.400 ;
        RECT 533.700 649.050 534.600 659.400 ;
        RECT 557.100 649.050 558.300 659.400 ;
        RECT 575.700 655.200 577.500 662.400 ;
        RECT 580.800 656.400 582.600 663.000 ;
        RECT 599.700 655.200 601.500 662.400 ;
        RECT 604.800 656.400 606.600 663.000 ;
        RECT 575.700 654.300 579.900 655.200 ;
        RECT 599.700 654.300 603.900 655.200 ;
        RECT 575.100 649.050 576.900 650.850 ;
        RECT 578.700 649.050 579.900 654.300 ;
        RECT 580.950 649.050 582.750 650.850 ;
        RECT 599.100 649.050 600.900 650.850 ;
        RECT 602.700 649.050 603.900 654.300 ;
        RECT 625.500 654.000 627.300 662.400 ;
        RECT 624.000 652.800 627.300 654.000 ;
        RECT 632.100 653.400 633.900 663.000 ;
        RECT 651.000 656.400 652.800 663.000 ;
        RECT 655.500 657.600 657.300 662.400 ;
        RECT 658.500 659.400 660.300 663.000 ;
        RECT 677.100 659.400 678.900 663.000 ;
        RECT 680.100 659.400 681.900 662.400 ;
        RECT 683.100 659.400 684.900 663.000 ;
        RECT 655.500 656.400 660.600 657.600 ;
        RECT 604.950 649.050 606.750 650.850 ;
        RECT 624.000 649.050 624.900 652.800 ;
        RECT 626.100 649.050 627.900 650.850 ;
        RECT 632.100 649.050 633.900 650.850 ;
        RECT 650.100 649.050 651.900 650.850 ;
        RECT 656.250 649.050 658.050 650.850 ;
        RECT 659.700 649.050 660.600 656.400 ;
        RECT 680.700 649.050 681.600 659.400 ;
        RECT 701.700 655.200 703.500 662.400 ;
        RECT 706.800 656.400 708.600 663.000 ;
        RECT 727.500 656.400 729.300 663.000 ;
        RECT 732.000 656.400 733.800 662.400 ;
        RECT 736.500 656.400 738.300 663.000 ;
        RECT 755.100 661.500 762.900 662.400 ;
        RECT 755.100 656.400 756.900 661.500 ;
        RECT 758.100 656.400 759.900 660.600 ;
        RECT 761.100 657.000 762.900 661.500 ;
        RECT 764.100 657.900 765.900 663.000 ;
        RECT 767.100 657.000 768.900 662.400 ;
        RECT 701.700 654.300 705.900 655.200 ;
        RECT 701.100 649.050 702.900 650.850 ;
        RECT 704.700 649.050 705.900 654.300 ;
        RECT 706.950 649.050 708.750 650.850 ;
        RECT 725.100 649.050 726.900 650.850 ;
        RECT 731.700 649.050 732.900 656.400 ;
        RECT 758.700 654.900 759.600 656.400 ;
        RECT 761.100 656.100 768.900 657.000 ;
        RECT 787.500 656.400 789.300 663.000 ;
        RECT 792.000 656.400 793.800 662.400 ;
        RECT 796.500 656.400 798.300 663.000 ;
        RECT 815.100 659.400 816.900 663.000 ;
        RECT 818.100 659.400 819.900 662.400 ;
        RECT 821.100 659.400 822.900 663.000 ;
        RECT 839.700 659.400 841.500 663.000 ;
        RECT 758.700 653.700 763.050 654.900 ;
        RECT 745.950 651.450 748.050 651.900 ;
        RECT 751.950 651.450 754.050 652.050 ;
        RECT 736.950 649.050 738.750 650.850 ;
        RECT 745.950 650.550 754.050 651.450 ;
        RECT 745.950 649.800 748.050 650.550 ;
        RECT 751.950 649.950 754.050 650.550 ;
        RECT 758.250 649.050 760.050 650.850 ;
        RECT 762.000 649.050 763.050 653.700 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 232.950 646.950 235.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 256.950 646.950 259.050 649.050 ;
        RECT 259.950 646.950 262.050 649.050 ;
        RECT 277.950 646.950 280.050 649.050 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 307.950 646.950 310.050 649.050 ;
        RECT 310.950 646.950 313.050 649.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 340.950 646.950 343.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 532.950 646.950 535.050 649.050 ;
        RECT 535.950 646.950 538.050 649.050 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 556.950 646.950 559.050 649.050 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 598.950 646.950 601.050 649.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 658.950 646.950 661.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 706.950 646.950 709.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 649.050 765.750 650.850 ;
        RECT 785.100 649.050 786.900 650.850 ;
        RECT 791.700 649.050 792.900 656.400 ;
        RECT 810.000 651.450 814.050 652.050 ;
        RECT 796.950 649.050 798.750 650.850 ;
        RECT 809.550 649.950 814.050 651.450 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 157.500 643.950 159.900 646.050 ;
        RECT 179.250 645.150 181.050 646.950 ;
        RECT 151.800 633.600 153.000 634.500 ;
        RECT 157.500 633.600 159.000 643.950 ;
        RECT 182.400 639.600 183.300 646.950 ;
        RECT 185.100 645.150 186.900 646.950 ;
        RECT 203.100 645.150 204.900 646.950 ;
        RECT 127.200 627.000 129.000 633.600 ;
        RECT 130.200 627.600 132.000 633.600 ;
        RECT 133.200 630.600 135.300 632.700 ;
        RECT 136.200 630.600 138.300 632.700 ;
        RECT 139.200 630.600 141.300 632.700 ;
        RECT 133.200 627.600 135.000 630.600 ;
        RECT 136.200 627.600 138.000 630.600 ;
        RECT 139.200 627.600 141.000 630.600 ;
        RECT 142.200 627.000 144.000 633.600 ;
        RECT 145.200 627.600 147.000 633.600 ;
        RECT 148.200 627.000 150.000 633.600 ;
        RECT 151.200 627.600 153.000 633.600 ;
        RECT 154.200 627.000 156.000 633.600 ;
        RECT 157.500 627.600 159.300 633.600 ;
        RECT 160.500 627.000 162.300 633.600 ;
        RECT 179.100 627.000 180.900 639.600 ;
        RECT 182.400 638.400 186.000 639.600 ;
        RECT 184.200 627.600 186.000 638.400 ;
        RECT 206.100 633.600 207.300 646.950 ;
        RECT 225.000 634.800 225.900 646.950 ;
        RECT 230.100 645.150 231.900 646.950 ;
        RECT 251.100 645.150 252.900 646.950 ;
        RECT 226.950 642.450 229.050 642.750 ;
        RECT 253.950 642.450 256.050 643.050 ;
        RECT 226.950 641.550 256.050 642.450 ;
        RECT 226.950 640.650 229.050 641.550 ;
        RECT 253.950 640.950 256.050 641.550 ;
        RECT 257.700 639.600 258.900 646.950 ;
        RECT 278.100 645.150 279.900 646.950 ;
        RECT 284.700 639.600 285.900 646.950 ;
        RECT 305.400 639.600 306.300 646.950 ;
        RECT 310.950 645.150 312.750 646.950 ;
        RECT 335.100 645.150 336.900 646.950 ;
        RECT 225.000 633.900 231.600 634.800 ;
        RECT 225.000 633.600 225.900 633.900 ;
        RECT 203.100 627.000 204.900 633.600 ;
        RECT 206.100 627.600 207.900 633.600 ;
        RECT 224.100 627.600 225.900 633.600 ;
        RECT 230.100 633.600 231.600 633.900 ;
        RECT 227.100 627.000 228.900 633.000 ;
        RECT 230.100 627.600 231.900 633.600 ;
        RECT 233.100 627.000 234.900 633.600 ;
        RECT 251.400 627.000 253.200 639.600 ;
        RECT 256.500 638.100 258.900 639.600 ;
        RECT 256.500 627.600 258.300 638.100 ;
        RECT 259.200 635.100 261.000 636.900 ;
        RECT 259.500 627.000 261.300 633.600 ;
        RECT 278.400 627.000 280.200 639.600 ;
        RECT 283.500 638.100 285.900 639.600 ;
        RECT 283.500 627.600 285.300 638.100 ;
        RECT 286.200 635.100 288.000 636.900 ;
        RECT 286.500 627.000 288.300 633.600 ;
        RECT 305.100 627.600 306.900 639.600 ;
        RECT 308.100 638.700 315.900 639.600 ;
        RECT 308.100 627.600 309.900 638.700 ;
        RECT 311.100 627.000 312.900 637.800 ;
        RECT 314.100 627.600 315.900 638.700 ;
        RECT 341.100 634.800 342.000 646.950 ;
        RECT 359.250 645.150 361.050 646.950 ;
        RECT 362.400 639.600 363.300 646.950 ;
        RECT 365.100 645.150 366.900 646.950 ;
        RECT 335.400 633.900 342.000 634.800 ;
        RECT 335.400 633.600 336.900 633.900 ;
        RECT 332.100 627.000 333.900 633.600 ;
        RECT 335.100 627.600 336.900 633.600 ;
        RECT 341.100 633.600 342.000 633.900 ;
        RECT 338.100 627.000 339.900 633.000 ;
        RECT 341.100 627.600 342.900 633.600 ;
        RECT 359.100 627.000 360.900 639.600 ;
        RECT 362.400 638.400 366.000 639.600 ;
        RECT 364.200 627.600 366.000 638.400 ;
        RECT 386.100 633.600 387.300 646.950 ;
        RECT 410.100 633.600 411.300 646.950 ;
        RECT 431.100 645.150 432.900 646.950 ;
        RECT 434.700 639.600 435.600 646.950 ;
        RECT 436.950 645.150 438.750 646.950 ;
        RECT 432.000 638.400 435.600 639.600 ;
        RECT 383.100 627.000 384.900 633.600 ;
        RECT 386.100 627.600 387.900 633.600 ;
        RECT 389.100 627.000 390.900 633.600 ;
        RECT 407.100 627.000 408.900 633.600 ;
        RECT 410.100 627.600 411.900 633.600 ;
        RECT 413.100 627.000 414.900 633.600 ;
        RECT 432.000 627.600 433.800 638.400 ;
        RECT 437.100 627.000 438.900 639.600 ;
        RECT 458.100 633.600 459.300 646.950 ;
        RECT 482.100 633.600 483.300 646.950 ;
        RECT 506.250 645.150 508.050 646.950 ;
        RECT 512.700 639.600 513.600 646.950 ;
        RECT 530.100 645.150 531.900 646.950 ;
        RECT 533.700 639.600 534.600 646.950 ;
        RECT 535.950 645.150 537.750 646.950 ;
        RECT 554.100 645.150 555.900 646.950 ;
        RECT 503.100 638.700 510.900 639.600 ;
        RECT 455.100 627.000 456.900 633.600 ;
        RECT 458.100 627.600 459.900 633.600 ;
        RECT 461.100 627.000 462.900 633.600 ;
        RECT 479.100 627.000 480.900 633.600 ;
        RECT 482.100 627.600 483.900 633.600 ;
        RECT 485.100 627.000 486.900 633.600 ;
        RECT 503.100 627.600 504.900 638.700 ;
        RECT 506.100 627.000 507.900 637.800 ;
        RECT 509.100 627.600 510.900 638.700 ;
        RECT 512.100 627.600 513.900 639.600 ;
        RECT 531.000 638.400 534.600 639.600 ;
        RECT 531.000 627.600 532.800 638.400 ;
        RECT 536.100 627.000 537.900 639.600 ;
        RECT 557.100 633.600 558.300 646.950 ;
        RECT 578.700 633.600 579.900 646.950 ;
        RECT 602.700 633.600 603.900 646.950 ;
        RECT 624.000 634.800 624.900 646.950 ;
        RECT 629.100 645.150 630.900 646.950 ;
        RECT 653.250 645.150 655.050 646.950 ;
        RECT 659.700 639.600 660.600 646.950 ;
        RECT 677.100 645.150 678.900 646.950 ;
        RECT 680.700 639.600 681.600 646.950 ;
        RECT 682.950 645.150 684.750 646.950 ;
        RECT 694.950 642.450 697.050 643.050 ;
        RECT 700.950 642.450 703.050 643.050 ;
        RECT 694.950 641.550 703.050 642.450 ;
        RECT 694.950 640.950 697.050 641.550 ;
        RECT 700.950 640.950 703.050 641.550 ;
        RECT 650.100 638.700 657.900 639.600 ;
        RECT 624.000 633.900 630.600 634.800 ;
        RECT 624.000 633.600 624.900 633.900 ;
        RECT 554.100 627.000 555.900 633.600 ;
        RECT 557.100 627.600 558.900 633.600 ;
        RECT 575.100 627.000 576.900 633.600 ;
        RECT 578.100 627.600 579.900 633.600 ;
        RECT 581.100 627.000 582.900 633.600 ;
        RECT 599.100 627.000 600.900 633.600 ;
        RECT 602.100 627.600 603.900 633.600 ;
        RECT 605.100 627.000 606.900 633.600 ;
        RECT 623.100 627.600 624.900 633.600 ;
        RECT 629.100 633.600 630.600 633.900 ;
        RECT 626.100 627.000 627.900 633.000 ;
        RECT 629.100 627.600 630.900 633.600 ;
        RECT 632.100 627.000 633.900 633.600 ;
        RECT 650.100 627.600 651.900 638.700 ;
        RECT 653.100 627.000 654.900 637.800 ;
        RECT 656.100 627.600 657.900 638.700 ;
        RECT 659.100 627.600 660.900 639.600 ;
        RECT 678.000 638.400 681.600 639.600 ;
        RECT 678.000 627.600 679.800 638.400 ;
        RECT 683.100 627.000 684.900 639.600 ;
        RECT 704.700 633.600 705.900 646.950 ;
        RECT 728.100 645.150 729.900 646.950 ;
        RECT 706.950 642.450 709.050 643.050 ;
        RECT 724.950 642.450 727.050 642.750 ;
        RECT 706.950 641.550 727.050 642.450 ;
        RECT 706.950 640.950 709.050 641.550 ;
        RECT 724.950 640.650 727.050 641.550 ;
        RECT 732.000 641.400 732.900 646.950 ;
        RECT 733.950 645.150 735.750 646.950 ;
        RECT 755.250 645.150 757.050 646.950 ;
        RECT 728.100 640.500 732.900 641.400 ;
        RECT 736.950 642.450 739.050 643.050 ;
        RECT 757.950 642.450 760.050 643.050 ;
        RECT 736.950 641.550 760.050 642.450 ;
        RECT 736.950 640.950 739.050 641.550 ;
        RECT 757.950 640.950 760.050 641.550 ;
        RECT 712.950 639.450 715.050 640.050 ;
        RECT 721.950 639.450 724.050 640.050 ;
        RECT 712.950 638.550 724.050 639.450 ;
        RECT 712.950 637.950 715.050 638.550 ;
        RECT 721.950 637.950 724.050 638.550 ;
        RECT 701.100 627.000 702.900 633.600 ;
        RECT 704.100 627.600 705.900 633.600 ;
        RECT 707.100 627.000 708.900 633.600 ;
        RECT 725.100 628.500 726.900 639.600 ;
        RECT 728.100 629.400 729.900 640.500 ;
        RECT 762.000 639.600 763.050 646.950 ;
        RECT 767.100 645.150 768.900 646.950 ;
        RECT 788.100 645.150 789.900 646.950 ;
        RECT 766.950 642.450 769.050 643.050 ;
        RECT 784.950 642.450 787.050 642.750 ;
        RECT 766.950 641.550 787.050 642.450 ;
        RECT 766.950 640.950 769.050 641.550 ;
        RECT 784.950 640.650 787.050 641.550 ;
        RECT 792.000 641.400 792.900 646.950 ;
        RECT 793.950 645.150 795.750 646.950 ;
        RECT 799.950 645.450 802.050 646.050 ;
        RECT 809.550 645.450 810.450 649.950 ;
        RECT 818.400 649.050 819.300 659.400 ;
        RECT 842.700 657.600 844.500 662.400 ;
        RECT 839.400 656.400 844.500 657.600 ;
        RECT 847.200 656.400 849.000 663.000 ;
        RECT 866.700 659.400 868.500 663.000 ;
        RECT 820.950 654.450 823.050 655.050 ;
        RECT 832.950 654.450 835.050 655.050 ;
        RECT 820.950 653.550 835.050 654.450 ;
        RECT 820.950 652.950 823.050 653.550 ;
        RECT 832.950 652.950 835.050 653.550 ;
        RECT 823.950 651.450 828.000 652.050 ;
        RECT 823.950 649.950 828.450 651.450 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 827.550 648.450 828.450 649.950 ;
        RECT 839.400 649.050 840.300 656.400 ;
        RECT 844.950 654.450 847.050 655.050 ;
        RECT 856.950 654.450 859.050 658.050 ;
        RECT 869.700 657.600 871.500 662.400 ;
        RECT 844.950 654.000 859.050 654.450 ;
        RECT 866.400 656.400 871.500 657.600 ;
        RECT 874.200 656.400 876.000 663.000 ;
        RECT 880.950 657.450 883.050 658.050 ;
        RECT 886.950 657.450 889.050 658.050 ;
        RECT 880.950 656.550 889.050 657.450 ;
        RECT 844.950 653.550 858.450 654.000 ;
        RECT 844.950 652.950 847.050 653.550 ;
        RECT 850.950 651.450 855.000 652.050 ;
        RECT 841.950 649.050 843.750 650.850 ;
        RECT 848.100 649.050 849.900 650.850 ;
        RECT 850.950 649.950 855.450 651.450 ;
        RECT 827.550 647.550 834.450 648.450 ;
        RECT 799.950 644.550 810.450 645.450 ;
        RECT 815.250 645.150 817.050 646.950 ;
        RECT 799.950 643.950 802.050 644.550 ;
        RECT 788.100 640.500 792.900 641.400 ;
        RECT 731.100 638.400 738.900 639.300 ;
        RECT 731.100 628.500 732.900 638.400 ;
        RECT 725.100 627.600 732.900 628.500 ;
        RECT 734.100 627.000 735.900 637.500 ;
        RECT 737.100 627.600 738.900 638.400 ;
        RECT 756.600 627.000 758.400 639.600 ;
        RECT 761.100 627.600 764.400 639.600 ;
        RECT 767.100 627.000 768.900 639.600 ;
        RECT 769.950 630.450 772.050 630.900 ;
        RECT 781.950 630.450 784.050 631.050 ;
        RECT 769.950 629.550 784.050 630.450 ;
        RECT 769.950 628.800 772.050 629.550 ;
        RECT 781.950 628.950 784.050 629.550 ;
        RECT 785.100 628.500 786.900 639.600 ;
        RECT 788.100 629.400 789.900 640.500 ;
        RECT 818.400 639.600 819.300 646.950 ;
        RECT 821.100 645.150 822.900 646.950 ;
        RECT 833.550 646.050 834.450 647.550 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 833.550 644.550 838.050 646.050 ;
        RECT 834.000 643.950 838.050 644.550 ;
        RECT 839.400 639.600 840.300 646.950 ;
        RECT 844.950 645.150 846.750 646.950 ;
        RECT 854.550 646.050 855.450 649.950 ;
        RECT 866.400 649.050 867.300 656.400 ;
        RECT 880.950 655.950 883.050 656.550 ;
        RECT 886.950 655.950 889.050 656.550 ;
        RECT 893.400 656.400 895.200 663.000 ;
        RECT 898.500 655.200 900.300 662.400 ;
        RECT 917.100 659.400 918.900 663.000 ;
        RECT 920.100 659.400 921.900 662.400 ;
        RECT 923.100 659.400 924.900 663.000 ;
        RECT 868.950 654.450 871.050 655.050 ;
        RECT 868.950 653.550 879.450 654.450 ;
        RECT 868.950 652.950 871.050 653.550 ;
        RECT 878.550 651.450 879.450 653.550 ;
        RECT 896.100 654.300 900.300 655.200 ;
        RECT 915.000 654.450 919.050 655.050 ;
        RECT 868.950 649.050 870.750 650.850 ;
        RECT 875.100 649.050 876.900 650.850 ;
        RECT 878.550 650.550 882.450 651.450 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 874.950 646.950 877.050 649.050 ;
        RECT 850.950 644.550 855.450 646.050 ;
        RECT 850.950 643.950 855.000 644.550 ;
        RECT 866.400 639.600 867.300 646.950 ;
        RECT 871.950 645.150 873.750 646.950 ;
        RECT 881.550 645.450 882.450 650.550 ;
        RECT 893.250 649.050 895.050 650.850 ;
        RECT 896.100 649.050 897.300 654.300 ;
        RECT 914.550 652.950 919.050 654.450 ;
        RECT 914.550 651.450 915.450 652.950 ;
        RECT 899.100 649.050 900.900 650.850 ;
        RECT 911.550 650.550 915.450 651.450 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 898.950 646.950 901.050 649.050 ;
        RECT 889.950 645.450 892.050 646.050 ;
        RECT 881.550 644.550 892.050 645.450 ;
        RECT 889.950 643.950 892.050 644.550 ;
        RECT 868.950 642.450 871.050 643.050 ;
        RECT 883.950 642.450 886.050 643.050 ;
        RECT 868.950 641.550 886.050 642.450 ;
        RECT 868.950 640.950 871.050 641.550 ;
        RECT 883.950 640.950 886.050 641.550 ;
        RECT 791.100 638.400 798.900 639.300 ;
        RECT 791.100 628.500 792.900 638.400 ;
        RECT 785.100 627.600 792.900 628.500 ;
        RECT 794.100 627.000 795.900 637.500 ;
        RECT 797.100 627.600 798.900 638.400 ;
        RECT 815.100 627.000 816.900 639.600 ;
        RECT 818.400 638.400 822.000 639.600 ;
        RECT 820.200 627.600 822.000 638.400 ;
        RECT 839.100 627.600 840.900 639.600 ;
        RECT 842.100 638.700 849.900 639.600 ;
        RECT 842.100 627.600 843.900 638.700 ;
        RECT 845.100 627.000 846.900 637.800 ;
        RECT 848.100 627.600 849.900 638.700 ;
        RECT 866.100 627.600 867.900 639.600 ;
        RECT 869.100 638.700 876.900 639.600 ;
        RECT 869.100 627.600 870.900 638.700 ;
        RECT 872.100 627.000 873.900 637.800 ;
        RECT 875.100 627.600 876.900 638.700 ;
        RECT 877.950 633.450 880.050 634.050 ;
        RECT 883.950 633.450 886.050 634.050 ;
        RECT 896.100 633.600 897.300 646.950 ;
        RECT 901.950 645.450 904.050 646.050 ;
        RECT 911.550 645.450 912.450 650.550 ;
        RECT 920.700 649.050 921.600 659.400 ;
        RECT 941.700 655.200 943.500 662.400 ;
        RECT 946.800 656.400 948.600 663.000 ;
        RECT 965.100 659.400 966.900 663.000 ;
        RECT 968.100 659.400 969.900 662.400 ;
        RECT 971.100 659.400 972.900 663.000 ;
        RECT 989.100 659.400 990.900 663.000 ;
        RECT 992.100 659.400 993.900 662.400 ;
        RECT 995.100 659.400 996.900 663.000 ;
        RECT 922.950 654.450 925.050 655.050 ;
        RECT 931.950 654.450 934.050 655.050 ;
        RECT 922.950 653.550 934.050 654.450 ;
        RECT 941.700 654.300 945.900 655.200 ;
        RECT 964.950 654.450 967.050 655.050 ;
        RECT 922.950 652.950 925.050 653.550 ;
        RECT 931.950 652.950 934.050 653.550 ;
        RECT 941.100 649.050 942.900 650.850 ;
        RECT 944.700 649.050 945.900 654.300 ;
        RECT 953.550 653.550 967.050 654.450 ;
        RECT 946.950 649.050 948.750 650.850 ;
        RECT 916.950 646.950 919.050 649.050 ;
        RECT 919.950 646.950 922.050 649.050 ;
        RECT 922.950 646.950 925.050 649.050 ;
        RECT 940.950 646.950 943.050 649.050 ;
        RECT 943.950 646.950 946.050 649.050 ;
        RECT 946.950 646.950 949.050 649.050 ;
        RECT 901.950 644.550 912.450 645.450 ;
        RECT 917.100 645.150 918.900 646.950 ;
        RECT 901.950 643.950 904.050 644.550 ;
        RECT 920.700 639.600 921.600 646.950 ;
        RECT 922.950 645.150 924.750 646.950 ;
        RECT 925.950 645.450 928.050 646.050 ;
        RECT 931.950 645.450 934.050 646.050 ;
        RECT 925.950 644.550 934.050 645.450 ;
        RECT 925.950 643.950 928.050 644.550 ;
        RECT 931.950 643.950 934.050 644.550 ;
        RECT 922.950 642.450 925.050 643.050 ;
        RECT 940.950 642.450 943.050 643.050 ;
        RECT 922.950 641.550 943.050 642.450 ;
        RECT 922.950 640.950 925.050 641.550 ;
        RECT 940.950 640.950 943.050 641.550 ;
        RECT 918.000 638.400 921.600 639.600 ;
        RECT 898.950 636.450 901.050 637.050 ;
        RECT 910.950 636.450 913.050 637.050 ;
        RECT 898.950 635.550 913.050 636.450 ;
        RECT 898.950 634.950 901.050 635.550 ;
        RECT 910.950 634.950 913.050 635.550 ;
        RECT 877.950 632.550 886.050 633.450 ;
        RECT 877.950 631.950 880.050 632.550 ;
        RECT 883.950 631.950 886.050 632.550 ;
        RECT 893.100 627.000 894.900 633.600 ;
        RECT 896.100 627.600 897.900 633.600 ;
        RECT 899.100 627.000 900.900 633.600 ;
        RECT 918.000 627.600 919.800 638.400 ;
        RECT 923.100 627.000 924.900 639.600 ;
        RECT 925.950 639.450 928.050 640.050 ;
        RECT 940.950 639.450 943.050 639.900 ;
        RECT 925.950 638.550 943.050 639.450 ;
        RECT 925.950 637.950 928.050 638.550 ;
        RECT 940.950 637.800 943.050 638.550 ;
        RECT 944.700 633.600 945.900 646.950 ;
        RECT 953.550 645.450 954.450 653.550 ;
        RECT 964.950 652.950 967.050 653.550 ;
        RECT 960.000 651.450 964.050 652.050 ;
        RECT 950.550 644.550 954.450 645.450 ;
        RECT 959.550 649.950 964.050 651.450 ;
        RECT 950.550 642.450 951.450 644.550 ;
        RECT 959.550 643.050 960.450 649.950 ;
        RECT 968.400 649.050 969.300 659.400 ;
        RECT 973.950 651.450 978.000 652.050 ;
        RECT 979.950 651.450 984.000 652.050 ;
        RECT 973.950 649.950 978.450 651.450 ;
        RECT 979.950 649.950 984.450 651.450 ;
        RECT 977.550 649.050 978.450 649.950 ;
        RECT 964.950 646.950 967.050 649.050 ;
        RECT 967.950 646.950 970.050 649.050 ;
        RECT 970.950 646.950 973.050 649.050 ;
        RECT 977.550 648.900 981.000 649.050 ;
        RECT 977.550 647.550 982.050 648.900 ;
        RECT 978.000 646.950 982.050 647.550 ;
        RECT 965.250 645.150 967.050 646.950 ;
        RECT 947.550 642.000 951.450 642.450 ;
        RECT 946.950 641.550 951.450 642.000 ;
        RECT 952.950 642.450 955.050 642.900 ;
        RECT 959.550 642.450 964.050 643.050 ;
        RECT 952.950 641.550 964.050 642.450 ;
        RECT 946.950 637.800 949.050 641.550 ;
        RECT 952.950 640.800 955.050 641.550 ;
        RECT 960.000 640.950 964.050 641.550 ;
        RECT 968.400 639.600 969.300 646.950 ;
        RECT 971.100 645.150 972.900 646.950 ;
        RECT 979.950 646.800 982.050 646.950 ;
        RECT 983.550 646.050 984.450 649.950 ;
        RECT 992.400 649.050 993.300 659.400 ;
        RECT 1013.700 655.200 1015.500 662.400 ;
        RECT 1018.800 656.400 1020.600 663.000 ;
        RECT 1013.700 654.300 1017.900 655.200 ;
        RECT 1013.100 649.050 1014.900 650.850 ;
        RECT 1016.700 649.050 1017.900 654.300 ;
        RECT 1018.950 649.050 1020.750 650.850 ;
        RECT 988.950 646.950 991.050 649.050 ;
        RECT 991.950 646.950 994.050 649.050 ;
        RECT 994.950 646.950 997.050 649.050 ;
        RECT 1012.950 646.950 1015.050 649.050 ;
        RECT 1015.950 646.950 1018.050 649.050 ;
        RECT 1018.950 646.950 1021.050 649.050 ;
        RECT 983.550 644.550 988.050 646.050 ;
        RECT 989.250 645.150 991.050 646.950 ;
        RECT 984.000 643.950 988.050 644.550 ;
        RECT 970.950 642.450 973.050 643.050 ;
        RECT 988.950 642.450 991.050 643.050 ;
        RECT 970.950 641.550 991.050 642.450 ;
        RECT 970.950 640.950 973.050 641.550 ;
        RECT 988.950 640.950 991.050 641.550 ;
        RECT 992.400 639.600 993.300 646.950 ;
        RECT 995.100 645.150 996.900 646.950 ;
        RECT 997.950 645.450 1000.050 646.050 ;
        RECT 1006.950 645.450 1009.050 646.050 ;
        RECT 997.950 644.550 1009.050 645.450 ;
        RECT 997.950 643.950 1000.050 644.550 ;
        RECT 1006.950 643.950 1009.050 644.550 ;
        RECT 941.100 627.000 942.900 633.600 ;
        RECT 944.100 627.600 945.900 633.600 ;
        RECT 947.100 627.000 948.900 633.600 ;
        RECT 965.100 627.000 966.900 639.600 ;
        RECT 968.400 638.400 972.000 639.600 ;
        RECT 970.200 627.600 972.000 638.400 ;
        RECT 989.100 627.000 990.900 639.600 ;
        RECT 992.400 638.400 996.000 639.600 ;
        RECT 994.200 627.600 996.000 638.400 ;
        RECT 1016.700 633.600 1017.900 646.950 ;
        RECT 1013.100 627.000 1014.900 633.600 ;
        RECT 1016.100 627.600 1017.900 633.600 ;
        RECT 1019.100 627.000 1020.900 633.600 ;
        RECT 17.100 611.400 18.900 623.400 ;
        RECT 20.100 613.200 21.900 624.000 ;
        RECT 23.100 617.400 24.900 623.400 ;
        RECT 41.700 617.400 43.500 624.000 ;
        RECT 17.100 604.050 18.300 611.400 ;
        RECT 23.700 610.500 24.900 617.400 ;
        RECT 42.000 614.100 43.800 615.900 ;
        RECT 44.700 612.900 46.500 623.400 ;
        RECT 19.200 609.600 24.900 610.500 ;
        RECT 44.100 611.400 46.500 612.900 ;
        RECT 49.800 611.400 51.600 624.000 ;
        RECT 53.700 617.400 55.500 624.000 ;
        RECT 56.700 618.300 58.500 623.400 ;
        RECT 56.400 617.400 58.500 618.300 ;
        RECT 59.700 617.400 61.500 624.000 ;
        RECT 56.400 616.500 57.300 617.400 ;
        RECT 53.700 615.600 57.300 616.500 ;
        RECT 19.200 608.700 21.000 609.600 ;
        RECT 17.100 601.950 19.200 604.050 ;
        RECT 17.100 594.600 18.300 601.950 ;
        RECT 20.100 597.300 21.000 608.700 ;
        RECT 31.950 609.450 34.050 610.050 ;
        RECT 40.950 609.450 43.050 610.200 ;
        RECT 31.950 608.550 43.050 609.450 ;
        RECT 31.950 607.950 34.050 608.550 ;
        RECT 40.950 608.100 43.050 608.550 ;
        RECT 22.800 604.050 24.600 605.850 ;
        RECT 44.100 604.050 45.300 611.400 ;
        RECT 50.100 604.050 51.900 605.850 ;
        RECT 22.500 601.950 24.600 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 46.950 601.950 49.050 604.050 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 41.100 600.150 42.900 601.950 ;
        RECT 19.200 596.400 21.000 597.300 ;
        RECT 25.950 597.450 28.050 598.050 ;
        RECT 31.950 597.450 34.050 598.050 ;
        RECT 44.100 597.600 45.300 601.950 ;
        RECT 47.100 600.150 48.900 601.950 ;
        RECT 25.950 596.550 34.050 597.450 ;
        RECT 19.200 595.500 24.900 596.400 ;
        RECT 25.950 595.950 28.050 596.550 ;
        RECT 31.950 595.950 34.050 596.550 ;
        RECT 41.700 596.700 45.300 597.600 ;
        RECT 53.700 599.400 54.900 615.600 ;
        RECT 58.200 614.400 60.000 614.700 ;
        RECT 62.700 614.400 64.500 623.400 ;
        RECT 65.700 617.400 67.500 624.000 ;
        RECT 69.300 620.400 71.100 623.400 ;
        RECT 72.300 620.400 74.100 623.400 ;
        RECT 69.300 618.300 71.400 620.400 ;
        RECT 72.300 618.300 74.400 620.400 ;
        RECT 75.300 617.400 77.100 623.400 ;
        RECT 78.300 617.400 80.100 624.000 ;
        RECT 74.700 615.300 76.800 617.400 ;
        RECT 82.200 615.900 84.000 623.400 ;
        RECT 85.200 617.400 87.000 624.000 ;
        RECT 88.200 617.400 90.000 623.400 ;
        RECT 91.200 620.400 93.000 623.400 ;
        RECT 94.200 620.400 96.000 623.400 ;
        RECT 97.200 620.400 99.000 623.400 ;
        RECT 91.200 618.300 93.300 620.400 ;
        RECT 94.200 618.300 96.300 620.400 ;
        RECT 97.200 618.300 99.300 620.400 ;
        RECT 100.200 617.400 102.000 624.000 ;
        RECT 103.200 617.400 105.000 623.400 ;
        RECT 106.200 617.400 108.000 624.000 ;
        RECT 109.200 617.400 111.000 623.400 ;
        RECT 112.200 617.400 114.000 624.000 ;
        RECT 115.500 617.400 117.300 623.400 ;
        RECT 118.500 617.400 120.300 624.000 ;
        RECT 137.700 617.400 139.500 624.000 ;
        RECT 58.200 613.200 77.400 614.400 ;
        RECT 82.200 613.800 85.500 615.900 ;
        RECT 88.200 613.500 90.900 617.400 ;
        RECT 94.200 616.500 96.300 617.400 ;
        RECT 94.200 615.300 102.300 616.500 ;
        RECT 100.500 614.700 102.300 615.300 ;
        RECT 103.200 614.400 104.400 617.400 ;
        RECT 109.800 616.500 111.000 617.400 ;
        RECT 109.800 615.600 113.700 616.500 ;
        RECT 107.100 614.400 108.900 615.000 ;
        RECT 58.200 612.900 60.000 613.200 ;
        RECT 76.200 612.600 77.400 613.200 ;
        RECT 91.800 612.600 93.900 613.500 ;
        RECT 61.500 611.700 63.300 612.300 ;
        RECT 71.400 611.700 73.500 612.300 ;
        RECT 61.500 610.500 73.500 611.700 ;
        RECT 76.200 611.400 93.900 612.600 ;
        RECT 97.200 612.300 99.300 613.500 ;
        RECT 103.200 613.200 108.900 614.400 ;
        RECT 112.800 612.300 113.700 615.600 ;
        RECT 97.200 611.400 113.700 612.300 ;
        RECT 71.400 610.200 73.500 610.500 ;
        RECT 76.200 609.300 111.900 610.500 ;
        RECT 76.200 608.700 77.400 609.300 ;
        RECT 110.100 608.700 111.900 609.300 ;
        RECT 63.900 607.800 77.400 608.700 ;
        RECT 88.800 607.800 90.900 608.100 ;
        RECT 63.900 607.050 65.700 607.800 ;
        RECT 55.800 604.950 57.900 607.050 ;
        RECT 61.800 605.250 65.700 607.050 ;
        RECT 83.400 606.300 85.500 607.200 ;
        RECT 61.800 604.950 63.900 605.250 ;
        RECT 74.400 605.100 85.500 606.300 ;
        RECT 87.000 606.000 90.900 607.800 ;
        RECT 95.100 606.300 96.900 608.100 ;
        RECT 96.000 605.100 96.900 606.300 ;
        RECT 56.100 603.300 57.900 604.950 ;
        RECT 74.400 604.500 76.200 605.100 ;
        RECT 83.400 604.200 96.900 605.100 ;
        RECT 99.600 604.800 104.700 606.600 ;
        RECT 106.800 604.950 108.900 607.050 ;
        RECT 99.600 603.300 100.500 604.800 ;
        RECT 56.100 602.100 100.500 603.300 ;
        RECT 106.800 602.100 108.300 604.950 ;
        RECT 71.400 599.400 73.200 601.200 ;
        RECT 79.800 600.000 81.900 601.050 ;
        RECT 101.700 600.600 108.300 602.100 ;
        RECT 53.700 598.200 70.500 599.400 ;
        RECT 17.100 588.600 18.900 594.600 ;
        RECT 20.100 588.000 21.900 594.600 ;
        RECT 23.700 591.600 24.900 595.500 ;
        RECT 41.700 594.600 42.900 596.700 ;
        RECT 23.100 588.600 24.900 591.600 ;
        RECT 41.100 588.600 42.900 594.600 ;
        RECT 44.100 593.700 51.900 595.050 ;
        RECT 44.100 588.600 45.900 593.700 ;
        RECT 47.100 588.000 48.900 592.800 ;
        RECT 50.100 588.600 51.900 593.700 ;
        RECT 53.700 594.600 54.900 598.200 ;
        RECT 68.400 597.300 70.500 598.200 ;
        RECT 57.900 596.700 59.700 597.300 ;
        RECT 57.900 595.500 66.300 596.700 ;
        RECT 64.800 594.600 66.300 595.500 ;
        RECT 71.400 596.400 72.300 599.400 ;
        RECT 76.800 599.100 81.900 600.000 ;
        RECT 76.800 598.200 78.600 599.100 ;
        RECT 79.800 598.950 81.900 599.100 ;
        RECT 86.100 599.100 103.200 600.600 ;
        RECT 86.100 598.500 88.200 599.100 ;
        RECT 86.100 596.700 87.900 598.500 ;
        RECT 104.100 597.900 111.900 599.700 ;
        RECT 71.400 595.200 78.600 596.400 ;
        RECT 73.800 594.600 75.600 595.200 ;
        RECT 77.700 594.600 78.600 595.200 ;
        RECT 93.300 594.600 99.900 596.400 ;
        RECT 104.100 594.600 105.600 597.900 ;
        RECT 112.800 594.600 113.700 611.400 ;
        RECT 53.700 588.600 55.500 594.600 ;
        RECT 59.100 588.000 60.900 594.600 ;
        RECT 64.500 588.600 66.300 594.600 ;
        RECT 68.700 591.600 70.800 593.700 ;
        RECT 71.700 591.600 73.800 593.700 ;
        RECT 74.700 591.600 76.800 593.700 ;
        RECT 77.700 593.400 80.400 594.600 ;
        RECT 78.600 592.500 80.400 593.400 ;
        RECT 82.200 592.500 84.900 594.600 ;
        RECT 68.700 588.600 70.500 591.600 ;
        RECT 71.700 588.600 73.500 591.600 ;
        RECT 74.700 588.600 76.500 591.600 ;
        RECT 77.700 588.000 79.500 591.600 ;
        RECT 82.200 588.600 84.000 592.500 ;
        RECT 88.200 591.600 90.300 593.700 ;
        RECT 91.200 591.600 93.300 593.700 ;
        RECT 94.200 591.600 96.300 593.700 ;
        RECT 97.200 591.600 99.300 593.700 ;
        RECT 101.400 593.400 105.600 594.600 ;
        RECT 85.200 588.000 87.000 591.600 ;
        RECT 88.200 588.600 90.000 591.600 ;
        RECT 91.200 588.600 93.000 591.600 ;
        RECT 94.200 588.600 96.000 591.600 ;
        RECT 97.200 588.600 99.000 591.600 ;
        RECT 101.400 588.600 103.200 593.400 ;
        RECT 106.500 588.000 108.300 594.600 ;
        RECT 111.900 588.600 113.700 594.600 ;
        RECT 115.500 607.050 117.000 617.400 ;
        RECT 138.000 614.100 139.800 615.900 ;
        RECT 140.700 612.900 142.500 623.400 ;
        RECT 140.100 611.400 142.500 612.900 ;
        RECT 145.800 611.400 147.600 624.000 ;
        RECT 164.100 612.300 165.900 623.400 ;
        RECT 167.100 613.200 168.900 624.000 ;
        RECT 170.100 612.300 171.900 623.400 ;
        RECT 164.100 611.400 171.900 612.300 ;
        RECT 173.100 611.400 174.900 623.400 ;
        RECT 191.100 617.400 192.900 624.000 ;
        RECT 194.100 617.400 195.900 623.400 ;
        RECT 115.500 604.950 117.900 607.050 ;
        RECT 115.500 591.600 117.000 604.950 ;
        RECT 140.100 604.050 141.300 611.400 ;
        RECT 154.950 609.450 157.050 610.050 ;
        RECT 169.950 609.450 172.050 610.050 ;
        RECT 154.950 608.550 172.050 609.450 ;
        RECT 154.950 607.950 157.050 608.550 ;
        RECT 169.950 607.950 172.050 608.550 ;
        RECT 146.100 604.050 147.900 605.850 ;
        RECT 167.250 604.050 169.050 605.850 ;
        RECT 173.700 604.050 174.600 611.400 ;
        RECT 191.100 604.050 192.900 605.850 ;
        RECT 194.100 604.050 195.300 617.400 ;
        RECT 212.100 611.400 213.900 623.400 ;
        RECT 215.100 612.300 216.900 623.400 ;
        RECT 218.100 613.200 219.900 624.000 ;
        RECT 221.100 612.300 222.900 623.400 ;
        RECT 215.100 611.400 222.900 612.300 ;
        RECT 239.100 611.400 240.900 624.000 ;
        RECT 244.200 612.600 246.000 623.400 ;
        RECT 242.400 611.400 246.000 612.600 ;
        RECT 263.100 612.300 264.900 623.400 ;
        RECT 266.100 613.200 267.900 624.000 ;
        RECT 269.100 612.300 270.900 623.400 ;
        RECT 263.100 611.400 270.900 612.300 ;
        RECT 272.100 611.400 273.900 623.400 ;
        RECT 290.100 617.400 291.900 624.000 ;
        RECT 293.100 617.400 294.900 623.400 ;
        RECT 296.100 618.000 297.900 624.000 ;
        RECT 293.400 617.100 294.900 617.400 ;
        RECT 299.100 617.400 300.900 623.400 ;
        RECT 317.100 617.400 318.900 623.400 ;
        RECT 320.100 618.000 321.900 624.000 ;
        RECT 299.100 617.100 300.000 617.400 ;
        RECT 293.400 616.200 300.000 617.100 ;
        RECT 212.400 604.050 213.300 611.400 ;
        RECT 229.950 609.450 232.050 610.050 ;
        RECT 238.950 609.450 241.050 610.050 ;
        RECT 229.950 608.550 241.050 609.450 ;
        RECT 229.950 607.950 232.050 608.550 ;
        RECT 238.950 607.950 241.050 608.550 ;
        RECT 217.950 604.050 219.750 605.850 ;
        RECT 239.250 604.050 241.050 605.850 ;
        RECT 242.400 604.050 243.300 611.400 ;
        RECT 256.950 609.450 259.050 610.050 ;
        RECT 268.950 609.450 271.050 610.200 ;
        RECT 256.950 608.550 271.050 609.450 ;
        RECT 256.950 607.950 259.050 608.550 ;
        RECT 268.950 608.100 271.050 608.550 ;
        RECT 245.100 604.050 246.900 605.850 ;
        RECT 266.250 604.050 268.050 605.850 ;
        RECT 272.700 604.050 273.600 611.400 ;
        RECT 293.100 604.050 294.900 605.850 ;
        RECT 299.100 604.050 300.000 616.200 ;
        RECT 318.000 617.100 318.900 617.400 ;
        RECT 323.100 617.400 324.900 623.400 ;
        RECT 326.100 617.400 327.900 624.000 ;
        RECT 323.100 617.100 324.600 617.400 ;
        RECT 318.000 616.200 324.600 617.100 ;
        RECT 318.000 604.050 318.900 616.200 ;
        RECT 345.000 612.600 346.800 623.400 ;
        RECT 345.000 611.400 348.600 612.600 ;
        RECT 350.100 611.400 351.900 624.000 ;
        RECT 368.100 617.400 369.900 624.000 ;
        RECT 371.100 617.400 372.900 623.400 ;
        RECT 323.100 604.050 324.900 605.850 ;
        RECT 344.100 604.050 345.900 605.850 ;
        RECT 347.700 604.050 348.600 611.400 ;
        RECT 352.950 606.450 355.050 607.050 ;
        RECT 358.950 606.450 361.050 607.050 ;
        RECT 349.950 604.050 351.750 605.850 ;
        RECT 352.950 605.550 361.050 606.450 ;
        RECT 352.950 604.950 355.050 605.550 ;
        RECT 358.950 604.950 361.050 605.550 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 368.100 601.950 370.200 604.050 ;
        RECT 137.100 600.150 138.900 601.950 ;
        RECT 140.100 597.600 141.300 601.950 ;
        RECT 143.100 600.150 144.900 601.950 ;
        RECT 164.100 600.150 165.900 601.950 ;
        RECT 170.250 600.150 172.050 601.950 ;
        RECT 137.700 596.700 141.300 597.600 ;
        RECT 137.700 594.600 138.900 596.700 ;
        RECT 115.500 588.600 117.300 591.600 ;
        RECT 118.500 588.000 120.300 591.600 ;
        RECT 137.100 588.600 138.900 594.600 ;
        RECT 140.100 593.700 147.900 595.050 ;
        RECT 173.700 594.600 174.600 601.950 ;
        RECT 140.100 588.600 141.900 593.700 ;
        RECT 143.100 588.000 144.900 592.800 ;
        RECT 146.100 588.600 147.900 593.700 ;
        RECT 165.000 588.000 166.800 594.600 ;
        RECT 169.500 593.400 174.600 594.600 ;
        RECT 169.500 588.600 171.300 593.400 ;
        RECT 194.100 591.600 195.300 601.950 ;
        RECT 212.400 594.600 213.300 601.950 ;
        RECT 214.950 600.150 216.750 601.950 ;
        RECT 221.100 600.150 222.900 601.950 ;
        RECT 217.950 597.450 220.050 598.050 ;
        RECT 235.950 597.450 238.050 598.050 ;
        RECT 217.950 596.550 238.050 597.450 ;
        RECT 217.950 595.950 220.050 596.550 ;
        RECT 235.950 595.950 238.050 596.550 ;
        RECT 212.400 593.400 217.500 594.600 ;
        RECT 172.500 588.000 174.300 591.600 ;
        RECT 191.100 588.000 192.900 591.600 ;
        RECT 194.100 588.600 195.900 591.600 ;
        RECT 212.700 588.000 214.500 591.600 ;
        RECT 215.700 588.600 217.500 593.400 ;
        RECT 220.200 588.000 222.000 594.600 ;
        RECT 242.400 591.600 243.300 601.950 ;
        RECT 263.100 600.150 264.900 601.950 ;
        RECT 269.250 600.150 271.050 601.950 ;
        RECT 272.700 594.600 273.600 601.950 ;
        RECT 290.100 600.150 291.900 601.950 ;
        RECT 296.100 600.150 297.900 601.950 ;
        RECT 299.100 598.200 300.000 601.950 ;
        RECT 239.100 588.000 240.900 591.600 ;
        RECT 242.100 588.600 243.900 591.600 ;
        RECT 245.100 588.000 246.900 591.600 ;
        RECT 264.000 588.000 265.800 594.600 ;
        RECT 268.500 593.400 273.600 594.600 ;
        RECT 268.500 588.600 270.300 593.400 ;
        RECT 271.500 588.000 273.300 591.600 ;
        RECT 290.100 588.000 291.900 597.600 ;
        RECT 296.700 597.000 300.000 598.200 ;
        RECT 318.000 598.200 318.900 601.950 ;
        RECT 320.100 600.150 321.900 601.950 ;
        RECT 326.100 600.150 327.900 601.950 ;
        RECT 318.000 597.000 321.300 598.200 ;
        RECT 296.700 588.600 298.500 597.000 ;
        RECT 319.500 588.600 321.300 597.000 ;
        RECT 326.100 588.000 327.900 597.600 ;
        RECT 347.700 591.600 348.600 601.950 ;
        RECT 368.250 600.150 370.050 601.950 ;
        RECT 371.100 597.300 372.000 617.400 ;
        RECT 374.100 612.000 375.900 624.000 ;
        RECT 377.100 611.400 378.900 623.400 ;
        RECT 392.100 617.400 393.900 623.400 ;
        RECT 395.100 618.000 396.900 624.000 ;
        RECT 393.000 617.100 393.900 617.400 ;
        RECT 398.100 617.400 399.900 623.400 ;
        RECT 401.100 617.400 402.900 624.000 ;
        RECT 419.100 617.400 420.900 624.000 ;
        RECT 422.100 617.400 423.900 623.400 ;
        RECT 425.100 618.000 426.900 624.000 ;
        RECT 398.100 617.100 399.600 617.400 ;
        RECT 393.000 616.200 399.600 617.100 ;
        RECT 422.400 617.100 423.900 617.400 ;
        RECT 428.100 617.400 429.900 623.400 ;
        RECT 446.100 617.400 447.900 624.000 ;
        RECT 449.100 617.400 450.900 623.400 ;
        RECT 467.700 617.400 469.500 624.000 ;
        RECT 428.100 617.100 429.000 617.400 ;
        RECT 422.400 616.200 429.000 617.100 ;
        RECT 373.200 604.050 375.000 605.850 ;
        RECT 377.400 604.050 378.300 611.400 ;
        RECT 393.000 604.050 393.900 616.200 ;
        RECT 412.950 612.450 415.050 613.050 ;
        RECT 421.950 612.450 424.050 613.050 ;
        RECT 412.950 611.550 424.050 612.450 ;
        RECT 412.950 610.950 415.050 611.550 ;
        RECT 421.950 610.950 424.050 611.550 ;
        RECT 400.950 609.450 403.050 610.050 ;
        RECT 424.950 609.450 427.050 610.050 ;
        RECT 400.950 608.550 427.050 609.450 ;
        RECT 400.950 607.950 403.050 608.550 ;
        RECT 424.950 607.950 427.050 608.550 ;
        RECT 398.100 604.050 399.900 605.850 ;
        RECT 422.100 604.050 423.900 605.850 ;
        RECT 428.100 604.050 429.000 616.200 ;
        RECT 446.100 604.050 447.900 605.850 ;
        RECT 449.100 604.050 450.300 617.400 ;
        RECT 468.000 614.100 469.800 615.900 ;
        RECT 470.700 612.900 472.500 623.400 ;
        RECT 470.100 611.400 472.500 612.900 ;
        RECT 475.800 611.400 477.600 624.000 ;
        RECT 494.100 617.400 495.900 624.000 ;
        RECT 497.100 617.400 498.900 623.400 ;
        RECT 500.100 617.400 501.900 624.000 ;
        RECT 470.100 604.050 471.300 611.400 ;
        RECT 476.100 604.050 477.900 605.850 ;
        RECT 497.100 604.050 498.300 617.400 ;
        RECT 518.100 611.400 519.900 624.000 ;
        RECT 523.200 612.600 525.000 623.400 ;
        RECT 542.100 617.400 543.900 624.000 ;
        RECT 545.100 617.400 546.900 623.400 ;
        RECT 548.100 617.400 549.900 624.000 ;
        RECT 566.100 617.400 567.900 624.000 ;
        RECT 569.100 617.400 570.900 623.400 ;
        RECT 572.100 617.400 573.900 624.000 ;
        RECT 590.100 622.500 597.900 623.400 ;
        RECT 521.400 611.400 525.000 612.600 ;
        RECT 518.250 604.050 520.050 605.850 ;
        RECT 521.400 604.050 522.300 611.400 ;
        RECT 523.950 609.450 526.050 610.050 ;
        RECT 541.950 609.450 544.050 609.900 ;
        RECT 523.950 608.550 544.050 609.450 ;
        RECT 523.950 607.950 526.050 608.550 ;
        RECT 541.950 607.800 544.050 608.550 ;
        RECT 524.100 604.050 525.900 605.850 ;
        RECT 545.700 604.050 546.900 617.400 ;
        RECT 569.100 604.050 570.300 617.400 ;
        RECT 590.100 611.400 591.900 622.500 ;
        RECT 593.100 610.500 594.900 621.600 ;
        RECT 596.100 612.600 597.900 622.500 ;
        RECT 599.100 613.500 600.900 624.000 ;
        RECT 602.100 612.600 603.900 623.400 ;
        RECT 596.100 611.700 603.900 612.600 ;
        RECT 620.100 611.400 621.900 624.000 ;
        RECT 623.100 611.400 624.900 623.400 ;
        RECT 641.100 611.400 642.900 624.000 ;
        RECT 646.200 612.600 648.000 623.400 ;
        RECT 644.400 611.400 648.000 612.600 ;
        RECT 665.100 612.600 666.900 623.400 ;
        RECT 668.100 613.500 669.900 624.000 ;
        RECT 671.100 622.500 678.900 623.400 ;
        RECT 671.100 612.600 672.900 622.500 ;
        RECT 665.100 611.700 672.900 612.600 ;
        RECT 593.100 609.600 597.900 610.500 ;
        RECT 593.100 604.050 594.900 605.850 ;
        RECT 597.000 604.050 597.900 609.600 ;
        RECT 598.950 604.050 600.750 605.850 ;
        RECT 623.100 604.050 624.300 611.400 ;
        RECT 641.250 604.050 643.050 605.850 ;
        RECT 644.400 604.050 645.300 611.400 ;
        RECT 674.100 610.500 675.900 621.600 ;
        RECT 677.100 611.400 678.900 622.500 ;
        RECT 696.600 611.400 698.400 624.000 ;
        RECT 701.100 611.400 704.400 623.400 ;
        RECT 707.100 611.400 708.900 624.000 ;
        RECT 725.100 612.600 726.900 623.400 ;
        RECT 728.100 613.500 729.900 624.000 ;
        RECT 731.100 622.500 738.900 623.400 ;
        RECT 731.100 612.600 732.900 622.500 ;
        RECT 725.100 611.700 732.900 612.600 ;
        RECT 671.100 609.600 675.900 610.500 ;
        RECT 647.100 604.050 648.900 605.850 ;
        RECT 668.250 604.050 670.050 605.850 ;
        RECT 671.100 604.050 672.000 609.600 ;
        RECT 679.950 606.450 684.000 607.050 ;
        RECT 679.950 606.000 684.450 606.450 ;
        RECT 674.100 604.050 675.900 605.850 ;
        RECT 679.950 604.950 685.050 606.000 ;
        RECT 373.500 601.950 375.600 604.050 ;
        RECT 376.800 601.950 378.900 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 418.950 601.950 421.050 604.050 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 496.950 601.950 499.050 604.050 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 520.950 601.950 523.050 604.050 ;
        RECT 523.950 601.950 526.050 604.050 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 571.950 601.950 574.050 604.050 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 682.950 601.950 685.050 604.950 ;
        RECT 695.250 604.050 697.050 605.850 ;
        RECT 702.000 604.050 703.050 611.400 ;
        RECT 734.100 610.500 735.900 621.600 ;
        RECT 737.100 611.400 738.900 622.500 ;
        RECT 755.100 611.400 756.900 623.400 ;
        RECT 758.100 612.300 759.900 623.400 ;
        RECT 761.100 613.200 762.900 624.000 ;
        RECT 764.100 612.300 765.900 623.400 ;
        RECT 783.600 612.900 785.400 623.400 ;
        RECT 758.100 611.400 765.900 612.300 ;
        RECT 783.000 611.400 785.400 612.900 ;
        RECT 786.600 611.400 788.400 624.000 ;
        RECT 791.100 611.400 792.900 623.400 ;
        RECT 809.100 617.400 810.900 624.000 ;
        RECT 812.100 617.400 813.900 623.400 ;
        RECT 815.100 617.400 816.900 624.000 ;
        RECT 706.950 609.450 709.050 610.050 ;
        RECT 712.950 609.450 715.050 610.050 ;
        RECT 727.950 609.450 730.050 610.050 ;
        RECT 706.950 608.550 715.050 609.450 ;
        RECT 706.950 607.950 709.050 608.550 ;
        RECT 712.950 607.950 715.050 608.550 ;
        RECT 719.550 608.550 730.050 609.450 ;
        RECT 707.100 604.050 708.900 605.850 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 697.950 601.950 700.050 604.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 368.100 596.400 376.500 597.300 ;
        RECT 344.100 588.000 345.900 591.600 ;
        RECT 347.100 588.600 348.900 591.600 ;
        RECT 350.100 588.000 351.900 591.600 ;
        RECT 368.100 588.600 369.900 596.400 ;
        RECT 374.700 595.500 376.500 596.400 ;
        RECT 377.400 594.600 378.300 601.950 ;
        RECT 393.000 598.200 393.900 601.950 ;
        RECT 395.100 600.150 396.900 601.950 ;
        RECT 401.100 600.150 402.900 601.950 ;
        RECT 419.100 600.150 420.900 601.950 ;
        RECT 425.100 600.150 426.900 601.950 ;
        RECT 428.100 598.200 429.000 601.950 ;
        RECT 393.000 597.000 396.300 598.200 ;
        RECT 372.600 588.000 374.400 594.600 ;
        RECT 375.600 592.800 378.300 594.600 ;
        RECT 375.600 588.600 377.400 592.800 ;
        RECT 394.500 588.600 396.300 597.000 ;
        RECT 401.100 588.000 402.900 597.600 ;
        RECT 419.100 588.000 420.900 597.600 ;
        RECT 425.700 597.000 429.000 598.200 ;
        RECT 425.700 588.600 427.500 597.000 ;
        RECT 449.100 591.600 450.300 601.950 ;
        RECT 467.100 600.150 468.900 601.950 ;
        RECT 470.100 597.600 471.300 601.950 ;
        RECT 473.100 600.150 474.900 601.950 ;
        RECT 494.250 600.150 496.050 601.950 ;
        RECT 467.700 596.700 471.300 597.600 ;
        RECT 497.100 596.700 498.300 601.950 ;
        RECT 500.100 600.150 501.900 601.950 ;
        RECT 467.700 594.600 468.900 596.700 ;
        RECT 497.100 595.800 501.300 596.700 ;
        RECT 446.100 588.000 447.900 591.600 ;
        RECT 449.100 588.600 450.900 591.600 ;
        RECT 467.100 588.600 468.900 594.600 ;
        RECT 470.100 593.700 477.900 595.050 ;
        RECT 470.100 588.600 471.900 593.700 ;
        RECT 473.100 588.000 474.900 592.800 ;
        RECT 476.100 588.600 477.900 593.700 ;
        RECT 494.400 588.000 496.200 594.600 ;
        RECT 499.500 588.600 501.300 595.800 ;
        RECT 521.400 591.600 522.300 601.950 ;
        RECT 542.100 600.150 543.900 601.950 ;
        RECT 545.700 596.700 546.900 601.950 ;
        RECT 547.950 600.150 549.750 601.950 ;
        RECT 566.250 600.150 568.050 601.950 ;
        RECT 542.700 595.800 546.900 596.700 ;
        RECT 569.100 596.700 570.300 601.950 ;
        RECT 572.100 600.150 573.900 601.950 ;
        RECT 590.100 600.150 591.900 601.950 ;
        RECT 569.100 595.800 573.300 596.700 ;
        RECT 518.100 588.000 519.900 591.600 ;
        RECT 521.100 588.600 522.900 591.600 ;
        RECT 524.100 588.000 525.900 591.600 ;
        RECT 542.700 588.600 544.500 595.800 ;
        RECT 547.800 588.000 549.600 594.600 ;
        RECT 566.400 588.000 568.200 594.600 ;
        RECT 571.500 588.600 573.300 595.800 ;
        RECT 596.700 594.600 597.900 601.950 ;
        RECT 601.950 600.150 603.750 601.950 ;
        RECT 620.100 600.150 621.900 601.950 ;
        RECT 623.100 594.600 624.300 601.950 ;
        RECT 592.500 588.000 594.300 594.600 ;
        RECT 597.000 588.600 598.800 594.600 ;
        RECT 601.500 588.000 603.300 594.600 ;
        RECT 620.100 588.000 621.900 594.600 ;
        RECT 623.100 588.600 624.900 594.600 ;
        RECT 644.400 591.600 645.300 601.950 ;
        RECT 665.250 600.150 667.050 601.950 ;
        RECT 646.950 597.450 649.050 598.050 ;
        RECT 652.950 597.450 655.050 597.900 ;
        RECT 646.950 596.550 655.050 597.450 ;
        RECT 646.950 595.950 649.050 596.550 ;
        RECT 652.950 595.800 655.050 596.550 ;
        RECT 671.100 594.600 672.300 601.950 ;
        RECT 677.100 600.150 678.900 601.950 ;
        RECT 679.950 600.450 682.050 601.050 ;
        RECT 679.950 599.550 693.450 600.450 ;
        RECT 698.250 600.150 700.050 601.950 ;
        RECT 679.950 598.950 682.050 599.550 ;
        RECT 676.950 597.450 679.050 598.050 ;
        RECT 688.950 597.450 691.050 598.050 ;
        RECT 676.950 596.550 691.050 597.450 ;
        RECT 676.950 595.950 679.050 596.550 ;
        RECT 688.950 595.950 691.050 596.550 ;
        RECT 692.550 595.050 693.450 599.550 ;
        RECT 702.000 597.300 703.050 601.950 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 703.950 600.150 705.750 601.950 ;
        RECT 719.550 601.050 720.450 608.550 ;
        RECT 727.950 607.950 730.050 608.550 ;
        RECT 731.100 609.600 735.900 610.500 ;
        RECT 728.250 604.050 730.050 605.850 ;
        RECT 731.100 604.050 732.000 609.600 ;
        RECT 734.100 604.050 735.900 605.850 ;
        RECT 755.400 604.050 756.300 611.400 ;
        RECT 760.950 604.050 762.750 605.850 ;
        RECT 783.000 604.050 784.200 611.400 ;
        RECT 791.700 609.900 792.900 611.400 ;
        RECT 785.100 608.700 792.900 609.900 ;
        RECT 785.100 608.100 786.900 608.700 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 763.950 601.950 766.050 604.050 ;
        RECT 782.100 601.950 784.200 604.050 ;
        RECT 711.000 600.450 715.050 601.050 ;
        RECT 698.700 596.100 703.050 597.300 ;
        RECT 710.550 598.950 715.050 600.450 ;
        RECT 719.550 599.550 724.050 601.050 ;
        RECT 725.250 600.150 727.050 601.950 ;
        RECT 720.000 598.950 724.050 599.550 ;
        RECT 641.100 588.000 642.900 591.600 ;
        RECT 644.100 588.600 645.900 591.600 ;
        RECT 647.100 588.000 648.900 591.600 ;
        RECT 665.700 588.000 667.500 594.600 ;
        RECT 670.200 588.600 672.000 594.600 ;
        RECT 674.700 588.000 676.500 594.600 ;
        RECT 691.950 592.950 694.050 595.050 ;
        RECT 698.700 594.600 699.600 596.100 ;
        RECT 695.100 589.500 696.900 594.600 ;
        RECT 698.100 590.400 699.900 594.600 ;
        RECT 701.100 594.000 708.900 594.900 ;
        RECT 701.100 589.500 702.900 594.000 ;
        RECT 695.100 588.600 702.900 589.500 ;
        RECT 704.100 588.000 705.900 593.100 ;
        RECT 707.100 588.600 708.900 594.000 ;
        RECT 710.550 594.450 711.450 598.950 ;
        RECT 712.950 597.450 715.050 597.900 ;
        RECT 727.950 597.450 730.050 597.750 ;
        RECT 712.950 596.550 730.050 597.450 ;
        RECT 712.950 595.800 715.050 596.550 ;
        RECT 727.950 595.650 730.050 596.550 ;
        RECT 721.950 594.450 724.050 595.050 ;
        RECT 731.100 594.600 732.300 601.950 ;
        RECT 737.100 600.150 738.900 601.950 ;
        RECT 755.400 594.600 756.300 601.950 ;
        RECT 757.950 600.150 759.750 601.950 ;
        RECT 764.100 600.150 765.900 601.950 ;
        RECT 763.950 597.450 766.050 598.050 ;
        RECT 778.950 597.450 781.050 598.050 ;
        RECT 763.950 596.550 781.050 597.450 ;
        RECT 763.950 595.950 766.050 596.550 ;
        RECT 778.950 595.950 781.050 596.550 ;
        RECT 710.550 593.550 724.050 594.450 ;
        RECT 721.950 592.950 724.050 593.550 ;
        RECT 725.700 588.000 727.500 594.600 ;
        RECT 730.200 588.600 732.000 594.600 ;
        RECT 734.700 588.000 736.500 594.600 ;
        RECT 755.400 593.400 760.500 594.600 ;
        RECT 755.700 588.000 757.500 591.600 ;
        RECT 758.700 588.600 760.500 593.400 ;
        RECT 763.200 588.000 765.000 594.600 ;
        RECT 766.950 594.450 769.050 595.050 ;
        RECT 772.950 594.450 775.050 595.050 ;
        RECT 766.950 593.550 775.050 594.450 ;
        RECT 766.950 592.950 769.050 593.550 ;
        RECT 772.950 592.950 775.050 593.550 ;
        RECT 782.100 594.600 783.000 601.950 ;
        RECT 785.400 597.600 786.300 608.100 ;
        RECT 804.000 606.450 808.050 607.050 ;
        RECT 787.200 604.050 789.000 605.850 ;
        RECT 803.550 604.950 808.050 606.450 ;
        RECT 787.500 601.950 789.600 604.050 ;
        RECT 790.800 601.950 792.900 604.050 ;
        RECT 790.800 600.150 792.600 601.950 ;
        RECT 803.550 601.050 804.450 604.950 ;
        RECT 812.700 604.050 813.900 617.400 ;
        RECT 834.000 612.600 835.800 623.400 ;
        RECT 834.000 611.400 837.600 612.600 ;
        RECT 839.100 611.400 840.900 624.000 ;
        RECT 857.100 617.400 858.900 624.000 ;
        RECT 860.100 617.400 861.900 623.400 ;
        RECT 863.100 617.400 864.900 624.000 ;
        RECT 881.100 617.400 882.900 623.400 ;
        RECT 884.100 618.000 885.900 624.000 ;
        RECT 833.100 604.050 834.900 605.850 ;
        RECT 836.700 604.050 837.600 611.400 ;
        RECT 841.950 606.450 846.000 607.050 ;
        RECT 838.950 604.050 840.750 605.850 ;
        RECT 841.950 604.950 846.450 606.450 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 803.550 599.550 808.050 601.050 ;
        RECT 809.100 600.150 810.900 601.950 ;
        RECT 804.000 598.950 808.050 599.550 ;
        RECT 784.200 596.700 786.300 597.600 ;
        RECT 812.700 596.700 813.900 601.950 ;
        RECT 814.950 600.150 816.750 601.950 ;
        RECT 823.950 600.450 826.050 601.050 ;
        RECT 829.950 600.450 832.050 601.050 ;
        RECT 823.950 599.550 832.050 600.450 ;
        RECT 823.950 598.950 826.050 599.550 ;
        RECT 829.950 598.950 832.050 599.550 ;
        RECT 784.200 595.800 789.600 596.700 ;
        RECT 782.100 588.600 783.900 594.600 ;
        RECT 785.100 588.000 786.900 594.000 ;
        RECT 788.700 591.600 789.600 595.800 ;
        RECT 809.700 595.800 813.900 596.700 ;
        RECT 814.950 597.450 817.050 598.050 ;
        RECT 832.950 597.450 835.050 598.050 ;
        RECT 814.950 596.550 835.050 597.450 ;
        RECT 814.950 595.950 817.050 596.550 ;
        RECT 832.950 595.950 835.050 596.550 ;
        RECT 788.100 588.600 789.900 591.600 ;
        RECT 791.100 588.600 792.900 591.600 ;
        RECT 809.700 588.600 811.500 595.800 ;
        RECT 791.700 588.000 792.900 588.600 ;
        RECT 814.800 588.000 816.600 594.600 ;
        RECT 817.950 591.450 820.050 592.050 ;
        RECT 829.950 591.450 832.050 592.050 ;
        RECT 836.700 591.600 837.600 601.950 ;
        RECT 845.550 601.050 846.450 604.950 ;
        RECT 860.700 604.050 861.900 617.400 ;
        RECT 882.000 617.100 882.900 617.400 ;
        RECT 887.100 617.400 888.900 623.400 ;
        RECT 890.100 617.400 891.900 624.000 ;
        RECT 887.100 617.100 888.600 617.400 ;
        RECT 882.000 616.200 888.600 617.100 ;
        RECT 871.950 606.450 874.050 607.050 ;
        RECT 877.950 606.450 880.050 607.050 ;
        RECT 871.950 605.550 880.050 606.450 ;
        RECT 871.950 604.950 874.050 605.550 ;
        RECT 877.950 604.950 880.050 605.550 ;
        RECT 882.000 604.050 882.900 616.200 ;
        RECT 908.400 611.400 910.200 624.000 ;
        RECT 913.500 612.900 915.300 623.400 ;
        RECT 916.500 617.400 918.300 624.000 ;
        RECT 935.100 617.400 936.900 624.000 ;
        RECT 938.100 617.400 939.900 623.400 ;
        RECT 941.100 617.400 942.900 624.000 ;
        RECT 916.200 614.100 918.000 615.900 ;
        RECT 913.500 611.400 915.900 612.900 ;
        RECT 887.100 604.050 888.900 605.850 ;
        RECT 908.100 604.050 909.900 605.850 ;
        RECT 914.700 604.050 915.900 611.400 ;
        RECT 916.950 612.450 919.050 613.050 ;
        RECT 934.950 612.450 937.050 613.050 ;
        RECT 916.950 611.550 937.050 612.450 ;
        RECT 916.950 610.950 919.050 611.550 ;
        RECT 934.950 610.950 937.050 611.550 ;
        RECT 938.100 604.050 939.300 617.400 ;
        RECT 959.100 611.400 960.900 623.400 ;
        RECT 962.100 611.400 963.900 624.000 ;
        RECT 980.100 611.400 981.900 624.000 ;
        RECT 985.200 612.600 987.000 623.400 ;
        RECT 983.400 611.400 987.000 612.600 ;
        RECT 1004.100 611.400 1005.900 624.000 ;
        RECT 1009.200 612.600 1011.000 623.400 ;
        RECT 1028.100 617.400 1029.900 623.400 ;
        RECT 1031.100 617.400 1032.900 624.000 ;
        RECT 1007.400 611.400 1011.000 612.600 ;
        RECT 1012.950 612.450 1015.050 613.050 ;
        RECT 1024.950 612.450 1027.050 613.050 ;
        RECT 1012.950 611.550 1027.050 612.450 ;
        RECT 943.950 606.450 946.050 607.050 ;
        RECT 943.950 605.550 954.450 606.450 ;
        RECT 943.950 604.950 946.050 605.550 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 916.950 601.950 919.050 604.050 ;
        RECT 934.950 601.950 937.050 604.050 ;
        RECT 937.950 601.950 940.050 604.050 ;
        RECT 940.950 601.950 943.050 604.050 ;
        RECT 841.950 599.550 846.450 601.050 ;
        RECT 857.100 600.150 858.900 601.950 ;
        RECT 841.950 598.950 846.000 599.550 ;
        RECT 838.950 597.450 841.050 598.050 ;
        RECT 850.950 597.450 853.050 598.050 ;
        RECT 838.950 596.550 853.050 597.450 ;
        RECT 860.700 596.700 861.900 601.950 ;
        RECT 862.950 600.150 864.750 601.950 ;
        RECT 882.000 598.200 882.900 601.950 ;
        RECT 884.100 600.150 885.900 601.950 ;
        RECT 890.100 600.150 891.900 601.950 ;
        RECT 911.100 600.150 912.900 601.950 ;
        RECT 882.000 597.000 885.300 598.200 ;
        RECT 914.700 597.600 915.900 601.950 ;
        RECT 917.100 600.150 918.900 601.950 ;
        RECT 935.250 600.150 937.050 601.950 ;
        RECT 838.950 595.950 841.050 596.550 ;
        RECT 850.950 595.950 853.050 596.550 ;
        RECT 857.700 595.800 861.900 596.700 ;
        RECT 817.950 590.550 832.050 591.450 ;
        RECT 817.950 589.950 820.050 590.550 ;
        RECT 829.950 589.950 832.050 590.550 ;
        RECT 833.100 588.000 834.900 591.600 ;
        RECT 836.100 588.600 837.900 591.600 ;
        RECT 839.100 588.000 840.900 591.600 ;
        RECT 844.950 591.450 847.050 591.900 ;
        RECT 853.950 591.450 856.050 592.050 ;
        RECT 844.950 590.550 856.050 591.450 ;
        RECT 844.950 589.800 847.050 590.550 ;
        RECT 853.950 589.950 856.050 590.550 ;
        RECT 857.700 588.600 859.500 595.800 ;
        RECT 862.800 588.000 864.600 594.600 ;
        RECT 883.500 588.600 885.300 597.000 ;
        RECT 890.100 588.000 891.900 597.600 ;
        RECT 914.700 596.700 918.300 597.600 ;
        RECT 908.100 593.700 915.900 595.050 ;
        RECT 908.100 588.600 909.900 593.700 ;
        RECT 911.100 588.000 912.900 592.800 ;
        RECT 914.100 588.600 915.900 593.700 ;
        RECT 917.100 594.600 918.300 596.700 ;
        RECT 938.100 596.700 939.300 601.950 ;
        RECT 941.100 600.150 942.900 601.950 ;
        RECT 953.550 601.050 954.450 605.550 ;
        RECT 959.700 604.050 960.900 611.400 ;
        RECT 961.950 609.450 964.050 610.050 ;
        RECT 976.950 609.450 979.050 610.050 ;
        RECT 961.950 608.550 979.050 609.450 ;
        RECT 961.950 607.950 964.050 608.550 ;
        RECT 976.950 607.950 979.050 608.550 ;
        RECT 980.250 604.050 982.050 605.850 ;
        RECT 983.400 604.050 984.300 611.400 ;
        RECT 985.950 609.450 988.050 610.050 ;
        RECT 994.950 609.450 997.050 610.050 ;
        RECT 985.950 608.550 997.050 609.450 ;
        RECT 985.950 607.950 988.050 608.550 ;
        RECT 994.950 607.950 997.050 608.550 ;
        RECT 988.950 606.450 991.050 607.050 ;
        RECT 997.950 606.450 1000.050 607.050 ;
        RECT 986.100 604.050 987.900 605.850 ;
        RECT 988.950 605.550 1000.050 606.450 ;
        RECT 988.950 604.950 991.050 605.550 ;
        RECT 997.950 604.950 1000.050 605.550 ;
        RECT 1004.250 604.050 1006.050 605.850 ;
        RECT 1007.400 604.050 1008.300 611.400 ;
        RECT 1012.950 610.950 1015.050 611.550 ;
        RECT 1024.950 610.950 1027.050 611.550 ;
        RECT 1010.100 604.050 1011.900 605.850 ;
        RECT 1028.700 604.050 1029.900 617.400 ;
        RECT 1031.100 604.050 1032.900 605.850 ;
        RECT 958.950 601.950 961.050 604.050 ;
        RECT 961.950 601.950 964.050 604.050 ;
        RECT 979.950 601.950 982.050 604.050 ;
        RECT 982.950 601.950 985.050 604.050 ;
        RECT 985.950 601.950 988.050 604.050 ;
        RECT 1003.950 601.950 1006.050 604.050 ;
        RECT 1006.950 601.950 1009.050 604.050 ;
        RECT 1009.950 601.950 1012.050 604.050 ;
        RECT 1027.950 601.950 1030.050 604.050 ;
        RECT 1030.950 601.950 1033.050 604.050 ;
        RECT 953.550 599.550 958.050 601.050 ;
        RECT 954.000 598.950 958.050 599.550 ;
        RECT 938.100 595.800 942.300 596.700 ;
        RECT 917.100 588.600 918.900 594.600 ;
        RECT 935.400 588.000 937.200 594.600 ;
        RECT 940.500 588.600 942.300 595.800 ;
        RECT 959.700 594.600 960.900 601.950 ;
        RECT 962.100 600.150 963.900 601.950 ;
        RECT 959.100 588.600 960.900 594.600 ;
        RECT 962.100 588.000 963.900 594.600 ;
        RECT 983.400 591.600 984.300 601.950 ;
        RECT 1007.400 591.600 1008.300 601.950 ;
        RECT 1015.950 597.450 1018.050 598.050 ;
        RECT 1010.550 597.000 1018.050 597.450 ;
        RECT 1009.950 596.550 1018.050 597.000 ;
        RECT 1009.950 592.950 1012.050 596.550 ;
        RECT 1015.950 595.950 1018.050 596.550 ;
        RECT 1028.700 591.600 1029.900 601.950 ;
        RECT 1030.950 597.450 1033.050 598.050 ;
        RECT 1039.950 597.450 1042.050 598.050 ;
        RECT 1030.950 596.550 1042.050 597.450 ;
        RECT 1030.950 595.950 1033.050 596.550 ;
        RECT 1039.950 595.950 1042.050 596.550 ;
        RECT 980.100 588.000 981.900 591.600 ;
        RECT 983.100 588.600 984.900 591.600 ;
        RECT 986.100 588.000 987.900 591.600 ;
        RECT 1004.100 588.000 1005.900 591.600 ;
        RECT 1007.100 588.600 1008.900 591.600 ;
        RECT 1010.100 588.000 1011.900 591.600 ;
        RECT 1028.100 588.600 1029.900 591.600 ;
        RECT 1031.100 588.000 1032.900 591.600 ;
        RECT 17.100 575.400 18.900 585.000 ;
        RECT 23.700 576.000 25.500 584.400 ;
        RECT 45.000 578.400 46.800 585.000 ;
        RECT 49.500 579.600 51.300 584.400 ;
        RECT 52.500 581.400 54.300 585.000 ;
        RECT 71.100 581.400 72.900 585.000 ;
        RECT 74.100 581.400 75.900 584.400 ;
        RECT 92.700 581.400 94.500 585.000 ;
        RECT 49.500 578.400 54.600 579.600 ;
        RECT 23.700 574.800 27.000 576.000 ;
        RECT 17.100 571.050 18.900 572.850 ;
        RECT 23.100 571.050 24.900 572.850 ;
        RECT 26.100 571.050 27.000 574.800 ;
        RECT 44.100 571.050 45.900 572.850 ;
        RECT 50.250 571.050 52.050 572.850 ;
        RECT 53.700 571.050 54.600 578.400 ;
        RECT 74.100 571.050 75.300 581.400 ;
        RECT 95.700 579.600 97.500 584.400 ;
        RECT 92.400 578.400 97.500 579.600 ;
        RECT 100.200 578.400 102.000 585.000 ;
        RECT 119.100 581.400 120.900 585.000 ;
        RECT 122.100 581.400 123.900 584.400 ;
        RECT 125.100 581.400 126.900 585.000 ;
        RECT 143.100 581.400 144.900 585.000 ;
        RECT 146.100 581.400 147.900 584.400 ;
        RECT 149.100 581.400 150.900 585.000 ;
        RECT 92.400 571.050 93.300 578.400 ;
        RECT 94.950 571.050 96.750 572.850 ;
        RECT 101.100 571.050 102.900 572.850 ;
        RECT 122.700 571.050 123.600 581.400 ;
        RECT 133.950 576.450 136.050 577.050 ;
        RECT 142.950 576.450 145.050 577.050 ;
        RECT 133.950 575.550 145.050 576.450 ;
        RECT 133.950 574.950 136.050 575.550 ;
        RECT 142.950 574.950 145.050 575.550 ;
        RECT 146.700 571.050 147.600 581.400 ;
        RECT 152.700 578.400 154.500 584.400 ;
        RECT 158.100 578.400 159.900 585.000 ;
        RECT 163.500 578.400 165.300 584.400 ;
        RECT 167.700 581.400 169.500 584.400 ;
        RECT 170.700 581.400 172.500 584.400 ;
        RECT 173.700 581.400 175.500 584.400 ;
        RECT 176.700 581.400 178.500 585.000 ;
        RECT 167.700 579.300 169.800 581.400 ;
        RECT 170.700 579.300 172.800 581.400 ;
        RECT 173.700 579.300 175.800 581.400 ;
        RECT 181.200 580.500 183.000 584.400 ;
        RECT 184.200 581.400 186.000 585.000 ;
        RECT 187.200 581.400 189.000 584.400 ;
        RECT 190.200 581.400 192.000 584.400 ;
        RECT 193.200 581.400 195.000 584.400 ;
        RECT 196.200 581.400 198.000 584.400 ;
        RECT 177.600 579.600 179.400 580.500 ;
        RECT 176.700 578.400 179.400 579.600 ;
        RECT 181.200 578.400 183.900 580.500 ;
        RECT 187.200 579.300 189.300 581.400 ;
        RECT 190.200 579.300 192.300 581.400 ;
        RECT 193.200 579.300 195.300 581.400 ;
        RECT 196.200 579.300 198.300 581.400 ;
        RECT 200.400 579.600 202.200 584.400 ;
        RECT 200.400 578.400 204.600 579.600 ;
        RECT 205.500 578.400 207.300 585.000 ;
        RECT 210.900 578.400 212.700 584.400 ;
        RECT 152.700 574.800 153.900 578.400 ;
        RECT 163.800 577.500 165.300 578.400 ;
        RECT 172.800 577.800 174.600 578.400 ;
        RECT 176.700 577.800 177.600 578.400 ;
        RECT 156.900 576.300 165.300 577.500 ;
        RECT 170.400 576.600 177.600 577.800 ;
        RECT 192.300 576.600 198.900 578.400 ;
        RECT 156.900 575.700 158.700 576.300 ;
        RECT 167.400 574.800 169.500 575.700 ;
        RECT 152.700 573.600 169.500 574.800 ;
        RECT 170.400 573.600 171.300 576.600 ;
        RECT 175.800 573.900 177.600 574.800 ;
        RECT 185.100 574.500 186.900 576.300 ;
        RECT 203.100 575.100 204.600 578.400 ;
        RECT 178.800 573.900 180.900 574.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 43.950 568.950 46.050 571.050 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 91.950 568.950 94.050 571.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 121.950 568.950 124.050 571.050 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 142.950 568.950 145.050 571.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 20.100 567.150 21.900 568.950 ;
        RECT 26.100 556.800 27.000 568.950 ;
        RECT 47.250 567.150 49.050 568.950 ;
        RECT 53.700 561.600 54.600 568.950 ;
        RECT 71.100 567.150 72.900 568.950 ;
        RECT 20.400 555.900 27.000 556.800 ;
        RECT 20.400 555.600 21.900 555.900 ;
        RECT 17.100 549.000 18.900 555.600 ;
        RECT 20.100 549.600 21.900 555.600 ;
        RECT 26.100 555.600 27.000 555.900 ;
        RECT 44.100 560.700 51.900 561.600 ;
        RECT 23.100 549.000 24.900 555.000 ;
        RECT 26.100 549.600 27.900 555.600 ;
        RECT 44.100 549.600 45.900 560.700 ;
        RECT 47.100 549.000 48.900 559.800 ;
        RECT 50.100 549.600 51.900 560.700 ;
        RECT 53.100 549.600 54.900 561.600 ;
        RECT 74.100 555.600 75.300 568.950 ;
        RECT 92.400 561.600 93.300 568.950 ;
        RECT 97.950 567.150 99.750 568.950 ;
        RECT 119.100 567.150 120.900 568.950 ;
        RECT 100.950 564.450 103.050 565.050 ;
        RECT 118.950 564.450 121.050 565.050 ;
        RECT 100.950 563.550 121.050 564.450 ;
        RECT 100.950 562.950 103.050 563.550 ;
        RECT 118.950 562.950 121.050 563.550 ;
        RECT 122.700 561.600 123.600 568.950 ;
        RECT 124.950 567.150 126.750 568.950 ;
        RECT 143.100 567.150 144.900 568.950 ;
        RECT 146.700 561.600 147.600 568.950 ;
        RECT 148.950 567.150 150.750 568.950 ;
        RECT 71.100 549.000 72.900 555.600 ;
        RECT 74.100 549.600 75.900 555.600 ;
        RECT 92.100 549.600 93.900 561.600 ;
        RECT 95.100 560.700 102.900 561.600 ;
        RECT 95.100 549.600 96.900 560.700 ;
        RECT 98.100 549.000 99.900 559.800 ;
        RECT 101.100 549.600 102.900 560.700 ;
        RECT 120.000 560.400 123.600 561.600 ;
        RECT 120.000 549.600 121.800 560.400 ;
        RECT 125.100 549.000 126.900 561.600 ;
        RECT 144.000 560.400 147.600 561.600 ;
        RECT 144.000 549.600 145.800 560.400 ;
        RECT 149.100 549.000 150.900 561.600 ;
        RECT 152.700 557.400 153.900 573.600 ;
        RECT 170.400 571.800 172.200 573.600 ;
        RECT 175.800 573.000 180.900 573.900 ;
        RECT 178.800 571.950 180.900 573.000 ;
        RECT 185.100 573.900 187.200 574.500 ;
        RECT 185.100 572.400 202.200 573.900 ;
        RECT 203.100 573.300 210.900 575.100 ;
        RECT 200.700 570.900 207.300 572.400 ;
        RECT 155.100 569.700 199.500 570.900 ;
        RECT 155.100 568.050 156.900 569.700 ;
        RECT 154.800 565.950 156.900 568.050 ;
        RECT 160.800 567.750 162.900 568.050 ;
        RECT 173.400 567.900 175.200 568.500 ;
        RECT 182.400 567.900 195.900 568.800 ;
        RECT 160.800 565.950 164.700 567.750 ;
        RECT 173.400 566.700 184.500 567.900 ;
        RECT 162.900 565.200 164.700 565.950 ;
        RECT 182.400 565.800 184.500 566.700 ;
        RECT 186.000 565.200 189.900 567.000 ;
        RECT 195.000 566.700 195.900 567.900 ;
        RECT 162.900 564.300 176.400 565.200 ;
        RECT 187.800 564.900 189.900 565.200 ;
        RECT 194.100 564.900 195.900 566.700 ;
        RECT 198.600 568.200 199.500 569.700 ;
        RECT 198.600 566.400 203.700 568.200 ;
        RECT 205.800 568.050 207.300 570.900 ;
        RECT 205.800 565.950 207.900 568.050 ;
        RECT 175.200 563.700 176.400 564.300 ;
        RECT 209.100 563.700 210.900 564.300 ;
        RECT 170.400 562.500 172.500 562.800 ;
        RECT 175.200 562.500 210.900 563.700 ;
        RECT 160.500 561.300 172.500 562.500 ;
        RECT 211.800 561.600 212.700 578.400 ;
        RECT 160.500 560.700 162.300 561.300 ;
        RECT 170.400 560.700 172.500 561.300 ;
        RECT 175.200 560.400 192.900 561.600 ;
        RECT 157.200 559.800 159.000 560.100 ;
        RECT 175.200 559.800 176.400 560.400 ;
        RECT 157.200 558.600 176.400 559.800 ;
        RECT 190.800 559.500 192.900 560.400 ;
        RECT 196.200 560.700 212.700 561.600 ;
        RECT 196.200 559.500 198.300 560.700 ;
        RECT 157.200 558.300 159.000 558.600 ;
        RECT 152.700 556.500 156.300 557.400 ;
        RECT 155.400 555.600 156.300 556.500 ;
        RECT 152.700 549.000 154.500 555.600 ;
        RECT 155.400 554.700 157.500 555.600 ;
        RECT 155.700 549.600 157.500 554.700 ;
        RECT 158.700 549.000 160.500 555.600 ;
        RECT 161.700 549.600 163.500 558.600 ;
        RECT 173.700 555.600 175.800 557.700 ;
        RECT 181.200 557.100 184.500 559.200 ;
        RECT 164.700 549.000 166.500 555.600 ;
        RECT 168.300 552.600 170.400 554.700 ;
        RECT 171.300 552.600 173.400 554.700 ;
        RECT 168.300 549.600 170.100 552.600 ;
        RECT 171.300 549.600 173.100 552.600 ;
        RECT 174.300 549.600 176.100 555.600 ;
        RECT 177.300 549.000 179.100 555.600 ;
        RECT 181.200 549.600 183.000 557.100 ;
        RECT 187.200 555.600 189.900 559.500 ;
        RECT 202.200 558.600 207.900 559.800 ;
        RECT 199.500 557.700 201.300 558.300 ;
        RECT 193.200 556.500 201.300 557.700 ;
        RECT 193.200 555.600 195.300 556.500 ;
        RECT 202.200 555.600 203.400 558.600 ;
        RECT 206.100 558.000 207.900 558.600 ;
        RECT 211.800 557.400 212.700 560.700 ;
        RECT 208.800 556.500 212.700 557.400 ;
        RECT 214.500 581.400 216.300 584.400 ;
        RECT 217.500 581.400 219.300 585.000 ;
        RECT 214.500 568.050 216.000 581.400 ;
        RECT 238.500 576.000 240.300 584.400 ;
        RECT 237.000 574.800 240.300 576.000 ;
        RECT 245.100 575.400 246.900 585.000 ;
        RECT 264.000 578.400 265.800 585.000 ;
        RECT 268.500 579.600 270.300 584.400 ;
        RECT 271.500 581.400 273.300 585.000 ;
        RECT 290.100 581.400 291.900 584.400 ;
        RECT 293.100 581.400 294.900 585.000 ;
        RECT 268.500 578.400 273.600 579.600 ;
        RECT 237.000 571.050 237.900 574.800 ;
        RECT 239.100 571.050 240.900 572.850 ;
        RECT 245.100 571.050 246.900 572.850 ;
        RECT 263.100 571.050 264.900 572.850 ;
        RECT 269.250 571.050 271.050 572.850 ;
        RECT 272.700 571.050 273.600 578.400 ;
        RECT 290.700 571.050 291.900 581.400 ;
        RECT 311.100 575.400 312.900 585.000 ;
        RECT 317.700 576.000 319.500 584.400 ;
        RECT 338.400 578.400 340.200 585.000 ;
        RECT 343.500 577.200 345.300 584.400 ;
        RECT 362.100 583.500 369.900 584.400 ;
        RECT 362.100 578.400 363.900 583.500 ;
        RECT 365.100 578.400 366.900 582.600 ;
        RECT 368.100 579.000 369.900 583.500 ;
        RECT 371.100 579.900 372.900 585.000 ;
        RECT 374.100 579.000 375.900 584.400 ;
        RECT 400.200 581.400 402.900 584.400 ;
        RECT 404.100 581.400 405.900 585.000 ;
        RECT 407.100 581.400 408.900 584.400 ;
        RECT 410.100 581.400 412.200 585.000 ;
        RECT 400.200 580.500 401.100 581.400 ;
        RECT 407.400 580.500 408.300 581.400 ;
        RECT 341.100 576.300 345.300 577.200 ;
        RECT 365.700 576.900 366.600 578.400 ;
        RECT 368.100 578.100 375.900 579.000 ;
        RECT 395.700 579.600 408.300 580.500 ;
        RECT 317.700 574.800 321.000 576.000 ;
        RECT 311.100 571.050 312.900 572.850 ;
        RECT 317.100 571.050 318.900 572.850 ;
        RECT 320.100 571.050 321.000 574.800 ;
        RECT 322.950 573.450 325.050 574.050 ;
        RECT 331.950 573.450 334.050 574.050 ;
        RECT 322.950 572.550 334.050 573.450 ;
        RECT 322.950 571.950 325.050 572.550 ;
        RECT 331.950 571.950 334.050 572.550 ;
        RECT 338.250 571.050 340.050 572.850 ;
        RECT 341.100 571.050 342.300 576.300 ;
        RECT 365.700 575.700 370.050 576.900 ;
        RECT 344.100 571.050 345.900 572.850 ;
        RECT 365.250 571.050 367.050 572.850 ;
        RECT 369.000 571.050 370.050 575.700 ;
        RECT 385.950 576.450 388.050 577.050 ;
        RECT 391.950 576.450 394.050 577.050 ;
        RECT 385.950 575.550 394.050 576.450 ;
        RECT 385.950 574.950 388.050 575.550 ;
        RECT 391.950 574.950 394.050 575.550 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 319.950 568.950 322.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 340.950 568.950 343.050 571.050 ;
        RECT 343.950 568.950 346.050 571.050 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 370.950 571.050 372.750 572.850 ;
        RECT 395.700 571.050 396.900 579.600 ;
        RECT 428.100 578.400 429.900 584.400 ;
        RECT 428.700 576.300 429.900 578.400 ;
        RECT 431.100 579.300 432.900 584.400 ;
        RECT 434.100 580.200 435.900 585.000 ;
        RECT 437.100 579.300 438.900 584.400 ;
        RECT 455.700 581.400 457.500 585.000 ;
        RECT 458.700 579.600 460.500 584.400 ;
        RECT 431.100 577.950 438.900 579.300 ;
        RECT 455.400 578.400 460.500 579.600 ;
        RECT 463.200 578.400 465.000 585.000 ;
        RECT 483.600 580.200 485.400 584.400 ;
        RECT 482.700 578.400 485.400 580.200 ;
        RECT 486.600 578.400 488.400 585.000 ;
        RECT 428.700 575.400 432.300 576.300 ;
        RECT 404.250 571.050 406.050 572.850 ;
        RECT 428.100 571.050 429.900 572.850 ;
        RECT 431.100 571.050 432.300 575.400 ;
        RECT 434.100 571.050 435.900 572.850 ;
        RECT 455.400 571.050 456.300 578.400 ;
        RECT 457.950 576.450 460.050 577.050 ;
        RECT 472.950 576.450 475.050 577.050 ;
        RECT 457.950 575.550 475.050 576.450 ;
        RECT 457.950 574.950 460.050 575.550 ;
        RECT 472.950 574.950 475.050 575.550 ;
        RECT 457.950 571.050 459.750 572.850 ;
        RECT 464.100 571.050 465.900 572.850 ;
        RECT 482.700 571.050 483.600 578.400 ;
        RECT 484.500 576.600 486.300 577.500 ;
        RECT 491.100 576.600 492.900 584.400 ;
        RECT 509.100 581.400 510.900 585.000 ;
        RECT 512.100 581.400 513.900 584.400 ;
        RECT 515.100 581.400 516.900 585.000 ;
        RECT 533.100 581.400 534.900 585.000 ;
        RECT 536.100 581.400 537.900 584.400 ;
        RECT 539.100 581.400 540.900 585.000 ;
        RECT 484.500 575.700 492.900 576.600 ;
        RECT 496.950 576.450 499.050 577.050 ;
        RECT 508.950 576.450 511.050 577.200 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 395.400 568.950 397.500 571.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 403.950 568.950 406.050 571.050 ;
        RECT 410.100 568.950 412.200 571.050 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 454.950 568.950 457.050 571.050 ;
        RECT 457.950 568.950 460.050 571.050 ;
        RECT 460.950 568.950 463.050 571.050 ;
        RECT 463.950 568.950 466.050 571.050 ;
        RECT 482.100 568.950 484.200 571.050 ;
        RECT 485.400 568.950 487.500 571.050 ;
        RECT 214.500 565.950 216.900 568.050 ;
        RECT 208.800 555.600 210.000 556.500 ;
        RECT 214.500 555.600 216.000 565.950 ;
        RECT 237.000 556.800 237.900 568.950 ;
        RECT 242.100 567.150 243.900 568.950 ;
        RECT 266.250 567.150 268.050 568.950 ;
        RECT 238.950 564.450 241.050 565.050 ;
        RECT 259.950 564.450 262.050 565.050 ;
        RECT 238.950 563.550 262.050 564.450 ;
        RECT 238.950 562.950 241.050 563.550 ;
        RECT 259.950 562.950 262.050 563.550 ;
        RECT 272.700 561.600 273.600 568.950 ;
        RECT 263.100 560.700 270.900 561.600 ;
        RECT 237.000 555.900 243.600 556.800 ;
        RECT 237.000 555.600 237.900 555.900 ;
        RECT 184.200 549.000 186.000 555.600 ;
        RECT 187.200 549.600 189.000 555.600 ;
        RECT 190.200 552.600 192.300 554.700 ;
        RECT 193.200 552.600 195.300 554.700 ;
        RECT 196.200 552.600 198.300 554.700 ;
        RECT 190.200 549.600 192.000 552.600 ;
        RECT 193.200 549.600 195.000 552.600 ;
        RECT 196.200 549.600 198.000 552.600 ;
        RECT 199.200 549.000 201.000 555.600 ;
        RECT 202.200 549.600 204.000 555.600 ;
        RECT 205.200 549.000 207.000 555.600 ;
        RECT 208.200 549.600 210.000 555.600 ;
        RECT 211.200 549.000 213.000 555.600 ;
        RECT 214.500 549.600 216.300 555.600 ;
        RECT 217.500 549.000 219.300 555.600 ;
        RECT 236.100 549.600 237.900 555.600 ;
        RECT 242.100 555.600 243.600 555.900 ;
        RECT 239.100 549.000 240.900 555.000 ;
        RECT 242.100 549.600 243.900 555.600 ;
        RECT 245.100 549.000 246.900 555.600 ;
        RECT 263.100 549.600 264.900 560.700 ;
        RECT 266.100 549.000 267.900 559.800 ;
        RECT 269.100 549.600 270.900 560.700 ;
        RECT 272.100 549.600 273.900 561.600 ;
        RECT 290.700 555.600 291.900 568.950 ;
        RECT 293.100 567.150 294.900 568.950 ;
        RECT 314.100 567.150 315.900 568.950 ;
        RECT 304.950 564.450 307.050 565.050 ;
        RECT 316.950 564.450 319.050 565.050 ;
        RECT 304.950 563.550 319.050 564.450 ;
        RECT 304.950 562.950 307.050 563.550 ;
        RECT 316.950 562.950 319.050 563.550 ;
        RECT 320.100 556.800 321.000 568.950 ;
        RECT 314.400 555.900 321.000 556.800 ;
        RECT 314.400 555.600 315.900 555.900 ;
        RECT 274.950 552.450 277.050 553.050 ;
        RECT 283.950 552.450 286.050 553.050 ;
        RECT 274.950 551.550 286.050 552.450 ;
        RECT 274.950 550.950 277.050 551.550 ;
        RECT 283.950 550.950 286.050 551.550 ;
        RECT 290.100 549.600 291.900 555.600 ;
        RECT 293.100 549.000 294.900 555.600 ;
        RECT 311.100 549.000 312.900 555.600 ;
        RECT 314.100 549.600 315.900 555.600 ;
        RECT 320.100 555.600 321.000 555.900 ;
        RECT 341.100 555.600 342.300 568.950 ;
        RECT 362.250 567.150 364.050 568.950 ;
        RECT 369.000 561.600 370.050 568.950 ;
        RECT 374.100 567.150 375.900 568.950 ;
        RECT 317.100 549.000 318.900 555.000 ;
        RECT 320.100 549.600 321.900 555.600 ;
        RECT 338.100 549.000 339.900 555.600 ;
        RECT 341.100 549.600 342.900 555.600 ;
        RECT 344.100 549.000 345.900 555.600 ;
        RECT 363.600 549.000 365.400 561.600 ;
        RECT 368.100 549.600 371.400 561.600 ;
        RECT 374.100 549.000 375.900 561.600 ;
        RECT 392.100 550.500 393.900 559.800 ;
        RECT 395.700 559.200 396.900 568.950 ;
        RECT 400.950 567.150 402.750 568.950 ;
        RECT 410.100 567.150 411.900 568.950 ;
        RECT 431.100 561.600 432.300 568.950 ;
        RECT 437.100 567.150 438.900 568.950 ;
        RECT 436.950 564.450 439.050 565.050 ;
        RECT 448.950 564.450 451.050 565.050 ;
        RECT 436.950 563.550 451.050 564.450 ;
        RECT 436.950 562.950 439.050 563.550 ;
        RECT 448.950 562.950 451.050 563.550 ;
        RECT 455.400 561.600 456.300 568.950 ;
        RECT 460.950 567.150 462.750 568.950 ;
        RECT 466.950 567.450 469.050 568.050 ;
        RECT 472.950 567.450 475.050 568.050 ;
        RECT 466.950 566.550 475.050 567.450 ;
        RECT 466.950 565.950 469.050 566.550 ;
        RECT 472.950 565.950 475.050 566.550 ;
        RECT 457.950 564.450 460.050 565.050 ;
        RECT 475.950 564.450 478.050 565.050 ;
        RECT 457.950 563.550 478.050 564.450 ;
        RECT 457.950 562.950 460.050 563.550 ;
        RECT 475.950 562.950 478.050 563.550 ;
        RECT 482.700 561.600 483.600 568.950 ;
        RECT 486.000 567.150 487.800 568.950 ;
        RECT 395.100 551.400 396.900 559.200 ;
        RECT 398.100 559.200 405.900 560.100 ;
        RECT 398.100 550.500 399.900 559.200 ;
        RECT 392.100 549.600 399.900 550.500 ;
        RECT 401.100 550.500 402.900 558.300 ;
        RECT 404.100 551.400 405.900 559.200 ;
        RECT 407.100 559.500 414.900 560.400 ;
        RECT 431.100 560.100 433.500 561.600 ;
        RECT 407.100 550.500 408.900 559.500 ;
        RECT 401.100 549.600 408.900 550.500 ;
        RECT 410.100 549.000 411.900 558.600 ;
        RECT 413.100 549.600 414.900 559.500 ;
        RECT 429.000 557.100 430.800 558.900 ;
        RECT 428.700 549.000 430.500 555.600 ;
        RECT 431.700 549.600 433.500 560.100 ;
        RECT 436.800 549.000 438.600 561.600 ;
        RECT 455.100 549.600 456.900 561.600 ;
        RECT 458.100 560.700 465.900 561.600 ;
        RECT 458.100 549.600 459.900 560.700 ;
        RECT 461.100 549.000 462.900 559.800 ;
        RECT 464.100 549.600 465.900 560.700 ;
        RECT 482.100 549.600 483.900 561.600 ;
        RECT 485.100 549.000 486.900 561.000 ;
        RECT 489.000 555.600 489.900 575.700 ;
        RECT 496.950 575.550 511.050 576.450 ;
        RECT 496.950 574.950 499.050 575.550 ;
        RECT 508.950 575.100 511.050 575.550 ;
        RECT 490.950 571.050 492.750 572.850 ;
        RECT 512.400 571.050 513.300 581.400 ;
        RECT 514.950 576.450 517.050 577.050 ;
        RECT 532.950 576.450 535.050 577.050 ;
        RECT 514.950 575.550 535.050 576.450 ;
        RECT 514.950 574.950 517.050 575.550 ;
        RECT 532.950 574.950 535.050 575.550 ;
        RECT 536.400 571.050 537.300 581.400 ;
        RECT 557.700 578.400 559.500 585.000 ;
        RECT 562.200 578.400 564.000 584.400 ;
        RECT 566.700 578.400 568.500 585.000 ;
        RECT 587.100 578.400 588.900 584.400 ;
        RECT 590.100 578.400 591.900 585.000 ;
        RECT 608.100 579.000 609.900 584.400 ;
        RECT 611.100 579.900 612.900 585.000 ;
        RECT 614.100 583.500 621.900 584.400 ;
        RECT 614.100 579.000 615.900 583.500 ;
        RECT 557.250 571.050 559.050 572.850 ;
        RECT 563.100 571.050 564.300 578.400 ;
        RECT 569.100 571.050 570.900 572.850 ;
        RECT 587.700 571.050 588.900 578.400 ;
        RECT 608.100 578.100 615.900 579.000 ;
        RECT 617.100 578.400 618.900 582.600 ;
        RECT 620.100 578.400 621.900 583.500 ;
        RECT 638.700 581.400 640.500 585.000 ;
        RECT 641.700 579.600 643.500 584.400 ;
        RECT 638.400 578.400 643.500 579.600 ;
        RECT 646.200 578.400 648.000 585.000 ;
        RECT 667.500 578.400 669.300 585.000 ;
        RECT 672.000 578.400 673.800 584.400 ;
        RECT 676.500 578.400 678.300 585.000 ;
        RECT 695.100 578.400 696.900 584.400 ;
        RECT 617.400 576.900 618.300 578.400 ;
        RECT 613.950 575.700 618.300 576.900 ;
        RECT 590.100 571.050 591.900 572.850 ;
        RECT 611.250 571.050 613.050 572.850 ;
        RECT 490.800 568.950 492.900 571.050 ;
        RECT 508.950 568.950 511.050 571.050 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 556.950 568.950 559.050 571.050 ;
        RECT 559.950 568.950 562.050 571.050 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 571.050 615.000 575.700 ;
        RECT 616.950 571.050 618.750 572.850 ;
        RECT 638.400 571.050 639.300 578.400 ;
        RECT 640.950 571.050 642.750 572.850 ;
        RECT 647.100 571.050 648.900 572.850 ;
        RECT 665.100 571.050 666.900 572.850 ;
        RECT 671.700 571.050 672.900 578.400 ;
        RECT 695.700 576.300 696.900 578.400 ;
        RECT 698.100 579.300 699.900 584.400 ;
        RECT 701.100 580.200 702.900 585.000 ;
        RECT 704.100 579.300 705.900 584.400 ;
        RECT 723.600 580.200 725.400 584.400 ;
        RECT 698.100 577.950 705.900 579.300 ;
        RECT 722.700 578.400 725.400 580.200 ;
        RECT 726.600 578.400 728.400 585.000 ;
        RECT 695.700 575.400 699.300 576.300 ;
        RECT 676.950 571.050 678.750 572.850 ;
        RECT 695.100 571.050 696.900 572.850 ;
        RECT 698.100 571.050 699.300 575.400 ;
        RECT 701.100 571.050 702.900 572.850 ;
        RECT 722.700 571.050 723.600 578.400 ;
        RECT 724.500 576.600 726.300 577.500 ;
        RECT 731.100 576.600 732.900 584.400 ;
        RECT 724.500 575.700 732.900 576.600 ;
        RECT 749.700 577.200 751.500 584.400 ;
        RECT 754.800 578.400 756.600 585.000 ;
        RECT 773.700 577.200 775.500 584.400 ;
        RECT 778.800 578.400 780.600 585.000 ;
        RECT 797.100 581.400 798.900 584.400 ;
        RECT 800.100 581.400 801.900 585.000 ;
        RECT 749.700 576.300 753.900 577.200 ;
        RECT 773.700 576.300 777.900 577.200 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 619.950 568.950 622.050 571.050 ;
        RECT 637.950 568.950 640.050 571.050 ;
        RECT 640.950 568.950 643.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 657.000 570.450 661.050 571.050 ;
        RECT 656.550 568.950 661.050 570.450 ;
        RECT 664.950 568.950 667.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 722.100 568.950 724.200 571.050 ;
        RECT 725.400 568.950 727.500 571.050 ;
        RECT 509.250 567.150 511.050 568.950 ;
        RECT 512.400 561.600 513.300 568.950 ;
        RECT 515.100 567.150 516.900 568.950 ;
        RECT 533.250 567.150 535.050 568.950 ;
        RECT 536.400 561.600 537.300 568.950 ;
        RECT 539.100 567.150 540.900 568.950 ;
        RECT 560.250 567.150 562.050 568.950 ;
        RECT 563.100 563.400 564.000 568.950 ;
        RECT 566.100 567.150 567.900 568.950 ;
        RECT 563.100 562.500 567.900 563.400 ;
        RECT 488.100 549.600 489.900 555.600 ;
        RECT 491.100 549.000 492.900 555.600 ;
        RECT 509.100 549.000 510.900 561.600 ;
        RECT 512.400 560.400 516.000 561.600 ;
        RECT 514.200 549.600 516.000 560.400 ;
        RECT 533.100 549.000 534.900 561.600 ;
        RECT 536.400 560.400 540.000 561.600 ;
        RECT 538.200 549.600 540.000 560.400 ;
        RECT 557.100 560.400 564.900 561.300 ;
        RECT 557.100 549.600 558.900 560.400 ;
        RECT 560.100 549.000 561.900 559.500 ;
        RECT 563.100 550.500 564.900 560.400 ;
        RECT 566.100 551.400 567.900 562.500 ;
        RECT 587.700 561.600 588.900 568.950 ;
        RECT 608.100 567.150 609.900 568.950 ;
        RECT 613.950 561.600 615.000 568.950 ;
        RECT 619.950 567.150 621.750 568.950 ;
        RECT 638.400 561.600 639.300 568.950 ;
        RECT 643.950 567.150 645.750 568.950 ;
        RECT 656.550 564.900 657.450 568.950 ;
        RECT 668.100 567.150 669.900 568.950 ;
        RECT 655.950 562.800 658.050 564.900 ;
        RECT 672.000 563.400 672.900 568.950 ;
        RECT 673.950 567.150 675.750 568.950 ;
        RECT 668.100 562.500 672.900 563.400 ;
        RECT 569.100 550.500 570.900 561.600 ;
        RECT 563.100 549.600 570.900 550.500 ;
        RECT 587.100 549.600 588.900 561.600 ;
        RECT 590.100 549.000 591.900 561.600 ;
        RECT 608.100 549.000 609.900 561.600 ;
        RECT 612.600 549.600 615.900 561.600 ;
        RECT 618.600 549.000 620.400 561.600 ;
        RECT 638.100 549.600 639.900 561.600 ;
        RECT 641.100 560.700 648.900 561.600 ;
        RECT 641.100 549.600 642.900 560.700 ;
        RECT 644.100 549.000 645.900 559.800 ;
        RECT 647.100 549.600 648.900 560.700 ;
        RECT 665.100 550.500 666.900 561.600 ;
        RECT 668.100 551.400 669.900 562.500 ;
        RECT 698.100 561.600 699.300 568.950 ;
        RECT 704.100 567.150 705.900 568.950 ;
        RECT 722.700 561.600 723.600 568.950 ;
        RECT 726.000 567.150 727.800 568.950 ;
        RECT 671.100 560.400 678.900 561.300 ;
        RECT 671.100 550.500 672.900 560.400 ;
        RECT 665.100 549.600 672.900 550.500 ;
        RECT 674.100 549.000 675.900 559.500 ;
        RECT 677.100 549.600 678.900 560.400 ;
        RECT 698.100 560.100 700.500 561.600 ;
        RECT 696.000 557.100 697.800 558.900 ;
        RECT 679.950 552.450 682.050 553.050 ;
        RECT 691.950 552.450 694.050 553.050 ;
        RECT 679.950 551.550 694.050 552.450 ;
        RECT 679.950 550.950 682.050 551.550 ;
        RECT 691.950 550.950 694.050 551.550 ;
        RECT 695.700 549.000 697.500 555.600 ;
        RECT 698.700 549.600 700.500 560.100 ;
        RECT 703.800 549.000 705.600 561.600 ;
        RECT 722.100 549.600 723.900 561.600 ;
        RECT 725.100 549.000 726.900 561.000 ;
        RECT 729.000 555.600 729.900 575.700 ;
        RECT 730.950 571.050 732.750 572.850 ;
        RECT 749.100 571.050 750.900 572.850 ;
        RECT 752.700 571.050 753.900 576.300 ;
        RECT 754.950 571.050 756.750 572.850 ;
        RECT 773.100 571.050 774.900 572.850 ;
        RECT 776.700 571.050 777.900 576.300 ;
        RECT 778.950 571.050 780.750 572.850 ;
        RECT 797.700 571.050 798.900 581.400 ;
        RECT 818.100 578.400 819.900 584.400 ;
        RECT 821.100 579.300 822.900 585.000 ;
        RECT 825.600 578.400 827.400 584.400 ;
        RECT 830.100 579.300 831.900 585.000 ;
        RECT 833.100 578.400 834.900 584.400 ;
        RECT 818.700 576.600 819.900 578.400 ;
        RECT 825.900 576.900 827.100 578.400 ;
        RECT 830.100 577.500 834.900 578.400 ;
        RECT 818.700 575.700 825.000 576.600 ;
        RECT 822.900 573.600 825.000 575.700 ;
        RECT 818.400 571.050 820.200 572.850 ;
        RECT 823.200 571.800 825.000 573.600 ;
        RECT 825.900 574.800 828.900 576.900 ;
        RECT 830.100 576.300 832.200 577.500 ;
        RECT 853.500 576.000 855.300 584.400 ;
        RECT 852.000 574.800 855.300 576.000 ;
        RECT 860.100 575.400 861.900 585.000 ;
        RECT 878.100 575.400 879.900 585.000 ;
        RECT 884.700 576.000 886.500 584.400 ;
        RECT 905.100 578.400 906.900 584.400 ;
        RECT 905.700 576.300 906.900 578.400 ;
        RECT 908.100 579.300 909.900 584.400 ;
        RECT 911.100 580.200 912.900 585.000 ;
        RECT 914.100 579.300 915.900 584.400 ;
        RECT 908.100 577.950 915.900 579.300 ;
        RECT 924.000 576.450 928.050 577.050 ;
        RECT 884.700 574.800 888.000 576.000 ;
        RECT 905.700 575.400 909.300 576.300 ;
        RECT 730.800 568.950 732.900 571.050 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 818.100 570.300 820.200 571.050 ;
        RECT 818.100 568.950 825.000 570.300 ;
        RECT 752.700 555.600 753.900 568.950 ;
        RECT 776.700 555.600 777.900 568.950 ;
        RECT 797.700 555.600 798.900 568.950 ;
        RECT 800.100 567.150 801.900 568.950 ;
        RECT 823.200 568.500 825.000 568.950 ;
        RECT 825.900 569.100 827.100 574.800 ;
        RECT 828.000 571.800 830.100 573.900 ;
        RECT 838.950 573.450 841.050 574.050 ;
        RECT 847.950 573.450 850.050 574.050 ;
        RECT 838.950 572.550 850.050 573.450 ;
        RECT 838.950 571.950 841.050 572.550 ;
        RECT 847.950 571.950 850.050 572.550 ;
        RECT 828.300 570.000 830.100 571.800 ;
        RECT 852.000 571.050 852.900 574.800 ;
        RECT 854.100 571.050 855.900 572.850 ;
        RECT 860.100 571.050 861.900 572.850 ;
        RECT 878.100 571.050 879.900 572.850 ;
        RECT 884.100 571.050 885.900 572.850 ;
        RECT 887.100 571.050 888.000 574.800 ;
        RECT 889.950 573.450 894.000 574.050 ;
        RECT 889.950 573.000 894.450 573.450 ;
        RECT 889.950 571.950 895.050 573.000 ;
        RECT 825.900 568.200 828.300 569.100 ;
        RECT 826.800 568.050 828.300 568.200 ;
        RECT 832.800 568.950 834.900 571.050 ;
        RECT 850.950 568.950 853.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 822.000 565.500 825.900 567.300 ;
        RECT 823.800 565.200 825.900 565.500 ;
        RECT 826.800 565.950 828.900 568.050 ;
        RECT 832.800 567.150 834.600 568.950 ;
        RECT 826.800 564.000 827.700 565.950 ;
        RECT 808.950 561.450 811.050 561.900 ;
        RECT 814.950 561.450 817.050 562.050 ;
        RECT 820.500 561.600 822.600 563.700 ;
        RECT 826.200 562.950 827.700 564.000 ;
        RECT 826.200 561.600 827.400 562.950 ;
        RECT 808.950 560.550 817.050 561.450 ;
        RECT 808.950 559.800 811.050 560.550 ;
        RECT 814.950 559.950 817.050 560.550 ;
        RECT 818.100 560.700 822.600 561.600 ;
        RECT 728.100 549.600 729.900 555.600 ;
        RECT 731.100 549.000 732.900 555.600 ;
        RECT 749.100 549.000 750.900 555.600 ;
        RECT 752.100 549.600 753.900 555.600 ;
        RECT 755.100 549.000 756.900 555.600 ;
        RECT 773.100 549.000 774.900 555.600 ;
        RECT 776.100 549.600 777.900 555.600 ;
        RECT 779.100 549.000 780.900 555.600 ;
        RECT 797.100 549.600 798.900 555.600 ;
        RECT 800.100 549.000 801.900 555.600 ;
        RECT 818.100 549.600 819.900 560.700 ;
        RECT 821.100 549.000 822.900 559.500 ;
        RECT 825.600 549.600 827.400 561.600 ;
        RECT 830.100 561.600 832.200 562.500 ;
        RECT 830.100 560.400 834.900 561.600 ;
        RECT 830.100 549.000 831.900 559.500 ;
        RECT 833.100 549.600 834.900 560.400 ;
        RECT 852.000 556.800 852.900 568.950 ;
        RECT 857.100 567.150 858.900 568.950 ;
        RECT 881.100 567.150 882.900 568.950 ;
        RECT 853.950 564.450 856.050 565.050 ;
        RECT 877.950 564.450 880.050 565.050 ;
        RECT 853.950 563.550 880.050 564.450 ;
        RECT 853.950 562.950 856.050 563.550 ;
        RECT 877.950 562.950 880.050 563.550 ;
        RECT 887.100 556.800 888.000 568.950 ;
        RECT 892.950 568.800 895.050 571.950 ;
        RECT 905.100 571.050 906.900 572.850 ;
        RECT 908.100 571.050 909.300 575.400 ;
        RECT 923.550 574.950 928.050 576.450 ;
        RECT 932.100 575.400 933.900 585.000 ;
        RECT 938.700 576.000 940.500 584.400 ;
        RECT 961.500 576.000 963.300 584.400 ;
        RECT 923.550 573.450 924.450 574.950 ;
        RECT 938.700 574.800 942.000 576.000 ;
        RECT 927.000 573.450 931.050 574.050 ;
        RECT 911.100 571.050 912.900 572.850 ;
        RECT 920.550 572.550 924.450 573.450 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 913.950 568.950 916.050 571.050 ;
        RECT 892.950 564.450 895.050 565.050 ;
        RECT 904.950 564.450 907.050 565.050 ;
        RECT 892.950 563.550 907.050 564.450 ;
        RECT 892.950 562.950 895.050 563.550 ;
        RECT 904.950 562.950 907.050 563.550 ;
        RECT 908.100 561.600 909.300 568.950 ;
        RECT 914.100 567.150 915.900 568.950 ;
        RECT 920.550 568.050 921.450 572.550 ;
        RECT 916.950 566.550 921.450 568.050 ;
        RECT 926.550 571.950 931.050 573.450 ;
        RECT 926.550 568.050 927.450 571.950 ;
        RECT 932.100 571.050 933.900 572.850 ;
        RECT 938.100 571.050 939.900 572.850 ;
        RECT 941.100 571.050 942.000 574.800 ;
        RECT 960.000 574.800 963.300 576.000 ;
        RECT 968.100 575.400 969.900 585.000 ;
        RECT 986.400 578.400 988.200 585.000 ;
        RECT 991.500 577.200 993.300 584.400 ;
        RECT 1010.100 581.400 1011.900 585.000 ;
        RECT 1013.100 581.400 1014.900 584.400 ;
        RECT 1016.100 581.400 1017.900 585.000 ;
        RECT 1034.100 581.400 1035.900 584.400 ;
        RECT 1037.100 581.400 1038.900 585.000 ;
        RECT 989.100 576.300 993.300 577.200 ;
        RECT 960.000 571.050 960.900 574.800 ;
        RECT 982.950 573.450 985.050 574.050 ;
        RECT 962.100 571.050 963.900 572.850 ;
        RECT 968.100 571.050 969.900 572.850 ;
        RECT 974.550 572.550 985.050 573.450 ;
        RECT 931.950 568.950 934.050 571.050 ;
        RECT 934.950 568.950 937.050 571.050 ;
        RECT 937.950 568.950 940.050 571.050 ;
        RECT 940.950 568.950 943.050 571.050 ;
        RECT 958.950 568.950 961.050 571.050 ;
        RECT 961.950 568.950 964.050 571.050 ;
        RECT 964.950 568.950 967.050 571.050 ;
        RECT 967.950 568.950 970.050 571.050 ;
        RECT 926.550 566.550 931.050 568.050 ;
        RECT 935.100 567.150 936.900 568.950 ;
        RECT 916.950 565.950 921.000 566.550 ;
        RECT 927.000 565.950 931.050 566.550 ;
        RECT 910.950 564.450 913.050 565.050 ;
        RECT 922.950 564.450 925.050 565.050 ;
        RECT 934.950 564.450 937.050 565.050 ;
        RECT 910.950 563.550 918.450 564.450 ;
        RECT 910.950 562.950 913.050 563.550 ;
        RECT 908.100 560.100 910.500 561.600 ;
        RECT 906.000 557.100 907.800 558.900 ;
        RECT 852.000 555.900 858.600 556.800 ;
        RECT 852.000 555.600 852.900 555.900 ;
        RECT 851.100 549.600 852.900 555.600 ;
        RECT 857.100 555.600 858.600 555.900 ;
        RECT 881.400 555.900 888.000 556.800 ;
        RECT 881.400 555.600 882.900 555.900 ;
        RECT 854.100 549.000 855.900 555.000 ;
        RECT 857.100 549.600 858.900 555.600 ;
        RECT 860.100 549.000 861.900 555.600 ;
        RECT 878.100 549.000 879.900 555.600 ;
        RECT 881.100 549.600 882.900 555.600 ;
        RECT 887.100 555.600 888.000 555.900 ;
        RECT 884.100 549.000 885.900 555.000 ;
        RECT 887.100 549.600 888.900 555.600 ;
        RECT 905.700 549.000 907.500 555.600 ;
        RECT 908.700 549.600 910.500 560.100 ;
        RECT 913.800 549.000 915.600 561.600 ;
        RECT 917.550 561.450 918.450 563.550 ;
        RECT 922.950 563.550 937.050 564.450 ;
        RECT 922.950 562.950 925.050 563.550 ;
        RECT 934.950 562.950 937.050 563.550 ;
        RECT 931.950 561.450 934.050 561.900 ;
        RECT 917.550 560.550 934.050 561.450 ;
        RECT 931.950 559.800 934.050 560.550 ;
        RECT 941.100 556.800 942.000 568.950 ;
        RECT 935.400 555.900 942.000 556.800 ;
        RECT 935.400 555.600 936.900 555.900 ;
        RECT 932.100 549.000 933.900 555.600 ;
        RECT 935.100 549.600 936.900 555.600 ;
        RECT 941.100 555.600 942.000 555.900 ;
        RECT 960.000 556.800 960.900 568.950 ;
        RECT 965.100 567.150 966.900 568.950 ;
        RECT 974.550 568.050 975.450 572.550 ;
        RECT 982.950 571.950 985.050 572.550 ;
        RECT 986.250 571.050 988.050 572.850 ;
        RECT 989.100 571.050 990.300 576.300 ;
        RECT 994.950 573.450 997.050 574.050 ;
        RECT 992.100 571.050 993.900 572.850 ;
        RECT 994.950 572.550 1005.450 573.450 ;
        RECT 994.950 571.950 997.050 572.550 ;
        RECT 985.950 568.950 988.050 571.050 ;
        RECT 988.950 568.950 991.050 571.050 ;
        RECT 991.950 568.950 994.050 571.050 ;
        RECT 970.950 566.550 975.450 568.050 ;
        RECT 970.950 565.950 975.000 566.550 ;
        RECT 961.950 561.450 964.050 562.050 ;
        RECT 976.950 561.450 979.050 562.050 ;
        RECT 961.950 560.550 979.050 561.450 ;
        RECT 961.950 559.950 964.050 560.550 ;
        RECT 976.950 559.950 979.050 560.550 ;
        RECT 960.000 555.900 966.600 556.800 ;
        RECT 960.000 555.600 960.900 555.900 ;
        RECT 938.100 549.000 939.900 555.000 ;
        RECT 941.100 549.600 942.900 555.600 ;
        RECT 959.100 549.600 960.900 555.600 ;
        RECT 965.100 555.600 966.600 555.900 ;
        RECT 989.100 555.600 990.300 568.950 ;
        RECT 1004.550 568.050 1005.450 572.550 ;
        RECT 1013.700 571.050 1014.600 581.400 ;
        RECT 1034.700 571.050 1035.900 581.400 ;
        RECT 1009.950 568.950 1012.050 571.050 ;
        RECT 1012.950 568.950 1015.050 571.050 ;
        RECT 1015.950 568.950 1018.050 571.050 ;
        RECT 1033.950 568.950 1036.050 571.050 ;
        RECT 1036.950 568.950 1039.050 571.050 ;
        RECT 1004.550 566.550 1009.050 568.050 ;
        RECT 1010.100 567.150 1011.900 568.950 ;
        RECT 1005.000 565.950 1009.050 566.550 ;
        RECT 1013.700 561.600 1014.600 568.950 ;
        RECT 1015.950 567.150 1017.750 568.950 ;
        RECT 1011.000 560.400 1014.600 561.600 ;
        RECT 962.100 549.000 963.900 555.000 ;
        RECT 965.100 549.600 966.900 555.600 ;
        RECT 968.100 549.000 969.900 555.600 ;
        RECT 986.100 549.000 987.900 555.600 ;
        RECT 989.100 549.600 990.900 555.600 ;
        RECT 992.100 549.000 993.900 555.600 ;
        RECT 994.950 552.450 997.050 553.050 ;
        RECT 1000.950 552.450 1003.050 553.050 ;
        RECT 994.950 551.550 1003.050 552.450 ;
        RECT 994.950 550.950 997.050 551.550 ;
        RECT 1000.950 550.950 1003.050 551.550 ;
        RECT 1011.000 549.600 1012.800 560.400 ;
        RECT 1016.100 549.000 1017.900 561.600 ;
        RECT 1034.700 555.600 1035.900 568.950 ;
        RECT 1037.100 567.150 1038.900 568.950 ;
        RECT 1034.100 549.600 1035.900 555.600 ;
        RECT 1037.100 549.000 1038.900 555.600 ;
        RECT 2.700 539.400 4.500 546.000 ;
        RECT 5.700 540.300 7.500 545.400 ;
        RECT 5.400 539.400 7.500 540.300 ;
        RECT 8.700 539.400 10.500 546.000 ;
        RECT 5.400 538.500 6.300 539.400 ;
        RECT 2.700 537.600 6.300 538.500 ;
        RECT 2.700 521.400 3.900 537.600 ;
        RECT 7.200 536.400 9.000 536.700 ;
        RECT 11.700 536.400 13.500 545.400 ;
        RECT 14.700 539.400 16.500 546.000 ;
        RECT 18.300 542.400 20.100 545.400 ;
        RECT 21.300 542.400 23.100 545.400 ;
        RECT 18.300 540.300 20.400 542.400 ;
        RECT 21.300 540.300 23.400 542.400 ;
        RECT 24.300 539.400 26.100 545.400 ;
        RECT 27.300 539.400 29.100 546.000 ;
        RECT 23.700 537.300 25.800 539.400 ;
        RECT 31.200 537.900 33.000 545.400 ;
        RECT 34.200 539.400 36.000 546.000 ;
        RECT 37.200 539.400 39.000 545.400 ;
        RECT 40.200 542.400 42.000 545.400 ;
        RECT 43.200 542.400 45.000 545.400 ;
        RECT 46.200 542.400 48.000 545.400 ;
        RECT 40.200 540.300 42.300 542.400 ;
        RECT 43.200 540.300 45.300 542.400 ;
        RECT 46.200 540.300 48.300 542.400 ;
        RECT 49.200 539.400 51.000 546.000 ;
        RECT 52.200 539.400 54.000 545.400 ;
        RECT 55.200 539.400 57.000 546.000 ;
        RECT 58.200 539.400 60.000 545.400 ;
        RECT 61.200 539.400 63.000 546.000 ;
        RECT 64.500 539.400 66.300 545.400 ;
        RECT 67.500 539.400 69.300 546.000 ;
        RECT 7.200 535.200 26.400 536.400 ;
        RECT 31.200 535.800 34.500 537.900 ;
        RECT 37.200 535.500 39.900 539.400 ;
        RECT 43.200 538.500 45.300 539.400 ;
        RECT 43.200 537.300 51.300 538.500 ;
        RECT 49.500 536.700 51.300 537.300 ;
        RECT 52.200 536.400 53.400 539.400 ;
        RECT 58.800 538.500 60.000 539.400 ;
        RECT 58.800 537.600 62.700 538.500 ;
        RECT 56.100 536.400 57.900 537.000 ;
        RECT 7.200 534.900 9.000 535.200 ;
        RECT 25.200 534.600 26.400 535.200 ;
        RECT 40.800 534.600 42.900 535.500 ;
        RECT 10.500 533.700 12.300 534.300 ;
        RECT 20.400 533.700 22.500 534.300 ;
        RECT 10.500 532.500 22.500 533.700 ;
        RECT 25.200 533.400 42.900 534.600 ;
        RECT 46.200 534.300 48.300 535.500 ;
        RECT 52.200 535.200 57.900 536.400 ;
        RECT 61.800 534.300 62.700 537.600 ;
        RECT 46.200 533.400 62.700 534.300 ;
        RECT 20.400 532.200 22.500 532.500 ;
        RECT 25.200 531.300 60.900 532.500 ;
        RECT 25.200 530.700 26.400 531.300 ;
        RECT 59.100 530.700 60.900 531.300 ;
        RECT 12.900 529.800 26.400 530.700 ;
        RECT 37.800 529.800 39.900 530.100 ;
        RECT 12.900 529.050 14.700 529.800 ;
        RECT 4.800 526.950 6.900 529.050 ;
        RECT 10.800 527.250 14.700 529.050 ;
        RECT 32.400 528.300 34.500 529.200 ;
        RECT 10.800 526.950 12.900 527.250 ;
        RECT 23.400 527.100 34.500 528.300 ;
        RECT 36.000 528.000 39.900 529.800 ;
        RECT 44.100 528.300 45.900 530.100 ;
        RECT 45.000 527.100 45.900 528.300 ;
        RECT 5.100 525.300 6.900 526.950 ;
        RECT 23.400 526.500 25.200 527.100 ;
        RECT 32.400 526.200 45.900 527.100 ;
        RECT 48.600 526.800 53.700 528.600 ;
        RECT 55.800 526.950 57.900 529.050 ;
        RECT 48.600 525.300 49.500 526.800 ;
        RECT 5.100 524.100 49.500 525.300 ;
        RECT 55.800 524.100 57.300 526.950 ;
        RECT 20.400 521.400 22.200 523.200 ;
        RECT 28.800 522.000 30.900 523.050 ;
        RECT 50.700 522.600 57.300 524.100 ;
        RECT 2.700 520.200 19.500 521.400 ;
        RECT 2.700 516.600 3.900 520.200 ;
        RECT 17.400 519.300 19.500 520.200 ;
        RECT 6.900 518.700 8.700 519.300 ;
        RECT 6.900 517.500 15.300 518.700 ;
        RECT 13.800 516.600 15.300 517.500 ;
        RECT 20.400 518.400 21.300 521.400 ;
        RECT 25.800 521.100 30.900 522.000 ;
        RECT 25.800 520.200 27.600 521.100 ;
        RECT 28.800 520.950 30.900 521.100 ;
        RECT 35.100 521.100 52.200 522.600 ;
        RECT 35.100 520.500 37.200 521.100 ;
        RECT 35.100 518.700 36.900 520.500 ;
        RECT 53.100 519.900 60.900 521.700 ;
        RECT 20.400 517.200 27.600 518.400 ;
        RECT 22.800 516.600 24.600 517.200 ;
        RECT 26.700 516.600 27.600 517.200 ;
        RECT 42.300 516.600 48.900 518.400 ;
        RECT 53.100 516.600 54.600 519.900 ;
        RECT 61.800 516.600 62.700 533.400 ;
        RECT 2.700 510.600 4.500 516.600 ;
        RECT 8.100 510.000 9.900 516.600 ;
        RECT 13.500 510.600 15.300 516.600 ;
        RECT 17.700 513.600 19.800 515.700 ;
        RECT 20.700 513.600 22.800 515.700 ;
        RECT 23.700 513.600 25.800 515.700 ;
        RECT 26.700 515.400 29.400 516.600 ;
        RECT 27.600 514.500 29.400 515.400 ;
        RECT 31.200 514.500 33.900 516.600 ;
        RECT 17.700 510.600 19.500 513.600 ;
        RECT 20.700 510.600 22.500 513.600 ;
        RECT 23.700 510.600 25.500 513.600 ;
        RECT 26.700 510.000 28.500 513.600 ;
        RECT 31.200 510.600 33.000 514.500 ;
        RECT 37.200 513.600 39.300 515.700 ;
        RECT 40.200 513.600 42.300 515.700 ;
        RECT 43.200 513.600 45.300 515.700 ;
        RECT 46.200 513.600 48.300 515.700 ;
        RECT 50.400 515.400 54.600 516.600 ;
        RECT 34.200 510.000 36.000 513.600 ;
        RECT 37.200 510.600 39.000 513.600 ;
        RECT 40.200 510.600 42.000 513.600 ;
        RECT 43.200 510.600 45.000 513.600 ;
        RECT 46.200 510.600 48.000 513.600 ;
        RECT 50.400 510.600 52.200 515.400 ;
        RECT 55.500 510.000 57.300 516.600 ;
        RECT 60.900 510.600 62.700 516.600 ;
        RECT 64.500 529.050 66.000 539.400 ;
        RECT 86.100 533.400 87.900 545.400 ;
        RECT 89.100 534.300 90.900 545.400 ;
        RECT 92.100 535.200 93.900 546.000 ;
        RECT 95.100 534.300 96.900 545.400 ;
        RECT 113.100 539.400 114.900 546.000 ;
        RECT 116.100 539.400 117.900 545.400 ;
        RECT 89.100 533.400 96.900 534.300 ;
        RECT 64.500 526.950 66.900 529.050 ;
        RECT 64.500 513.600 66.000 526.950 ;
        RECT 86.400 526.050 87.300 533.400 ;
        RECT 88.950 531.450 91.050 532.050 ;
        RECT 112.950 531.450 115.050 532.050 ;
        RECT 88.950 530.550 115.050 531.450 ;
        RECT 88.950 529.950 91.050 530.550 ;
        RECT 112.950 529.950 115.050 530.550 ;
        RECT 91.950 526.050 93.750 527.850 ;
        RECT 113.100 526.050 114.900 527.850 ;
        RECT 116.100 526.050 117.300 539.400 ;
        RECT 134.100 533.400 135.900 545.400 ;
        RECT 137.100 534.300 138.900 545.400 ;
        RECT 140.100 535.200 141.900 546.000 ;
        RECT 143.100 534.300 144.900 545.400 ;
        RECT 161.100 539.400 162.900 546.000 ;
        RECT 164.100 539.400 165.900 545.400 ;
        RECT 182.100 539.400 183.900 546.000 ;
        RECT 185.100 539.400 186.900 545.400 ;
        RECT 188.100 539.400 189.900 546.000 ;
        RECT 193.950 543.450 196.050 544.050 ;
        RECT 202.950 543.450 205.050 544.050 ;
        RECT 193.950 542.550 205.050 543.450 ;
        RECT 193.950 541.950 196.050 542.550 ;
        RECT 202.950 541.950 205.050 542.550 ;
        RECT 137.100 533.400 144.900 534.300 ;
        RECT 134.400 526.050 135.300 533.400 ;
        RECT 139.950 526.050 141.750 527.850 ;
        RECT 161.100 526.050 162.900 527.850 ;
        RECT 164.100 526.050 165.300 539.400 ;
        RECT 177.000 528.450 181.050 529.050 ;
        RECT 176.550 526.950 181.050 528.450 ;
        RECT 85.950 523.950 88.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 86.400 516.600 87.300 523.950 ;
        RECT 88.950 522.150 90.750 523.950 ;
        RECT 95.100 522.150 96.900 523.950 ;
        RECT 86.400 515.400 91.500 516.600 ;
        RECT 64.500 510.600 66.300 513.600 ;
        RECT 67.500 510.000 69.300 513.600 ;
        RECT 86.700 510.000 88.500 513.600 ;
        RECT 89.700 510.600 91.500 515.400 ;
        RECT 94.200 510.000 96.000 516.600 ;
        RECT 116.100 513.600 117.300 523.950 ;
        RECT 134.400 516.600 135.300 523.950 ;
        RECT 136.950 522.150 138.750 523.950 ;
        RECT 143.100 522.150 144.900 523.950 ;
        RECT 134.400 515.400 139.500 516.600 ;
        RECT 113.100 510.000 114.900 513.600 ;
        RECT 116.100 510.600 117.900 513.600 ;
        RECT 134.700 510.000 136.500 513.600 ;
        RECT 137.700 510.600 139.500 515.400 ;
        RECT 142.200 510.000 144.000 516.600 ;
        RECT 164.100 513.600 165.300 523.950 ;
        RECT 176.550 523.050 177.450 526.950 ;
        RECT 185.700 526.050 186.900 539.400 ;
        RECT 206.400 533.400 208.200 546.000 ;
        RECT 211.500 534.900 213.300 545.400 ;
        RECT 214.500 539.400 216.300 546.000 ;
        RECT 233.100 539.400 234.900 546.000 ;
        RECT 236.100 539.400 237.900 545.400 ;
        RECT 239.100 540.000 240.900 546.000 ;
        RECT 236.400 539.100 237.900 539.400 ;
        RECT 242.100 539.400 243.900 545.400 ;
        RECT 242.100 539.100 243.000 539.400 ;
        RECT 236.400 538.200 243.000 539.100 ;
        RECT 214.200 536.100 216.000 537.900 ;
        RECT 211.500 533.400 213.900 534.900 ;
        RECT 206.100 526.050 207.900 527.850 ;
        RECT 212.700 526.050 213.900 533.400 ;
        RECT 217.950 528.450 220.050 529.050 ;
        RECT 226.950 528.450 229.050 529.050 ;
        RECT 217.950 527.550 229.050 528.450 ;
        RECT 217.950 526.950 220.050 527.550 ;
        RECT 226.950 526.950 229.050 527.550 ;
        RECT 236.100 526.050 237.900 527.850 ;
        RECT 242.100 526.050 243.000 538.200 ;
        RECT 260.100 533.400 261.900 546.000 ;
        RECT 265.200 534.600 267.000 545.400 ;
        RECT 271.950 540.450 274.050 541.050 ;
        RECT 280.950 540.450 283.050 541.050 ;
        RECT 271.950 539.550 283.050 540.450 ;
        RECT 271.950 538.950 274.050 539.550 ;
        RECT 280.950 538.950 283.050 539.550 ;
        RECT 263.400 533.400 267.000 534.600 ;
        RECT 284.100 534.600 285.900 545.400 ;
        RECT 287.100 535.500 288.900 546.000 ;
        RECT 290.100 544.500 297.900 545.400 ;
        RECT 290.100 534.600 291.900 544.500 ;
        RECT 284.100 533.700 291.900 534.600 ;
        RECT 260.250 526.050 262.050 527.850 ;
        RECT 263.400 526.050 264.300 533.400 ;
        RECT 293.100 532.500 294.900 543.600 ;
        RECT 296.100 533.400 297.900 544.500 ;
        RECT 314.100 539.400 315.900 545.400 ;
        RECT 317.100 540.000 318.900 546.000 ;
        RECT 315.000 539.100 315.900 539.400 ;
        RECT 320.100 539.400 321.900 545.400 ;
        RECT 323.100 539.400 324.900 546.000 ;
        RECT 320.100 539.100 321.600 539.400 ;
        RECT 315.000 538.200 321.600 539.100 ;
        RECT 290.100 531.600 294.900 532.500 ;
        RECT 266.100 526.050 267.900 527.850 ;
        RECT 287.250 526.050 289.050 527.850 ;
        RECT 290.100 526.050 291.000 531.600 ;
        RECT 293.100 526.050 294.900 527.850 ;
        RECT 315.000 526.050 315.900 538.200 ;
        RECT 319.950 534.450 322.050 535.050 ;
        RECT 337.950 534.450 340.050 535.050 ;
        RECT 319.950 533.550 340.050 534.450 ;
        RECT 319.950 532.950 322.050 533.550 ;
        RECT 337.950 532.950 340.050 533.550 ;
        RECT 342.000 534.600 343.800 545.400 ;
        RECT 342.000 533.400 345.600 534.600 ;
        RECT 347.100 533.400 348.900 546.000 ;
        RECT 365.100 539.400 366.900 546.000 ;
        RECT 368.100 539.400 369.900 545.400 ;
        RECT 320.100 526.050 321.900 527.850 ;
        RECT 341.100 526.050 342.900 527.850 ;
        RECT 344.700 526.050 345.600 533.400 ;
        RECT 346.950 526.050 348.750 527.850 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 211.950 523.950 214.050 526.050 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 343.950 523.950 346.050 526.050 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 365.100 523.950 367.200 526.050 ;
        RECT 176.550 521.550 181.050 523.050 ;
        RECT 182.100 522.150 183.900 523.950 ;
        RECT 177.000 520.950 181.050 521.550 ;
        RECT 185.700 518.700 186.900 523.950 ;
        RECT 187.950 522.150 189.750 523.950 ;
        RECT 209.100 522.150 210.900 523.950 ;
        RECT 212.700 519.600 213.900 523.950 ;
        RECT 215.100 522.150 216.900 523.950 ;
        RECT 233.100 522.150 234.900 523.950 ;
        RECT 239.100 522.150 240.900 523.950 ;
        RECT 242.100 520.200 243.000 523.950 ;
        RECT 212.700 518.700 216.300 519.600 ;
        RECT 182.700 517.800 186.900 518.700 ;
        RECT 161.100 510.000 162.900 513.600 ;
        RECT 164.100 510.600 165.900 513.600 ;
        RECT 182.700 510.600 184.500 517.800 ;
        RECT 187.800 510.000 189.600 516.600 ;
        RECT 206.100 515.700 213.900 517.050 ;
        RECT 206.100 510.600 207.900 515.700 ;
        RECT 209.100 510.000 210.900 514.800 ;
        RECT 212.100 510.600 213.900 515.700 ;
        RECT 215.100 516.600 216.300 518.700 ;
        RECT 215.100 510.600 216.900 516.600 ;
        RECT 233.100 510.000 234.900 519.600 ;
        RECT 239.700 519.000 243.000 520.200 ;
        RECT 239.700 510.600 241.500 519.000 ;
        RECT 263.400 513.600 264.300 523.950 ;
        RECT 284.250 522.150 286.050 523.950 ;
        RECT 290.100 516.600 291.300 523.950 ;
        RECT 296.100 522.150 297.900 523.950 ;
        RECT 304.950 522.450 307.050 523.050 ;
        RECT 310.950 522.450 313.050 523.050 ;
        RECT 304.950 521.550 313.050 522.450 ;
        RECT 304.950 520.950 307.050 521.550 ;
        RECT 310.950 520.950 313.050 521.550 ;
        RECT 315.000 520.200 315.900 523.950 ;
        RECT 317.100 522.150 318.900 523.950 ;
        RECT 323.100 522.150 324.900 523.950 ;
        RECT 315.000 519.000 318.300 520.200 ;
        RECT 260.100 510.000 261.900 513.600 ;
        RECT 263.100 510.600 264.900 513.600 ;
        RECT 266.100 510.000 267.900 513.600 ;
        RECT 284.700 510.000 286.500 516.600 ;
        RECT 289.200 510.600 291.000 516.600 ;
        RECT 293.700 510.000 295.500 516.600 ;
        RECT 316.500 510.600 318.300 519.000 ;
        RECT 323.100 510.000 324.900 519.600 ;
        RECT 344.700 513.600 345.600 523.950 ;
        RECT 365.250 522.150 367.050 523.950 ;
        RECT 368.100 519.300 369.000 539.400 ;
        RECT 371.100 534.000 372.900 546.000 ;
        RECT 374.100 533.400 375.900 545.400 ;
        RECT 392.100 539.400 393.900 545.400 ;
        RECT 395.100 540.000 396.900 546.000 ;
        RECT 393.000 539.100 393.900 539.400 ;
        RECT 398.100 539.400 399.900 545.400 ;
        RECT 401.100 539.400 402.900 546.000 ;
        RECT 419.700 539.400 421.500 546.000 ;
        RECT 398.100 539.100 399.600 539.400 ;
        RECT 393.000 538.200 399.600 539.100 ;
        RECT 370.200 526.050 372.000 527.850 ;
        RECT 374.400 526.050 375.300 533.400 ;
        RECT 393.000 526.050 393.900 538.200 ;
        RECT 420.000 536.100 421.800 537.900 ;
        RECT 412.950 534.450 415.050 535.050 ;
        RECT 418.950 534.450 421.050 535.050 ;
        RECT 422.700 534.900 424.500 545.400 ;
        RECT 412.950 533.550 421.050 534.450 ;
        RECT 412.950 532.950 415.050 533.550 ;
        RECT 418.950 532.950 421.050 533.550 ;
        RECT 422.100 533.400 424.500 534.900 ;
        RECT 427.800 533.400 429.600 546.000 ;
        RECT 446.100 539.400 447.900 546.000 ;
        RECT 449.100 539.400 450.900 545.400 ;
        RECT 398.100 526.050 399.900 527.850 ;
        RECT 422.100 526.050 423.300 533.400 ;
        RECT 428.100 526.050 429.900 527.850 ;
        RECT 446.100 526.050 447.900 527.850 ;
        RECT 449.100 526.050 450.300 539.400 ;
        RECT 467.100 533.400 468.900 545.400 ;
        RECT 470.100 534.300 471.900 545.400 ;
        RECT 473.100 535.200 474.900 546.000 ;
        RECT 476.100 534.300 477.900 545.400 ;
        RECT 494.700 539.400 496.500 546.000 ;
        RECT 495.000 536.100 496.800 537.900 ;
        RECT 497.700 534.900 499.500 545.400 ;
        RECT 470.100 533.400 477.900 534.300 ;
        RECT 497.100 533.400 499.500 534.900 ;
        RECT 502.800 533.400 504.600 546.000 ;
        RECT 521.700 539.400 523.500 546.000 ;
        RECT 522.000 536.100 523.800 537.900 ;
        RECT 524.700 534.900 526.500 545.400 ;
        RECT 524.100 533.400 526.500 534.900 ;
        RECT 529.800 533.400 531.600 546.000 ;
        RECT 533.700 539.400 535.500 546.000 ;
        RECT 536.700 539.400 538.500 545.400 ;
        RECT 540.000 539.400 541.800 546.000 ;
        RECT 543.000 539.400 544.800 545.400 ;
        RECT 546.000 539.400 547.800 546.000 ;
        RECT 549.000 539.400 550.800 545.400 ;
        RECT 552.000 539.400 553.800 546.000 ;
        RECT 555.000 542.400 556.800 545.400 ;
        RECT 558.000 542.400 559.800 545.400 ;
        RECT 561.000 542.400 562.800 545.400 ;
        RECT 554.700 540.300 556.800 542.400 ;
        RECT 557.700 540.300 559.800 542.400 ;
        RECT 560.700 540.300 562.800 542.400 ;
        RECT 564.000 539.400 565.800 545.400 ;
        RECT 567.000 539.400 568.800 546.000 ;
        RECT 467.400 526.050 468.300 533.400 ;
        RECT 472.950 526.050 474.750 527.850 ;
        RECT 497.100 526.050 498.300 533.400 ;
        RECT 499.950 531.450 502.050 532.050 ;
        RECT 511.950 531.450 514.050 532.050 ;
        RECT 499.950 530.550 514.050 531.450 ;
        RECT 499.950 529.950 502.050 530.550 ;
        RECT 511.950 529.950 514.050 530.550 ;
        RECT 503.100 526.050 504.900 527.850 ;
        RECT 524.100 526.050 525.300 533.400 ;
        RECT 537.000 529.050 538.500 539.400 ;
        RECT 543.000 538.500 544.200 539.400 ;
        RECT 530.100 526.050 531.900 527.850 ;
        RECT 536.100 526.950 538.500 529.050 ;
        RECT 370.500 523.950 372.600 526.050 ;
        RECT 373.800 523.950 375.900 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 397.950 523.950 400.050 526.050 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 448.950 523.950 451.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 475.950 523.950 478.050 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 365.100 518.400 373.500 519.300 ;
        RECT 341.100 510.000 342.900 513.600 ;
        RECT 344.100 510.600 345.900 513.600 ;
        RECT 347.100 510.000 348.900 513.600 ;
        RECT 365.100 510.600 366.900 518.400 ;
        RECT 371.700 517.500 373.500 518.400 ;
        RECT 374.400 516.600 375.300 523.950 ;
        RECT 393.000 520.200 393.900 523.950 ;
        RECT 395.100 522.150 396.900 523.950 ;
        RECT 401.100 522.150 402.900 523.950 ;
        RECT 419.100 522.150 420.900 523.950 ;
        RECT 393.000 519.000 396.300 520.200 ;
        RECT 422.100 519.600 423.300 523.950 ;
        RECT 425.100 522.150 426.900 523.950 ;
        RECT 369.600 510.000 371.400 516.600 ;
        RECT 372.600 514.800 375.300 516.600 ;
        RECT 372.600 510.600 374.400 514.800 ;
        RECT 394.500 510.600 396.300 519.000 ;
        RECT 401.100 510.000 402.900 519.600 ;
        RECT 419.700 518.700 423.300 519.600 ;
        RECT 419.700 516.600 420.900 518.700 ;
        RECT 419.100 510.600 420.900 516.600 ;
        RECT 422.100 515.700 429.900 517.050 ;
        RECT 422.100 510.600 423.900 515.700 ;
        RECT 425.100 510.000 426.900 514.800 ;
        RECT 428.100 510.600 429.900 515.700 ;
        RECT 449.100 513.600 450.300 523.950 ;
        RECT 467.400 516.600 468.300 523.950 ;
        RECT 469.950 522.150 471.750 523.950 ;
        RECT 476.100 522.150 477.900 523.950 ;
        RECT 478.950 522.450 481.050 523.050 ;
        RECT 484.950 522.450 487.050 523.050 ;
        RECT 478.950 521.550 487.050 522.450 ;
        RECT 494.100 522.150 495.900 523.950 ;
        RECT 478.950 520.950 481.050 521.550 ;
        RECT 484.950 520.950 487.050 521.550 ;
        RECT 469.950 519.450 472.050 520.050 ;
        RECT 481.950 519.450 484.050 519.900 ;
        RECT 497.100 519.600 498.300 523.950 ;
        RECT 500.100 522.150 501.900 523.950 ;
        RECT 521.100 522.150 522.900 523.950 ;
        RECT 524.100 519.600 525.300 523.950 ;
        RECT 527.100 522.150 528.900 523.950 ;
        RECT 469.950 518.550 484.050 519.450 ;
        RECT 469.950 517.950 472.050 518.550 ;
        RECT 481.950 517.800 484.050 518.550 ;
        RECT 494.700 518.700 498.300 519.600 ;
        RECT 521.700 518.700 525.300 519.600 ;
        RECT 494.700 516.600 495.900 518.700 ;
        RECT 467.400 515.400 472.500 516.600 ;
        RECT 446.100 510.000 447.900 513.600 ;
        RECT 449.100 510.600 450.900 513.600 ;
        RECT 467.700 510.000 469.500 513.600 ;
        RECT 470.700 510.600 472.500 515.400 ;
        RECT 475.200 510.000 477.000 516.600 ;
        RECT 494.100 510.600 495.900 516.600 ;
        RECT 497.100 515.700 504.900 517.050 ;
        RECT 521.700 516.600 522.900 518.700 ;
        RECT 497.100 510.600 498.900 515.700 ;
        RECT 500.100 510.000 501.900 514.800 ;
        RECT 503.100 510.600 504.900 515.700 ;
        RECT 521.100 510.600 522.900 516.600 ;
        RECT 524.100 515.700 531.900 517.050 ;
        RECT 524.100 510.600 525.900 515.700 ;
        RECT 527.100 510.000 528.900 514.800 ;
        RECT 530.100 510.600 531.900 515.700 ;
        RECT 537.000 513.600 538.500 526.950 ;
        RECT 533.700 510.000 535.500 513.600 ;
        RECT 536.700 510.600 538.500 513.600 ;
        RECT 540.300 537.600 544.200 538.500 ;
        RECT 540.300 534.300 541.200 537.600 ;
        RECT 545.100 536.400 546.900 537.000 ;
        RECT 549.600 536.400 550.800 539.400 ;
        RECT 557.700 538.500 559.800 539.400 ;
        RECT 551.700 537.300 559.800 538.500 ;
        RECT 551.700 536.700 553.500 537.300 ;
        RECT 545.100 535.200 550.800 536.400 ;
        RECT 563.100 535.500 565.800 539.400 ;
        RECT 570.000 537.900 571.800 545.400 ;
        RECT 573.900 539.400 575.700 546.000 ;
        RECT 576.900 539.400 578.700 545.400 ;
        RECT 579.900 542.400 581.700 545.400 ;
        RECT 582.900 542.400 584.700 545.400 ;
        RECT 579.600 540.300 581.700 542.400 ;
        RECT 582.600 540.300 584.700 542.400 ;
        RECT 586.500 539.400 588.300 546.000 ;
        RECT 568.500 535.800 571.800 537.900 ;
        RECT 577.200 537.300 579.300 539.400 ;
        RECT 589.500 536.400 591.300 545.400 ;
        RECT 592.500 539.400 594.300 546.000 ;
        RECT 595.500 540.300 597.300 545.400 ;
        RECT 595.500 539.400 597.600 540.300 ;
        RECT 598.500 539.400 600.300 546.000 ;
        RECT 596.700 538.500 597.600 539.400 ;
        RECT 596.700 537.600 600.300 538.500 ;
        RECT 594.000 536.400 595.800 536.700 ;
        RECT 554.700 534.300 556.800 535.500 ;
        RECT 540.300 533.400 556.800 534.300 ;
        RECT 560.100 534.600 562.200 535.500 ;
        RECT 576.600 535.200 595.800 536.400 ;
        RECT 576.600 534.600 577.800 535.200 ;
        RECT 594.000 534.900 595.800 535.200 ;
        RECT 560.100 533.400 577.800 534.600 ;
        RECT 580.500 533.700 582.600 534.300 ;
        RECT 590.700 533.700 592.500 534.300 ;
        RECT 540.300 516.600 541.200 533.400 ;
        RECT 580.500 532.500 592.500 533.700 ;
        RECT 542.100 531.300 577.800 532.500 ;
        RECT 580.500 532.200 582.600 532.500 ;
        RECT 542.100 530.700 543.900 531.300 ;
        RECT 576.600 530.700 577.800 531.300 ;
        RECT 545.100 526.950 547.200 529.050 ;
        RECT 545.700 524.100 547.200 526.950 ;
        RECT 549.300 526.800 554.400 528.600 ;
        RECT 553.500 525.300 554.400 526.800 ;
        RECT 557.100 528.300 558.900 530.100 ;
        RECT 563.100 529.800 565.200 530.100 ;
        RECT 576.600 529.800 590.100 530.700 ;
        RECT 557.100 527.100 558.000 528.300 ;
        RECT 563.100 528.000 567.000 529.800 ;
        RECT 568.500 528.300 570.600 529.200 ;
        RECT 588.300 529.050 590.100 529.800 ;
        RECT 568.500 527.100 579.600 528.300 ;
        RECT 588.300 527.250 592.200 529.050 ;
        RECT 557.100 526.200 570.600 527.100 ;
        RECT 577.800 526.500 579.600 527.100 ;
        RECT 590.100 526.950 592.200 527.250 ;
        RECT 596.100 526.950 598.200 529.050 ;
        RECT 596.100 525.300 597.900 526.950 ;
        RECT 553.500 524.100 597.900 525.300 ;
        RECT 545.700 522.600 552.300 524.100 ;
        RECT 542.100 519.900 549.900 521.700 ;
        RECT 550.800 521.100 567.900 522.600 ;
        RECT 565.800 520.500 567.900 521.100 ;
        RECT 572.100 522.000 574.200 523.050 ;
        RECT 572.100 521.100 577.200 522.000 ;
        RECT 580.800 521.400 582.600 523.200 ;
        RECT 599.100 521.400 600.300 537.600 ;
        RECT 617.100 534.600 618.900 545.400 ;
        RECT 620.100 535.500 621.900 546.000 ;
        RECT 617.100 533.400 621.900 534.600 ;
        RECT 619.800 532.500 621.900 533.400 ;
        RECT 624.600 533.400 626.400 545.400 ;
        RECT 629.100 535.500 630.900 546.000 ;
        RECT 632.100 534.300 633.900 545.400 ;
        RECT 629.400 533.400 633.900 534.300 ;
        RECT 650.100 534.600 651.900 545.400 ;
        RECT 653.100 535.500 654.900 546.000 ;
        RECT 656.100 544.500 663.900 545.400 ;
        RECT 656.100 534.600 657.900 544.500 ;
        RECT 650.100 533.700 657.900 534.600 ;
        RECT 624.600 532.050 625.800 533.400 ;
        RECT 624.300 531.000 625.800 532.050 ;
        RECT 629.400 531.300 631.500 533.400 ;
        RECT 659.100 532.500 660.900 543.600 ;
        RECT 662.100 533.400 663.900 544.500 ;
        RECT 680.700 539.400 682.500 546.000 ;
        RECT 681.000 536.100 682.800 537.900 ;
        RECT 683.700 534.900 685.500 545.400 ;
        RECT 683.100 533.400 685.500 534.900 ;
        RECT 688.800 533.400 690.600 546.000 ;
        RECT 691.950 540.450 694.050 541.050 ;
        RECT 703.950 540.450 706.050 540.900 ;
        RECT 691.950 539.550 706.050 540.450 ;
        RECT 691.950 538.950 694.050 539.550 ;
        RECT 703.950 538.800 706.050 539.550 ;
        RECT 708.600 533.400 710.400 546.000 ;
        RECT 713.100 533.400 716.400 545.400 ;
        RECT 719.100 533.400 720.900 546.000 ;
        RECT 737.100 534.300 738.900 545.400 ;
        RECT 740.100 535.500 741.900 546.000 ;
        RECT 737.100 533.400 741.600 534.300 ;
        RECT 744.600 533.400 746.400 545.400 ;
        RECT 749.100 535.500 750.900 546.000 ;
        RECT 752.100 534.600 753.900 545.400 ;
        RECT 771.600 534.900 773.400 545.400 ;
        RECT 656.100 531.600 660.900 532.500 ;
        RECT 624.300 529.050 625.200 531.000 ;
        RECT 617.400 526.050 619.200 527.850 ;
        RECT 623.100 526.950 625.200 529.050 ;
        RECT 626.100 529.500 628.200 529.800 ;
        RECT 626.100 527.700 630.000 529.500 ;
        RECT 617.100 523.950 619.200 526.050 ;
        RECT 623.700 526.800 625.200 526.950 ;
        RECT 623.700 525.900 626.100 526.800 ;
        RECT 572.100 520.950 574.200 521.100 ;
        RECT 548.400 516.600 549.900 519.900 ;
        RECT 566.100 518.700 567.900 520.500 ;
        RECT 575.400 520.200 577.200 521.100 ;
        RECT 581.700 518.400 582.600 521.400 ;
        RECT 583.500 520.200 600.300 521.400 ;
        RECT 621.900 523.200 623.700 525.000 ;
        RECT 621.900 521.100 624.000 523.200 ;
        RECT 624.900 520.200 626.100 525.900 ;
        RECT 627.000 526.050 628.800 526.500 ;
        RECT 653.250 526.050 655.050 527.850 ;
        RECT 656.100 526.050 657.000 531.600 ;
        RECT 667.950 531.450 670.050 532.050 ;
        RECT 676.950 531.450 679.050 532.050 ;
        RECT 667.950 530.550 679.050 531.450 ;
        RECT 667.950 529.950 670.050 530.550 ;
        RECT 676.950 529.950 679.050 530.550 ;
        RECT 664.950 528.450 667.050 529.050 ;
        RECT 659.100 526.050 660.900 527.850 ;
        RECT 664.950 527.550 672.450 528.450 ;
        RECT 664.950 526.950 667.050 527.550 ;
        RECT 627.000 524.700 633.900 526.050 ;
        RECT 631.800 523.950 633.900 524.700 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 671.550 525.450 672.450 527.550 ;
        RECT 683.100 526.050 684.300 533.400 ;
        RECT 685.950 531.450 688.050 532.050 ;
        RECT 694.950 531.450 697.050 532.050 ;
        RECT 685.950 530.550 697.050 531.450 ;
        RECT 685.950 529.950 688.050 530.550 ;
        RECT 694.950 529.950 697.050 530.550 ;
        RECT 689.100 526.050 690.900 527.850 ;
        RECT 707.250 526.050 709.050 527.850 ;
        RECT 714.000 526.050 715.050 533.400 ;
        RECT 718.950 531.450 721.050 531.900 ;
        RECT 733.950 531.450 736.050 532.050 ;
        RECT 718.950 530.550 736.050 531.450 ;
        RECT 739.500 531.300 741.600 533.400 ;
        RECT 745.200 532.050 746.400 533.400 ;
        RECT 749.100 533.400 753.900 534.600 ;
        RECT 771.000 533.400 773.400 534.900 ;
        RECT 774.600 533.400 776.400 546.000 ;
        RECT 779.100 533.400 780.900 545.400 ;
        RECT 797.100 533.400 798.900 546.000 ;
        RECT 802.200 534.600 804.000 545.400 ;
        RECT 800.400 533.400 804.000 534.600 ;
        RECT 821.100 533.400 822.900 545.400 ;
        RECT 824.100 534.300 825.900 545.400 ;
        RECT 827.100 535.200 828.900 546.000 ;
        RECT 830.100 534.300 831.900 545.400 ;
        RECT 824.100 533.400 831.900 534.300 ;
        RECT 848.100 533.400 849.900 546.000 ;
        RECT 853.200 534.600 855.000 545.400 ;
        RECT 872.100 539.400 873.900 546.000 ;
        RECT 875.100 539.400 876.900 545.400 ;
        RECT 878.100 539.400 879.900 546.000 ;
        RECT 896.100 539.400 897.900 546.000 ;
        RECT 899.100 539.400 900.900 545.400 ;
        RECT 902.100 540.000 903.900 546.000 ;
        RECT 851.400 533.400 855.000 534.600 ;
        RECT 749.100 532.500 751.200 533.400 ;
        RECT 745.200 531.000 746.700 532.050 ;
        RECT 718.950 529.800 721.050 530.550 ;
        RECT 733.950 529.950 736.050 530.550 ;
        RECT 742.800 529.500 744.900 529.800 ;
        RECT 719.100 526.050 720.900 527.850 ;
        RECT 741.000 527.700 744.900 529.500 ;
        RECT 745.800 529.050 746.700 531.000 ;
        RECT 745.800 526.950 747.900 529.050 ;
        RECT 745.800 526.800 747.300 526.950 ;
        RECT 742.200 526.050 744.000 526.500 ;
        RECT 671.550 524.550 675.450 525.450 ;
        RECT 583.500 519.300 585.600 520.200 ;
        RECT 594.300 518.700 596.100 519.300 ;
        RECT 554.100 516.600 560.700 518.400 ;
        RECT 575.400 517.200 582.600 518.400 ;
        RECT 587.700 517.500 596.100 518.700 ;
        RECT 575.400 516.600 576.300 517.200 ;
        RECT 578.400 516.600 580.200 517.200 ;
        RECT 587.700 516.600 589.200 517.500 ;
        RECT 599.100 516.600 600.300 520.200 ;
        RECT 619.800 517.500 621.900 518.700 ;
        RECT 623.100 518.100 626.100 520.200 ;
        RECT 627.000 521.400 628.800 523.200 ;
        RECT 631.800 522.150 633.600 523.950 ;
        RECT 650.250 522.150 652.050 523.950 ;
        RECT 627.000 519.300 629.100 521.400 ;
        RECT 627.000 518.400 633.300 519.300 ;
        RECT 540.300 510.600 542.100 516.600 ;
        RECT 545.700 510.000 547.500 516.600 ;
        RECT 548.400 515.400 552.600 516.600 ;
        RECT 550.800 510.600 552.600 515.400 ;
        RECT 554.700 513.600 556.800 515.700 ;
        RECT 557.700 513.600 559.800 515.700 ;
        RECT 560.700 513.600 562.800 515.700 ;
        RECT 563.700 513.600 565.800 515.700 ;
        RECT 569.100 514.500 571.800 516.600 ;
        RECT 573.600 515.400 576.300 516.600 ;
        RECT 573.600 514.500 575.400 515.400 ;
        RECT 555.000 510.600 556.800 513.600 ;
        RECT 558.000 510.600 559.800 513.600 ;
        RECT 561.000 510.600 562.800 513.600 ;
        RECT 564.000 510.600 565.800 513.600 ;
        RECT 567.000 510.000 568.800 513.600 ;
        RECT 570.000 510.600 571.800 514.500 ;
        RECT 577.200 513.600 579.300 515.700 ;
        RECT 580.200 513.600 582.300 515.700 ;
        RECT 583.200 513.600 585.300 515.700 ;
        RECT 574.500 510.000 576.300 513.600 ;
        RECT 577.500 510.600 579.300 513.600 ;
        RECT 580.500 510.600 582.300 513.600 ;
        RECT 583.500 510.600 585.300 513.600 ;
        RECT 587.700 510.600 589.500 516.600 ;
        RECT 593.100 510.000 594.900 516.600 ;
        RECT 598.500 510.600 600.300 516.600 ;
        RECT 617.100 516.600 621.900 517.500 ;
        RECT 624.900 516.600 626.100 518.100 ;
        RECT 632.100 516.600 633.300 518.400 ;
        RECT 656.100 516.600 657.300 523.950 ;
        RECT 662.100 522.150 663.900 523.950 ;
        RECT 674.550 523.050 675.450 524.550 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 674.550 521.550 679.050 523.050 ;
        RECT 680.100 522.150 681.900 523.950 ;
        RECT 675.000 520.950 679.050 521.550 ;
        RECT 683.100 519.600 684.300 523.950 ;
        RECT 686.100 522.150 687.900 523.950 ;
        RECT 710.250 522.150 712.050 523.950 ;
        RECT 680.700 518.700 684.300 519.600 ;
        RECT 714.000 519.300 715.050 523.950 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 737.100 524.700 744.000 526.050 ;
        RECT 744.900 525.900 747.300 526.800 ;
        RECT 751.800 526.050 753.600 527.850 ;
        RECT 771.000 526.050 772.200 533.400 ;
        RECT 779.700 531.900 780.900 533.400 ;
        RECT 773.100 530.700 780.900 531.900 ;
        RECT 773.100 530.100 774.900 530.700 ;
        RECT 737.100 523.950 739.200 524.700 ;
        RECT 715.950 522.150 717.750 523.950 ;
        RECT 737.400 522.150 739.200 523.950 ;
        RECT 742.200 521.400 744.000 523.200 ;
        RECT 741.900 519.300 744.000 521.400 ;
        RECT 680.700 516.600 681.900 518.700 ;
        RECT 710.700 518.100 715.050 519.300 ;
        RECT 737.700 518.400 744.000 519.300 ;
        RECT 744.900 520.200 746.100 525.900 ;
        RECT 747.300 523.200 749.100 525.000 ;
        RECT 751.800 523.950 753.900 526.050 ;
        RECT 770.100 523.950 772.200 526.050 ;
        RECT 747.000 521.100 749.100 523.200 ;
        RECT 617.100 510.600 618.900 516.600 ;
        RECT 620.100 510.000 621.900 515.700 ;
        RECT 624.600 510.600 626.400 516.600 ;
        RECT 629.100 510.000 630.900 515.700 ;
        RECT 632.100 510.600 633.900 516.600 ;
        RECT 650.700 510.000 652.500 516.600 ;
        RECT 655.200 510.600 657.000 516.600 ;
        RECT 659.700 510.000 661.500 516.600 ;
        RECT 680.100 510.600 681.900 516.600 ;
        RECT 683.100 515.700 690.900 517.050 ;
        RECT 710.700 516.600 711.600 518.100 ;
        RECT 683.100 510.600 684.900 515.700 ;
        RECT 686.100 510.000 687.900 514.800 ;
        RECT 689.100 510.600 690.900 515.700 ;
        RECT 707.100 511.500 708.900 516.600 ;
        RECT 710.100 512.400 711.900 516.600 ;
        RECT 713.100 516.000 720.900 516.900 ;
        RECT 737.700 516.600 738.900 518.400 ;
        RECT 744.900 518.100 747.900 520.200 ;
        RECT 744.900 516.600 746.100 518.100 ;
        RECT 749.100 517.500 751.200 518.700 ;
        RECT 749.100 516.600 753.900 517.500 ;
        RECT 713.100 511.500 714.900 516.000 ;
        RECT 707.100 510.600 714.900 511.500 ;
        RECT 716.100 510.000 717.900 515.100 ;
        RECT 719.100 510.600 720.900 516.000 ;
        RECT 737.100 510.600 738.900 516.600 ;
        RECT 740.100 510.000 741.900 515.700 ;
        RECT 744.600 510.600 746.400 516.600 ;
        RECT 749.100 510.000 750.900 515.700 ;
        RECT 752.100 510.600 753.900 516.600 ;
        RECT 770.100 516.600 771.000 523.950 ;
        RECT 773.400 519.600 774.300 530.100 ;
        RECT 775.200 526.050 777.000 527.850 ;
        RECT 797.250 526.050 799.050 527.850 ;
        RECT 800.400 526.050 801.300 533.400 ;
        RECT 803.100 526.050 804.900 527.850 ;
        RECT 821.400 526.050 822.300 533.400 ;
        RECT 835.950 529.950 838.050 532.050 ;
        RECT 847.950 531.450 850.050 532.050 ;
        RECT 842.550 530.550 850.050 531.450 ;
        RECT 826.950 526.050 828.750 527.850 ;
        RECT 775.500 523.950 777.600 526.050 ;
        RECT 778.800 523.950 780.900 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 826.950 523.950 829.050 526.050 ;
        RECT 829.950 523.950 832.050 526.050 ;
        RECT 778.800 522.150 780.600 523.950 ;
        RECT 781.950 522.450 784.050 523.050 ;
        RECT 793.950 522.450 796.050 523.050 ;
        RECT 781.950 521.550 796.050 522.450 ;
        RECT 781.950 520.950 784.050 521.550 ;
        RECT 793.950 520.950 796.050 521.550 ;
        RECT 772.200 518.700 774.300 519.600 ;
        RECT 778.950 519.450 781.050 520.050 ;
        RECT 796.950 519.450 799.050 520.050 ;
        RECT 772.200 517.800 777.600 518.700 ;
        RECT 778.950 518.550 799.050 519.450 ;
        RECT 778.950 517.950 781.050 518.550 ;
        RECT 796.950 517.950 799.050 518.550 ;
        RECT 770.100 510.600 771.900 516.600 ;
        RECT 773.100 510.000 774.900 516.000 ;
        RECT 776.700 513.600 777.600 517.800 ;
        RECT 800.400 513.600 801.300 523.950 ;
        RECT 808.950 522.450 811.050 523.050 ;
        RECT 817.950 522.450 820.050 523.050 ;
        RECT 808.950 521.550 820.050 522.450 ;
        RECT 808.950 520.950 811.050 521.550 ;
        RECT 817.950 520.950 820.050 521.550 ;
        RECT 821.400 516.600 822.300 523.950 ;
        RECT 823.950 522.150 825.750 523.950 ;
        RECT 830.100 522.150 831.900 523.950 ;
        RECT 829.950 519.450 832.050 520.050 ;
        RECT 836.550 519.450 837.450 529.950 ;
        RECT 842.550 523.050 843.450 530.550 ;
        RECT 847.950 529.950 850.050 530.550 ;
        RECT 848.250 526.050 850.050 527.850 ;
        RECT 851.400 526.050 852.300 533.400 ;
        RECT 854.100 526.050 855.900 527.850 ;
        RECT 875.100 526.050 876.300 539.400 ;
        RECT 899.400 539.100 900.900 539.400 ;
        RECT 905.100 539.400 906.900 545.400 ;
        RECT 910.950 540.450 913.050 541.050 ;
        RECT 916.950 540.450 919.050 541.050 ;
        RECT 910.950 539.550 919.050 540.450 ;
        RECT 905.100 539.100 906.000 539.400 ;
        RECT 899.400 538.200 906.000 539.100 ;
        RECT 910.950 538.950 913.050 539.550 ;
        RECT 916.950 538.950 919.050 539.550 ;
        RECT 923.100 539.400 924.900 545.400 ;
        RECT 926.100 540.000 927.900 546.000 ;
        RECT 924.000 539.100 924.900 539.400 ;
        RECT 929.100 539.400 930.900 545.400 ;
        RECT 932.100 539.400 933.900 546.000 ;
        RECT 950.700 539.400 952.500 546.000 ;
        RECT 929.100 539.100 930.600 539.400 ;
        RECT 886.950 534.450 889.050 535.050 ;
        RECT 901.950 534.450 904.050 535.050 ;
        RECT 886.950 533.550 904.050 534.450 ;
        RECT 886.950 532.950 889.050 533.550 ;
        RECT 901.950 532.950 904.050 533.550 ;
        RECT 899.100 526.050 900.900 527.850 ;
        RECT 905.100 526.050 906.000 538.200 ;
        RECT 924.000 538.200 930.600 539.100 ;
        RECT 918.000 528.450 922.050 529.050 ;
        RECT 917.550 526.950 922.050 528.450 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 850.950 523.950 853.050 526.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 842.550 521.550 847.050 523.050 ;
        RECT 843.000 520.950 847.050 521.550 ;
        RECT 829.950 518.550 837.450 519.450 ;
        RECT 829.950 517.950 832.050 518.550 ;
        RECT 821.400 515.400 826.500 516.600 ;
        RECT 776.100 510.600 777.900 513.600 ;
        RECT 779.100 510.600 780.900 513.600 ;
        RECT 779.700 510.000 780.900 510.600 ;
        RECT 797.100 510.000 798.900 513.600 ;
        RECT 800.100 510.600 801.900 513.600 ;
        RECT 803.100 510.000 804.900 513.600 ;
        RECT 821.700 510.000 823.500 513.600 ;
        RECT 824.700 510.600 826.500 515.400 ;
        RECT 829.200 510.000 831.000 516.600 ;
        RECT 838.950 513.450 841.050 514.050 ;
        RECT 844.950 513.450 847.050 514.050 ;
        RECT 851.400 513.600 852.300 523.950 ;
        RECT 872.250 522.150 874.050 523.950 ;
        RECT 875.100 518.700 876.300 523.950 ;
        RECT 878.100 522.150 879.900 523.950 ;
        RECT 896.100 522.150 897.900 523.950 ;
        RECT 902.100 522.150 903.900 523.950 ;
        RECT 905.100 520.200 906.000 523.950 ;
        RECT 917.550 523.050 918.450 526.950 ;
        RECT 924.000 526.050 924.900 538.200 ;
        RECT 951.000 536.100 952.800 537.900 ;
        RECT 953.700 534.900 955.500 545.400 ;
        RECT 953.100 533.400 955.500 534.900 ;
        RECT 958.800 533.400 960.600 546.000 ;
        RECT 977.100 539.400 978.900 545.400 ;
        RECT 980.100 540.000 981.900 546.000 ;
        RECT 978.000 539.100 978.900 539.400 ;
        RECT 983.100 539.400 984.900 545.400 ;
        RECT 986.100 539.400 987.900 546.000 ;
        RECT 1004.100 539.400 1005.900 545.400 ;
        RECT 1007.100 540.000 1008.900 546.000 ;
        RECT 983.100 539.100 984.600 539.400 ;
        RECT 978.000 538.200 984.600 539.100 ;
        RECT 1005.000 539.100 1005.900 539.400 ;
        RECT 1010.100 539.400 1011.900 545.400 ;
        RECT 1013.100 539.400 1014.900 546.000 ;
        RECT 1031.100 539.400 1032.900 546.000 ;
        RECT 1034.100 539.400 1035.900 545.400 ;
        RECT 1037.100 539.400 1038.900 546.000 ;
        RECT 1010.100 539.100 1011.600 539.400 ;
        RECT 1005.000 538.200 1011.600 539.100 ;
        RECT 967.950 534.450 970.050 535.050 ;
        RECT 973.950 534.450 976.050 535.050 ;
        RECT 967.950 533.550 976.050 534.450 ;
        RECT 931.950 531.450 934.050 532.050 ;
        RECT 949.950 531.450 952.050 532.200 ;
        RECT 931.950 530.550 952.050 531.450 ;
        RECT 931.950 529.950 934.050 530.550 ;
        RECT 949.950 530.100 952.050 530.550 ;
        RECT 929.100 526.050 930.900 527.850 ;
        RECT 953.100 526.050 954.300 533.400 ;
        RECT 967.950 532.950 970.050 533.550 ;
        RECT 973.950 532.950 976.050 533.550 ;
        RECT 972.000 528.450 976.050 529.050 ;
        RECT 959.100 526.050 960.900 527.850 ;
        RECT 971.550 526.950 976.050 528.450 ;
        RECT 922.950 523.950 925.050 526.050 ;
        RECT 925.950 523.950 928.050 526.050 ;
        RECT 928.950 523.950 931.050 526.050 ;
        RECT 931.950 523.950 934.050 526.050 ;
        RECT 949.950 523.950 952.050 526.050 ;
        RECT 952.950 523.950 955.050 526.050 ;
        RECT 955.950 523.950 958.050 526.050 ;
        RECT 958.950 523.950 961.050 526.050 ;
        RECT 917.550 521.550 922.050 523.050 ;
        RECT 918.000 520.950 922.050 521.550 ;
        RECT 875.100 517.800 879.300 518.700 ;
        RECT 838.950 512.550 847.050 513.450 ;
        RECT 838.950 511.950 841.050 512.550 ;
        RECT 844.950 511.950 847.050 512.550 ;
        RECT 848.100 510.000 849.900 513.600 ;
        RECT 851.100 510.600 852.900 513.600 ;
        RECT 854.100 510.000 855.900 513.600 ;
        RECT 872.400 510.000 874.200 516.600 ;
        RECT 877.500 510.600 879.300 517.800 ;
        RECT 896.100 510.000 897.900 519.600 ;
        RECT 902.700 519.000 906.000 520.200 ;
        RECT 924.000 520.200 924.900 523.950 ;
        RECT 926.100 522.150 927.900 523.950 ;
        RECT 932.100 522.150 933.900 523.950 ;
        RECT 934.950 522.450 937.050 523.050 ;
        RECT 946.950 522.450 949.050 523.050 ;
        RECT 934.950 521.550 949.050 522.450 ;
        RECT 950.100 522.150 951.900 523.950 ;
        RECT 934.950 520.950 937.050 521.550 ;
        RECT 946.950 520.950 949.050 521.550 ;
        RECT 924.000 519.000 927.300 520.200 ;
        RECT 953.100 519.600 954.300 523.950 ;
        RECT 956.100 522.150 957.900 523.950 ;
        RECT 971.550 523.050 972.450 526.950 ;
        RECT 978.000 526.050 978.900 538.200 ;
        RECT 985.950 537.450 988.050 538.050 ;
        RECT 991.950 537.450 994.050 538.050 ;
        RECT 985.950 536.550 994.050 537.450 ;
        RECT 985.950 535.950 988.050 536.550 ;
        RECT 991.950 535.950 994.050 536.550 ;
        RECT 979.950 531.450 982.050 532.200 ;
        RECT 985.950 531.450 988.050 532.050 ;
        RECT 997.950 531.450 1000.050 532.050 ;
        RECT 979.950 530.550 1000.050 531.450 ;
        RECT 979.950 530.100 982.050 530.550 ;
        RECT 985.950 529.950 988.050 530.550 ;
        RECT 997.950 529.950 1000.050 530.550 ;
        RECT 983.100 526.050 984.900 527.850 ;
        RECT 1005.000 526.050 1005.900 538.200 ;
        RECT 1006.950 534.450 1009.050 535.050 ;
        RECT 1030.950 534.450 1033.050 535.050 ;
        RECT 1006.950 533.550 1033.050 534.450 ;
        RECT 1006.950 532.950 1009.050 533.550 ;
        RECT 1030.950 532.950 1033.050 533.550 ;
        RECT 1006.950 531.450 1009.050 531.900 ;
        RECT 1031.550 531.450 1032.450 532.950 ;
        RECT 1006.950 530.550 1017.450 531.450 ;
        RECT 1006.950 529.800 1009.050 530.550 ;
        RECT 1016.550 528.450 1017.450 530.550 ;
        RECT 1025.550 530.550 1032.450 531.450 ;
        RECT 1010.100 526.050 1011.900 527.850 ;
        RECT 1016.550 527.550 1020.450 528.450 ;
        RECT 976.950 523.950 979.050 526.050 ;
        RECT 979.950 523.950 982.050 526.050 ;
        RECT 982.950 523.950 985.050 526.050 ;
        RECT 985.950 523.950 988.050 526.050 ;
        RECT 1003.950 523.950 1006.050 526.050 ;
        RECT 1006.950 523.950 1009.050 526.050 ;
        RECT 1009.950 523.950 1012.050 526.050 ;
        RECT 1012.950 523.950 1015.050 526.050 ;
        RECT 971.550 521.550 976.050 523.050 ;
        RECT 972.000 520.950 976.050 521.550 ;
        RECT 902.700 510.600 904.500 519.000 ;
        RECT 925.500 510.600 927.300 519.000 ;
        RECT 932.100 510.000 933.900 519.600 ;
        RECT 950.700 518.700 954.300 519.600 ;
        RECT 978.000 520.200 978.900 523.950 ;
        RECT 980.100 522.150 981.900 523.950 ;
        RECT 986.100 522.150 987.900 523.950 ;
        RECT 1005.000 520.200 1005.900 523.950 ;
        RECT 1007.100 522.150 1008.900 523.950 ;
        RECT 1013.100 522.150 1014.900 523.950 ;
        RECT 1019.550 523.050 1020.450 527.550 ;
        RECT 1015.950 521.550 1020.450 523.050 ;
        RECT 1025.550 523.050 1026.450 530.550 ;
        RECT 1034.700 526.050 1035.900 539.400 ;
        RECT 1030.950 523.950 1033.050 526.050 ;
        RECT 1033.950 523.950 1036.050 526.050 ;
        RECT 1036.950 523.950 1039.050 526.050 ;
        RECT 1025.550 521.550 1030.050 523.050 ;
        RECT 1031.100 522.150 1032.900 523.950 ;
        RECT 1015.950 520.950 1020.000 521.550 ;
        RECT 1026.000 520.950 1030.050 521.550 ;
        RECT 978.000 519.000 981.300 520.200 ;
        RECT 950.700 516.600 951.900 518.700 ;
        RECT 950.100 510.600 951.900 516.600 ;
        RECT 953.100 515.700 960.900 517.050 ;
        RECT 953.100 510.600 954.900 515.700 ;
        RECT 956.100 510.000 957.900 514.800 ;
        RECT 959.100 510.600 960.900 515.700 ;
        RECT 979.500 510.600 981.300 519.000 ;
        RECT 986.100 510.000 987.900 519.600 ;
        RECT 1005.000 519.000 1008.300 520.200 ;
        RECT 1006.500 510.600 1008.300 519.000 ;
        RECT 1013.100 510.000 1014.900 519.600 ;
        RECT 1034.700 518.700 1035.900 523.950 ;
        RECT 1036.950 522.150 1038.750 523.950 ;
        RECT 1031.700 517.800 1035.900 518.700 ;
        RECT 1031.700 510.600 1033.500 517.800 ;
        RECT 1036.800 510.000 1038.600 516.600 ;
        RECT 17.100 503.400 18.900 507.000 ;
        RECT 20.100 503.400 21.900 506.400 ;
        RECT 38.100 503.400 39.900 506.400 ;
        RECT 41.100 503.400 42.900 507.000 ;
        RECT 4.950 495.450 7.050 496.050 ;
        RECT 13.950 495.450 16.050 496.050 ;
        RECT 4.950 494.550 16.050 495.450 ;
        RECT 4.950 493.950 7.050 494.550 ;
        RECT 13.950 493.950 16.050 494.550 ;
        RECT 20.100 493.050 21.300 503.400 ;
        RECT 38.700 493.050 39.900 503.400 ;
        RECT 59.400 500.400 61.200 507.000 ;
        RECT 64.500 499.200 66.300 506.400 ;
        RECT 62.100 498.300 66.300 499.200 ;
        RECT 59.250 493.050 61.050 494.850 ;
        RECT 62.100 493.050 63.300 498.300 ;
        RECT 85.500 498.000 87.300 506.400 ;
        RECT 84.000 496.800 87.300 498.000 ;
        RECT 92.100 497.400 93.900 507.000 ;
        RECT 112.500 498.000 114.300 506.400 ;
        RECT 111.000 496.800 114.300 498.000 ;
        RECT 119.100 497.400 120.900 507.000 ;
        RECT 137.400 500.400 139.200 507.000 ;
        RECT 142.500 499.200 144.300 506.400 ;
        RECT 166.200 503.400 168.900 506.400 ;
        RECT 170.100 503.400 171.900 507.000 ;
        RECT 173.100 503.400 174.900 506.400 ;
        RECT 176.100 503.400 178.200 507.000 ;
        RECT 197.100 503.400 198.900 507.000 ;
        RECT 200.100 503.400 201.900 506.400 ;
        RECT 203.100 503.400 204.900 507.000 ;
        RECT 166.200 502.500 167.100 503.400 ;
        RECT 173.400 502.500 174.300 503.400 ;
        RECT 140.100 498.300 144.300 499.200 ;
        RECT 161.700 501.600 174.300 502.500 ;
        RECT 65.100 493.050 66.900 494.850 ;
        RECT 84.000 493.050 84.900 496.800 ;
        RECT 86.100 493.050 87.900 494.850 ;
        RECT 92.100 493.050 93.900 494.850 ;
        RECT 111.000 493.050 111.900 496.800 ;
        RECT 113.100 493.050 114.900 494.850 ;
        RECT 119.100 493.050 120.900 494.850 ;
        RECT 137.250 493.050 139.050 494.850 ;
        RECT 140.100 493.050 141.300 498.300 ;
        RECT 143.100 493.050 144.900 494.850 ;
        RECT 161.700 493.050 162.900 501.600 ;
        RECT 187.950 501.450 190.050 502.050 ;
        RECT 193.950 501.450 196.050 502.050 ;
        RECT 187.950 500.550 196.050 501.450 ;
        RECT 187.950 499.950 190.050 500.550 ;
        RECT 193.950 499.950 196.050 500.550 ;
        RECT 166.950 498.450 169.050 499.050 ;
        RECT 172.950 498.450 175.050 499.050 ;
        RECT 196.950 498.450 199.050 499.200 ;
        RECT 166.950 497.550 199.050 498.450 ;
        RECT 166.950 496.950 169.050 497.550 ;
        RECT 172.950 496.950 175.050 497.550 ;
        RECT 196.950 497.100 199.050 497.550 ;
        RECT 178.950 495.450 181.050 496.050 ;
        RECT 193.950 495.450 196.050 496.050 ;
        RECT 170.250 493.050 172.050 494.850 ;
        RECT 178.950 494.550 196.050 495.450 ;
        RECT 178.950 493.950 181.050 494.550 ;
        RECT 193.950 493.950 196.050 494.550 ;
        RECT 200.400 493.050 201.300 503.400 ;
        RECT 221.100 500.400 222.900 506.400 ;
        RECT 224.100 500.400 225.900 507.000 ;
        RECT 242.400 500.400 244.200 507.000 ;
        RECT 221.700 493.050 222.900 500.400 ;
        RECT 247.500 499.200 249.300 506.400 ;
        RECT 266.100 503.400 267.900 507.000 ;
        RECT 269.100 503.400 270.900 506.400 ;
        RECT 272.100 503.400 273.900 507.000 ;
        RECT 253.950 501.450 256.050 502.050 ;
        RECT 265.950 501.450 268.050 501.900 ;
        RECT 253.950 500.550 268.050 501.450 ;
        RECT 253.950 499.950 256.050 500.550 ;
        RECT 265.950 499.800 268.050 500.550 ;
        RECT 245.100 498.300 249.300 499.200 ;
        RECT 224.100 493.050 225.900 494.850 ;
        RECT 242.250 493.050 244.050 494.850 ;
        RECT 245.100 493.050 246.300 498.300 ;
        RECT 250.950 495.450 253.050 496.050 ;
        RECT 259.950 495.450 262.050 496.050 ;
        RECT 248.100 493.050 249.900 494.850 ;
        RECT 250.950 494.550 262.050 495.450 ;
        RECT 250.950 493.950 253.050 494.550 ;
        RECT 259.950 493.950 262.050 494.550 ;
        RECT 269.400 493.050 270.300 503.400 ;
        RECT 292.500 498.000 294.300 506.400 ;
        RECT 291.000 496.800 294.300 498.000 ;
        RECT 299.100 497.400 300.900 507.000 ;
        RECT 317.100 500.400 318.900 507.000 ;
        RECT 320.100 500.400 321.900 506.400 ;
        RECT 291.000 493.050 291.900 496.800 ;
        RECT 293.100 493.050 294.900 494.850 ;
        RECT 299.100 493.050 300.900 494.850 ;
        RECT 317.100 493.050 318.900 494.850 ;
        RECT 320.100 493.050 321.300 500.400 ;
        RECT 338.100 497.400 339.900 507.000 ;
        RECT 365.100 506.400 366.300 507.000 ;
        RECT 344.700 498.000 346.500 506.400 ;
        RECT 365.100 503.400 366.900 506.400 ;
        RECT 368.100 503.400 369.900 506.400 ;
        RECT 368.400 499.200 369.300 503.400 ;
        RECT 371.100 501.000 372.900 507.000 ;
        RECT 374.100 500.400 375.900 506.400 ;
        RECT 392.100 503.400 393.900 507.000 ;
        RECT 395.100 503.400 396.900 506.400 ;
        RECT 398.100 503.400 399.900 507.000 ;
        RECT 416.100 503.400 417.900 507.000 ;
        RECT 419.100 503.400 420.900 506.400 ;
        RECT 422.100 503.400 423.900 507.000 ;
        RECT 368.400 498.300 373.800 499.200 ;
        RECT 344.700 496.800 348.000 498.000 ;
        RECT 322.950 495.450 325.050 496.050 ;
        RECT 334.950 495.450 337.050 496.050 ;
        RECT 322.950 494.550 337.050 495.450 ;
        RECT 322.950 493.950 325.050 494.550 ;
        RECT 334.950 493.950 337.050 494.550 ;
        RECT 338.100 493.050 339.900 494.850 ;
        RECT 344.100 493.050 345.900 494.850 ;
        RECT 347.100 493.050 348.000 496.800 ;
        RECT 371.700 497.400 373.800 498.300 ;
        RECT 365.400 493.050 367.200 494.850 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 64.950 490.950 67.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 88.950 490.950 91.050 493.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 115.950 490.950 118.050 493.050 ;
        RECT 118.950 490.950 121.050 493.050 ;
        RECT 136.950 490.950 139.050 493.050 ;
        RECT 139.950 490.950 142.050 493.050 ;
        RECT 142.950 490.950 145.050 493.050 ;
        RECT 161.400 490.950 163.500 493.050 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 176.100 490.950 178.200 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 268.950 490.950 271.050 493.050 ;
        RECT 271.950 490.950 274.050 493.050 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 295.950 490.950 298.050 493.050 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 365.100 490.950 367.200 493.050 ;
        RECT 368.400 490.950 370.500 493.050 ;
        RECT 17.100 489.150 18.900 490.950 ;
        RECT 20.100 477.600 21.300 490.950 ;
        RECT 38.700 477.600 39.900 490.950 ;
        RECT 41.100 489.150 42.900 490.950 ;
        RECT 62.100 477.600 63.300 490.950 ;
        RECT 84.000 478.800 84.900 490.950 ;
        RECT 89.100 489.150 90.900 490.950 ;
        RECT 111.000 478.800 111.900 490.950 ;
        RECT 116.100 489.150 117.900 490.950 ;
        RECT 112.950 486.450 115.050 487.050 ;
        RECT 121.950 486.450 124.050 487.050 ;
        RECT 112.950 485.550 124.050 486.450 ;
        RECT 112.950 484.950 115.050 485.550 ;
        RECT 121.950 484.950 124.050 485.550 ;
        RECT 84.000 477.900 90.600 478.800 ;
        RECT 84.000 477.600 84.900 477.900 ;
        RECT 17.100 471.000 18.900 477.600 ;
        RECT 20.100 471.600 21.900 477.600 ;
        RECT 38.100 471.600 39.900 477.600 ;
        RECT 41.100 471.000 42.900 477.600 ;
        RECT 59.100 471.000 60.900 477.600 ;
        RECT 62.100 471.600 63.900 477.600 ;
        RECT 65.100 471.000 66.900 477.600 ;
        RECT 83.100 471.600 84.900 477.600 ;
        RECT 89.100 477.600 90.600 477.900 ;
        RECT 111.000 477.900 117.600 478.800 ;
        RECT 111.000 477.600 111.900 477.900 ;
        RECT 86.100 471.000 87.900 477.000 ;
        RECT 89.100 471.600 90.900 477.600 ;
        RECT 92.100 471.000 93.900 477.600 ;
        RECT 110.100 471.600 111.900 477.600 ;
        RECT 116.100 477.600 117.600 477.900 ;
        RECT 140.100 477.600 141.300 490.950 ;
        RECT 113.100 471.000 114.900 477.000 ;
        RECT 116.100 471.600 117.900 477.600 ;
        RECT 119.100 471.000 120.900 477.600 ;
        RECT 137.100 471.000 138.900 477.600 ;
        RECT 140.100 471.600 141.900 477.600 ;
        RECT 143.100 471.000 144.900 477.600 ;
        RECT 158.100 472.500 159.900 481.800 ;
        RECT 161.700 481.200 162.900 490.950 ;
        RECT 166.950 489.150 168.750 490.950 ;
        RECT 176.100 489.150 177.900 490.950 ;
        RECT 197.250 489.150 199.050 490.950 ;
        RECT 169.950 486.450 172.050 487.050 ;
        RECT 184.950 486.450 187.050 487.050 ;
        RECT 169.950 485.550 187.050 486.450 ;
        RECT 169.950 484.950 172.050 485.550 ;
        RECT 184.950 484.950 187.050 485.550 ;
        RECT 200.400 483.600 201.300 490.950 ;
        RECT 203.100 489.150 204.900 490.950 ;
        RECT 221.700 483.600 222.900 490.950 ;
        RECT 223.950 486.450 226.050 487.050 ;
        RECT 229.950 486.450 232.050 487.050 ;
        RECT 223.950 485.550 232.050 486.450 ;
        RECT 223.950 484.950 226.050 485.550 ;
        RECT 229.950 484.950 232.050 485.550 ;
        RECT 161.100 473.400 162.900 481.200 ;
        RECT 164.100 481.200 171.900 482.100 ;
        RECT 164.100 472.500 165.900 481.200 ;
        RECT 158.100 471.600 165.900 472.500 ;
        RECT 167.100 472.500 168.900 480.300 ;
        RECT 170.100 473.400 171.900 481.200 ;
        RECT 173.100 481.500 180.900 482.400 ;
        RECT 173.100 472.500 174.900 481.500 ;
        RECT 167.100 471.600 174.900 472.500 ;
        RECT 176.100 471.000 177.900 480.600 ;
        RECT 179.100 471.600 180.900 481.500 ;
        RECT 197.100 471.000 198.900 483.600 ;
        RECT 200.400 482.400 204.000 483.600 ;
        RECT 202.200 471.600 204.000 482.400 ;
        RECT 221.100 471.600 222.900 483.600 ;
        RECT 224.100 471.000 225.900 483.600 ;
        RECT 245.100 477.600 246.300 490.950 ;
        RECT 266.250 489.150 268.050 490.950 ;
        RECT 269.400 483.600 270.300 490.950 ;
        RECT 272.100 489.150 273.900 490.950 ;
        RECT 242.100 471.000 243.900 477.600 ;
        RECT 245.100 471.600 246.900 477.600 ;
        RECT 248.100 471.000 249.900 477.600 ;
        RECT 266.100 471.000 267.900 483.600 ;
        RECT 269.400 482.400 273.000 483.600 ;
        RECT 271.200 471.600 273.000 482.400 ;
        RECT 291.000 478.800 291.900 490.950 ;
        RECT 296.100 489.150 297.900 490.950 ;
        RECT 320.100 483.600 321.300 490.950 ;
        RECT 341.100 489.150 342.900 490.950 ;
        RECT 291.000 477.900 297.600 478.800 ;
        RECT 291.000 477.600 291.900 477.900 ;
        RECT 290.100 471.600 291.900 477.600 ;
        RECT 296.100 477.600 297.600 477.900 ;
        RECT 293.100 471.000 294.900 477.000 ;
        RECT 296.100 471.600 297.900 477.600 ;
        RECT 299.100 471.000 300.900 477.600 ;
        RECT 317.100 471.000 318.900 483.600 ;
        RECT 320.100 471.600 321.900 483.600 ;
        RECT 347.100 478.800 348.000 490.950 ;
        RECT 369.000 489.150 370.800 490.950 ;
        RECT 371.700 486.900 372.600 497.400 ;
        RECT 375.000 493.050 375.900 500.400 ;
        RECT 395.700 493.050 396.600 503.400 ;
        RECT 419.700 493.050 420.600 503.400 ;
        RECT 440.100 500.400 441.900 506.400 ;
        RECT 440.700 498.300 441.900 500.400 ;
        RECT 443.100 501.300 444.900 506.400 ;
        RECT 446.100 502.200 447.900 507.000 ;
        RECT 449.100 501.300 450.900 506.400 ;
        RECT 467.700 503.400 469.500 507.000 ;
        RECT 470.700 501.600 472.500 506.400 ;
        RECT 443.100 499.950 450.900 501.300 ;
        RECT 467.400 500.400 472.500 501.600 ;
        RECT 475.200 500.400 477.000 507.000 ;
        RECT 494.100 500.400 495.900 506.400 ;
        RECT 440.700 497.400 444.300 498.300 ;
        RECT 440.100 493.050 441.900 494.850 ;
        RECT 443.100 493.050 444.300 497.400 ;
        RECT 446.100 493.050 447.900 494.850 ;
        RECT 467.400 493.050 468.300 500.400 ;
        RECT 469.950 498.450 472.050 499.050 ;
        RECT 487.950 498.450 490.050 498.900 ;
        RECT 469.950 497.550 490.050 498.450 ;
        RECT 469.950 496.950 472.050 497.550 ;
        RECT 487.950 496.800 490.050 497.550 ;
        RECT 494.700 498.300 495.900 500.400 ;
        RECT 497.100 501.300 498.900 506.400 ;
        RECT 500.100 502.200 501.900 507.000 ;
        RECT 503.100 501.300 504.900 506.400 ;
        RECT 497.100 499.950 504.900 501.300 ;
        RECT 521.100 500.400 522.900 506.400 ;
        RECT 524.100 501.300 525.900 507.000 ;
        RECT 528.600 500.400 530.400 506.400 ;
        RECT 533.100 501.300 534.900 507.000 ;
        RECT 536.100 500.400 537.900 506.400 ;
        RECT 539.700 503.400 541.500 507.000 ;
        RECT 542.700 503.400 544.500 506.400 ;
        RECT 521.100 499.500 525.900 500.400 ;
        RECT 523.800 498.300 525.900 499.500 ;
        RECT 528.900 498.900 530.100 500.400 ;
        RECT 494.700 497.400 498.300 498.300 ;
        RECT 469.950 493.050 471.750 494.850 ;
        RECT 476.100 493.050 477.900 494.850 ;
        RECT 494.100 493.050 495.900 494.850 ;
        RECT 497.100 493.050 498.300 497.400 ;
        RECT 527.100 496.800 530.100 498.900 ;
        RECT 536.100 498.600 537.300 500.400 ;
        RECT 500.100 493.050 501.900 494.850 ;
        RECT 525.900 493.800 528.000 495.900 ;
        RECT 373.800 490.950 375.900 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 466.950 490.950 469.050 493.050 ;
        RECT 469.950 490.950 472.050 493.050 ;
        RECT 472.950 490.950 475.050 493.050 ;
        RECT 475.950 490.950 478.050 493.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 499.950 490.950 502.050 493.050 ;
        RECT 502.950 490.950 505.050 493.050 ;
        RECT 521.100 490.950 523.200 493.050 ;
        RECT 525.900 492.000 527.700 493.800 ;
        RECT 528.900 491.100 530.100 496.800 ;
        RECT 531.000 497.700 537.300 498.600 ;
        RECT 531.000 495.600 533.100 497.700 ;
        RECT 531.000 493.800 532.800 495.600 ;
        RECT 535.800 493.050 537.600 494.850 ;
        RECT 535.800 492.300 537.900 493.050 ;
        RECT 371.100 486.300 372.900 486.900 ;
        RECT 341.400 477.900 348.000 478.800 ;
        RECT 341.400 477.600 342.900 477.900 ;
        RECT 338.100 471.000 339.900 477.600 ;
        RECT 341.100 471.600 342.900 477.600 ;
        RECT 347.100 477.600 348.000 477.900 ;
        RECT 365.100 485.100 372.900 486.300 ;
        RECT 365.100 483.600 366.300 485.100 ;
        RECT 373.800 483.600 375.000 490.950 ;
        RECT 392.100 489.150 393.900 490.950 ;
        RECT 395.700 483.600 396.600 490.950 ;
        RECT 397.950 489.150 399.750 490.950 ;
        RECT 416.100 489.150 417.900 490.950 ;
        RECT 419.700 483.600 420.600 490.950 ;
        RECT 421.950 489.150 423.750 490.950 ;
        RECT 443.100 483.600 444.300 490.950 ;
        RECT 449.100 489.150 450.900 490.950 ;
        RECT 467.400 483.600 468.300 490.950 ;
        RECT 472.950 489.150 474.750 490.950 ;
        RECT 497.100 483.600 498.300 490.950 ;
        RECT 503.100 489.150 504.900 490.950 ;
        RECT 521.400 489.150 523.200 490.950 ;
        RECT 527.700 490.200 530.100 491.100 ;
        RECT 531.000 490.950 537.900 492.300 ;
        RECT 531.000 490.500 532.800 490.950 ;
        RECT 527.700 490.050 529.200 490.200 ;
        RECT 543.000 490.050 544.500 503.400 ;
        RECT 527.100 487.950 529.200 490.050 ;
        RECT 502.950 486.450 505.050 487.050 ;
        RECT 517.950 486.450 520.050 487.050 ;
        RECT 502.950 485.550 520.050 486.450 ;
        RECT 502.950 484.950 505.050 485.550 ;
        RECT 517.950 484.950 520.050 485.550 ;
        RECT 528.300 486.000 529.200 487.950 ;
        RECT 530.100 487.500 534.000 489.300 ;
        RECT 542.100 487.950 544.500 490.050 ;
        RECT 530.100 487.200 532.200 487.500 ;
        RECT 528.300 484.950 529.800 486.000 ;
        RECT 523.800 483.600 525.900 484.500 ;
        RECT 344.100 471.000 345.900 477.000 ;
        RECT 347.100 471.600 348.900 477.600 ;
        RECT 365.100 471.600 366.900 483.600 ;
        RECT 369.600 471.000 371.400 483.600 ;
        RECT 372.600 482.100 375.000 483.600 ;
        RECT 393.000 482.400 396.600 483.600 ;
        RECT 372.600 471.600 374.400 482.100 ;
        RECT 393.000 471.600 394.800 482.400 ;
        RECT 398.100 471.000 399.900 483.600 ;
        RECT 417.000 482.400 420.600 483.600 ;
        RECT 417.000 471.600 418.800 482.400 ;
        RECT 422.100 471.000 423.900 483.600 ;
        RECT 443.100 482.100 445.500 483.600 ;
        RECT 441.000 479.100 442.800 480.900 ;
        RECT 440.700 471.000 442.500 477.600 ;
        RECT 443.700 471.600 445.500 482.100 ;
        RECT 448.800 471.000 450.600 483.600 ;
        RECT 467.100 471.600 468.900 483.600 ;
        RECT 470.100 482.700 477.900 483.600 ;
        RECT 470.100 471.600 471.900 482.700 ;
        RECT 473.100 471.000 474.900 481.800 ;
        RECT 476.100 471.600 477.900 482.700 ;
        RECT 497.100 482.100 499.500 483.600 ;
        RECT 495.000 479.100 496.800 480.900 ;
        RECT 494.700 471.000 496.500 477.600 ;
        RECT 497.700 471.600 499.500 482.100 ;
        RECT 502.800 471.000 504.600 483.600 ;
        RECT 521.100 482.400 525.900 483.600 ;
        RECT 528.600 483.600 529.800 484.950 ;
        RECT 533.400 483.600 535.500 485.700 ;
        RECT 521.100 471.600 522.900 482.400 ;
        RECT 524.100 471.000 525.900 481.500 ;
        RECT 528.600 471.600 530.400 483.600 ;
        RECT 533.400 482.700 537.900 483.600 ;
        RECT 533.100 471.000 534.900 481.500 ;
        RECT 536.100 471.600 537.900 482.700 ;
        RECT 543.000 477.600 544.500 487.950 ;
        RECT 546.300 500.400 548.100 506.400 ;
        RECT 551.700 500.400 553.500 507.000 ;
        RECT 556.800 501.600 558.600 506.400 ;
        RECT 561.000 503.400 562.800 506.400 ;
        RECT 564.000 503.400 565.800 506.400 ;
        RECT 567.000 503.400 568.800 506.400 ;
        RECT 570.000 503.400 571.800 506.400 ;
        RECT 573.000 503.400 574.800 507.000 ;
        RECT 554.400 500.400 558.600 501.600 ;
        RECT 560.700 501.300 562.800 503.400 ;
        RECT 563.700 501.300 565.800 503.400 ;
        RECT 566.700 501.300 568.800 503.400 ;
        RECT 569.700 501.300 571.800 503.400 ;
        RECT 576.000 502.500 577.800 506.400 ;
        RECT 580.500 503.400 582.300 507.000 ;
        RECT 583.500 503.400 585.300 506.400 ;
        RECT 586.500 503.400 588.300 506.400 ;
        RECT 589.500 503.400 591.300 506.400 ;
        RECT 575.100 500.400 577.800 502.500 ;
        RECT 579.600 501.600 581.400 502.500 ;
        RECT 579.600 500.400 582.300 501.600 ;
        RECT 583.200 501.300 585.300 503.400 ;
        RECT 586.200 501.300 588.300 503.400 ;
        RECT 589.200 501.300 591.300 503.400 ;
        RECT 593.700 500.400 595.500 506.400 ;
        RECT 599.100 500.400 600.900 507.000 ;
        RECT 604.500 500.400 606.300 506.400 ;
        RECT 623.100 500.400 624.900 506.400 ;
        RECT 626.100 501.300 627.900 507.000 ;
        RECT 630.600 500.400 632.400 506.400 ;
        RECT 635.100 501.300 636.900 507.000 ;
        RECT 638.100 500.400 639.900 506.400 ;
        RECT 546.300 483.600 547.200 500.400 ;
        RECT 554.400 497.100 555.900 500.400 ;
        RECT 560.100 498.600 566.700 500.400 ;
        RECT 581.400 499.800 582.300 500.400 ;
        RECT 584.400 499.800 586.200 500.400 ;
        RECT 581.400 498.600 588.600 499.800 ;
        RECT 548.100 495.300 555.900 497.100 ;
        RECT 572.100 496.500 573.900 498.300 ;
        RECT 571.800 495.900 573.900 496.500 ;
        RECT 556.800 494.400 573.900 495.900 ;
        RECT 578.100 495.900 580.200 496.050 ;
        RECT 581.400 495.900 583.200 496.800 ;
        RECT 578.100 495.000 583.200 495.900 ;
        RECT 587.700 495.600 588.600 498.600 ;
        RECT 593.700 499.500 595.200 500.400 ;
        RECT 593.700 498.300 602.100 499.500 ;
        RECT 600.300 497.700 602.100 498.300 ;
        RECT 589.500 496.800 591.600 497.700 ;
        RECT 605.100 496.800 606.300 500.400 ;
        RECT 607.950 498.450 610.050 499.050 ;
        RECT 613.950 498.450 616.050 499.050 ;
        RECT 607.950 497.550 616.050 498.450 ;
        RECT 623.700 498.600 624.900 500.400 ;
        RECT 630.900 498.900 632.100 500.400 ;
        RECT 635.100 499.500 639.900 500.400 ;
        RECT 641.700 500.400 643.500 506.400 ;
        RECT 647.100 500.400 648.900 507.000 ;
        RECT 652.500 500.400 654.300 506.400 ;
        RECT 656.700 503.400 658.500 506.400 ;
        RECT 659.700 503.400 661.500 506.400 ;
        RECT 662.700 503.400 664.500 506.400 ;
        RECT 665.700 503.400 667.500 507.000 ;
        RECT 656.700 501.300 658.800 503.400 ;
        RECT 659.700 501.300 661.800 503.400 ;
        RECT 662.700 501.300 664.800 503.400 ;
        RECT 670.200 502.500 672.000 506.400 ;
        RECT 673.200 503.400 675.000 507.000 ;
        RECT 676.200 503.400 678.000 506.400 ;
        RECT 679.200 503.400 681.000 506.400 ;
        RECT 682.200 503.400 684.000 506.400 ;
        RECT 685.200 503.400 687.000 506.400 ;
        RECT 666.600 501.600 668.400 502.500 ;
        RECT 665.700 500.400 668.400 501.600 ;
        RECT 670.200 500.400 672.900 502.500 ;
        RECT 676.200 501.300 678.300 503.400 ;
        RECT 679.200 501.300 681.300 503.400 ;
        RECT 682.200 501.300 684.300 503.400 ;
        RECT 685.200 501.300 687.300 503.400 ;
        RECT 689.400 501.600 691.200 506.400 ;
        RECT 689.400 500.400 693.600 501.600 ;
        RECT 694.500 500.400 696.300 507.000 ;
        RECT 699.900 500.400 701.700 506.400 ;
        RECT 623.700 497.700 630.000 498.600 ;
        RECT 607.950 496.950 610.050 497.550 ;
        RECT 613.950 496.950 616.050 497.550 ;
        RECT 589.500 495.600 606.300 496.800 ;
        RECT 627.900 495.600 630.000 497.700 ;
        RECT 551.700 492.900 558.300 494.400 ;
        RECT 578.100 493.950 580.200 495.000 ;
        RECT 586.800 493.800 588.600 495.600 ;
        RECT 551.700 490.050 553.200 492.900 ;
        RECT 559.500 491.700 603.900 492.900 ;
        RECT 559.500 490.200 560.400 491.700 ;
        RECT 551.100 487.950 553.200 490.050 ;
        RECT 555.300 488.400 560.400 490.200 ;
        RECT 563.100 489.900 576.600 490.800 ;
        RECT 583.800 489.900 585.600 490.500 ;
        RECT 602.100 490.050 603.900 491.700 ;
        RECT 563.100 488.700 564.000 489.900 ;
        RECT 563.100 486.900 564.900 488.700 ;
        RECT 569.100 487.200 573.000 489.000 ;
        RECT 574.500 488.700 585.600 489.900 ;
        RECT 596.100 489.750 598.200 490.050 ;
        RECT 574.500 487.800 576.600 488.700 ;
        RECT 594.300 487.950 598.200 489.750 ;
        RECT 602.100 487.950 604.200 490.050 ;
        RECT 594.300 487.200 596.100 487.950 ;
        RECT 569.100 486.900 571.200 487.200 ;
        RECT 582.600 486.300 596.100 487.200 ;
        RECT 548.100 485.700 549.900 486.300 ;
        RECT 582.600 485.700 583.800 486.300 ;
        RECT 548.100 484.500 583.800 485.700 ;
        RECT 586.500 484.500 588.600 484.800 ;
        RECT 546.300 482.700 562.800 483.600 ;
        RECT 546.300 479.400 547.200 482.700 ;
        RECT 551.100 480.600 556.800 481.800 ;
        RECT 560.700 481.500 562.800 482.700 ;
        RECT 566.100 482.400 583.800 483.600 ;
        RECT 586.500 483.300 598.500 484.500 ;
        RECT 586.500 482.700 588.600 483.300 ;
        RECT 596.700 482.700 598.500 483.300 ;
        RECT 566.100 481.500 568.200 482.400 ;
        RECT 582.600 481.800 583.800 482.400 ;
        RECT 600.000 481.800 601.800 482.100 ;
        RECT 551.100 480.000 552.900 480.600 ;
        RECT 546.300 478.500 550.200 479.400 ;
        RECT 549.000 477.600 550.200 478.500 ;
        RECT 555.600 477.600 556.800 480.600 ;
        RECT 557.700 479.700 559.500 480.300 ;
        RECT 557.700 478.500 565.800 479.700 ;
        RECT 563.700 477.600 565.800 478.500 ;
        RECT 569.100 477.600 571.800 481.500 ;
        RECT 574.500 479.100 577.800 481.200 ;
        RECT 582.600 480.600 601.800 481.800 ;
        RECT 539.700 471.000 541.500 477.600 ;
        RECT 542.700 471.600 544.500 477.600 ;
        RECT 546.000 471.000 547.800 477.600 ;
        RECT 549.000 471.600 550.800 477.600 ;
        RECT 552.000 471.000 553.800 477.600 ;
        RECT 555.000 471.600 556.800 477.600 ;
        RECT 558.000 471.000 559.800 477.600 ;
        RECT 560.700 474.600 562.800 476.700 ;
        RECT 563.700 474.600 565.800 476.700 ;
        RECT 566.700 474.600 568.800 476.700 ;
        RECT 561.000 471.600 562.800 474.600 ;
        RECT 564.000 471.600 565.800 474.600 ;
        RECT 567.000 471.600 568.800 474.600 ;
        RECT 570.000 471.600 571.800 477.600 ;
        RECT 573.000 471.000 574.800 477.600 ;
        RECT 576.000 471.600 577.800 479.100 ;
        RECT 583.200 477.600 585.300 479.700 ;
        RECT 579.900 471.000 581.700 477.600 ;
        RECT 582.900 471.600 584.700 477.600 ;
        RECT 585.600 474.600 587.700 476.700 ;
        RECT 588.600 474.600 590.700 476.700 ;
        RECT 585.900 471.600 587.700 474.600 ;
        RECT 588.900 471.600 590.700 474.600 ;
        RECT 592.500 471.000 594.300 477.600 ;
        RECT 595.500 471.600 597.300 480.600 ;
        RECT 600.000 480.300 601.800 480.600 ;
        RECT 605.100 479.400 606.300 495.600 ;
        RECT 623.400 493.050 625.200 494.850 ;
        RECT 628.200 493.800 630.000 495.600 ;
        RECT 630.900 496.800 633.900 498.900 ;
        RECT 635.100 498.300 637.200 499.500 ;
        RECT 641.700 496.800 642.900 500.400 ;
        RECT 652.800 499.500 654.300 500.400 ;
        RECT 661.800 499.800 663.600 500.400 ;
        RECT 665.700 499.800 666.600 500.400 ;
        RECT 645.900 498.300 654.300 499.500 ;
        RECT 659.400 498.600 666.600 499.800 ;
        RECT 681.300 498.600 687.900 500.400 ;
        RECT 645.900 497.700 647.700 498.300 ;
        RECT 656.400 496.800 658.500 497.700 ;
        RECT 623.100 492.300 625.200 493.050 ;
        RECT 623.100 490.950 630.000 492.300 ;
        RECT 628.200 490.500 630.000 490.950 ;
        RECT 630.900 491.100 632.100 496.800 ;
        RECT 633.000 493.800 635.100 495.900 ;
        RECT 633.300 492.000 635.100 493.800 ;
        RECT 641.700 495.600 658.500 496.800 ;
        RECT 659.400 495.600 660.300 498.600 ;
        RECT 664.800 495.900 666.600 496.800 ;
        RECT 674.100 496.500 675.900 498.300 ;
        RECT 692.100 497.100 693.600 500.400 ;
        RECT 667.800 495.900 669.900 496.050 ;
        RECT 630.900 490.200 633.300 491.100 ;
        RECT 631.800 490.050 633.300 490.200 ;
        RECT 637.800 490.950 639.900 493.050 ;
        RECT 627.000 487.500 630.900 489.300 ;
        RECT 628.800 487.200 630.900 487.500 ;
        RECT 631.800 487.950 633.900 490.050 ;
        RECT 637.800 489.150 639.600 490.950 ;
        RECT 631.800 486.000 632.700 487.950 ;
        RECT 625.500 483.600 627.600 485.700 ;
        RECT 631.200 484.950 632.700 486.000 ;
        RECT 631.200 483.600 632.400 484.950 ;
        RECT 602.700 478.500 606.300 479.400 ;
        RECT 623.100 482.700 627.600 483.600 ;
        RECT 602.700 477.600 603.600 478.500 ;
        RECT 598.500 471.000 600.300 477.600 ;
        RECT 601.500 476.700 603.600 477.600 ;
        RECT 601.500 471.600 603.300 476.700 ;
        RECT 604.500 471.000 606.300 477.600 ;
        RECT 623.100 471.600 624.900 482.700 ;
        RECT 626.100 471.000 627.900 481.500 ;
        RECT 630.600 471.600 632.400 483.600 ;
        RECT 635.100 483.600 637.200 484.500 ;
        RECT 635.100 482.400 639.900 483.600 ;
        RECT 635.100 471.000 636.900 481.500 ;
        RECT 638.100 471.600 639.900 482.400 ;
        RECT 641.700 479.400 642.900 495.600 ;
        RECT 659.400 493.800 661.200 495.600 ;
        RECT 664.800 495.000 669.900 495.900 ;
        RECT 667.800 493.950 669.900 495.000 ;
        RECT 674.100 495.900 676.200 496.500 ;
        RECT 674.100 494.400 691.200 495.900 ;
        RECT 692.100 495.300 699.900 497.100 ;
        RECT 689.700 492.900 696.300 494.400 ;
        RECT 644.100 491.700 688.500 492.900 ;
        RECT 644.100 490.050 645.900 491.700 ;
        RECT 643.800 487.950 645.900 490.050 ;
        RECT 649.800 489.750 651.900 490.050 ;
        RECT 662.400 489.900 664.200 490.500 ;
        RECT 671.400 489.900 684.900 490.800 ;
        RECT 649.800 487.950 653.700 489.750 ;
        RECT 662.400 488.700 673.500 489.900 ;
        RECT 651.900 487.200 653.700 487.950 ;
        RECT 671.400 487.800 673.500 488.700 ;
        RECT 675.000 487.200 678.900 489.000 ;
        RECT 684.000 488.700 684.900 489.900 ;
        RECT 651.900 486.300 665.400 487.200 ;
        RECT 676.800 486.900 678.900 487.200 ;
        RECT 683.100 486.900 684.900 488.700 ;
        RECT 687.600 490.200 688.500 491.700 ;
        RECT 687.600 488.400 692.700 490.200 ;
        RECT 694.800 490.050 696.300 492.900 ;
        RECT 694.800 487.950 696.900 490.050 ;
        RECT 664.200 485.700 665.400 486.300 ;
        RECT 698.100 485.700 699.900 486.300 ;
        RECT 659.400 484.500 661.500 484.800 ;
        RECT 664.200 484.500 699.900 485.700 ;
        RECT 649.500 483.300 661.500 484.500 ;
        RECT 700.800 483.600 701.700 500.400 ;
        RECT 649.500 482.700 651.300 483.300 ;
        RECT 659.400 482.700 661.500 483.300 ;
        RECT 664.200 482.400 681.900 483.600 ;
        RECT 646.200 481.800 648.000 482.100 ;
        RECT 664.200 481.800 665.400 482.400 ;
        RECT 646.200 480.600 665.400 481.800 ;
        RECT 679.800 481.500 681.900 482.400 ;
        RECT 685.200 482.700 701.700 483.600 ;
        RECT 685.200 481.500 687.300 482.700 ;
        RECT 646.200 480.300 648.000 480.600 ;
        RECT 641.700 478.500 645.300 479.400 ;
        RECT 644.400 477.600 645.300 478.500 ;
        RECT 641.700 471.000 643.500 477.600 ;
        RECT 644.400 476.700 646.500 477.600 ;
        RECT 644.700 471.600 646.500 476.700 ;
        RECT 647.700 471.000 649.500 477.600 ;
        RECT 650.700 471.600 652.500 480.600 ;
        RECT 662.700 477.600 664.800 479.700 ;
        RECT 670.200 479.100 673.500 481.200 ;
        RECT 653.700 471.000 655.500 477.600 ;
        RECT 657.300 474.600 659.400 476.700 ;
        RECT 660.300 474.600 662.400 476.700 ;
        RECT 657.300 471.600 659.100 474.600 ;
        RECT 660.300 471.600 662.100 474.600 ;
        RECT 663.300 471.600 665.100 477.600 ;
        RECT 666.300 471.000 668.100 477.600 ;
        RECT 670.200 471.600 672.000 479.100 ;
        RECT 676.200 477.600 678.900 481.500 ;
        RECT 691.200 480.600 696.900 481.800 ;
        RECT 688.500 479.700 690.300 480.300 ;
        RECT 682.200 478.500 690.300 479.700 ;
        RECT 682.200 477.600 684.300 478.500 ;
        RECT 691.200 477.600 692.400 480.600 ;
        RECT 695.100 480.000 696.900 480.600 ;
        RECT 700.800 479.400 701.700 482.700 ;
        RECT 697.800 478.500 701.700 479.400 ;
        RECT 703.500 503.400 705.300 506.400 ;
        RECT 706.500 503.400 708.300 507.000 ;
        RECT 703.500 490.050 705.000 503.400 ;
        RECT 725.100 500.400 726.900 507.000 ;
        RECT 728.100 499.500 729.900 506.400 ;
        RECT 731.100 500.400 732.900 507.000 ;
        RECT 734.100 499.500 735.900 506.400 ;
        RECT 737.100 500.400 738.900 507.000 ;
        RECT 740.100 499.500 741.900 506.400 ;
        RECT 743.100 500.400 744.900 507.000 ;
        RECT 746.100 499.500 747.900 506.400 ;
        RECT 749.100 500.400 750.900 507.000 ;
        RECT 752.700 500.400 754.500 506.400 ;
        RECT 758.100 500.400 759.900 507.000 ;
        RECT 763.500 500.400 765.300 506.400 ;
        RECT 767.700 503.400 769.500 506.400 ;
        RECT 770.700 503.400 772.500 506.400 ;
        RECT 773.700 503.400 775.500 506.400 ;
        RECT 776.700 503.400 778.500 507.000 ;
        RECT 767.700 501.300 769.800 503.400 ;
        RECT 770.700 501.300 772.800 503.400 ;
        RECT 773.700 501.300 775.800 503.400 ;
        RECT 781.200 502.500 783.000 506.400 ;
        RECT 784.200 503.400 786.000 507.000 ;
        RECT 787.200 503.400 789.000 506.400 ;
        RECT 790.200 503.400 792.000 506.400 ;
        RECT 793.200 503.400 795.000 506.400 ;
        RECT 796.200 503.400 798.000 506.400 ;
        RECT 777.600 501.600 779.400 502.500 ;
        RECT 776.700 500.400 779.400 501.600 ;
        RECT 781.200 500.400 783.900 502.500 ;
        RECT 787.200 501.300 789.300 503.400 ;
        RECT 790.200 501.300 792.300 503.400 ;
        RECT 793.200 501.300 795.300 503.400 ;
        RECT 796.200 501.300 798.300 503.400 ;
        RECT 800.400 501.600 802.200 506.400 ;
        RECT 800.400 500.400 804.600 501.600 ;
        RECT 805.500 500.400 807.300 507.000 ;
        RECT 810.900 500.400 812.700 506.400 ;
        RECT 727.050 498.300 729.900 499.500 ;
        RECT 732.000 498.300 735.900 499.500 ;
        RECT 738.000 498.300 741.900 499.500 ;
        RECT 744.000 498.300 747.900 499.500 ;
        RECT 727.050 493.050 728.100 498.300 ;
        RECT 732.000 497.400 733.200 498.300 ;
        RECT 738.000 497.400 739.200 498.300 ;
        RECT 744.000 497.400 745.200 498.300 ;
        RECT 729.000 496.200 733.200 497.400 ;
        RECT 729.000 495.600 730.800 496.200 ;
        RECT 727.050 490.950 730.200 493.050 ;
        RECT 703.500 487.950 705.900 490.050 ;
        RECT 697.800 477.600 699.000 478.500 ;
        RECT 703.500 477.600 705.000 487.950 ;
        RECT 727.050 485.700 728.100 490.950 ;
        RECT 732.000 485.700 733.200 496.200 ;
        RECT 735.000 496.200 739.200 497.400 ;
        RECT 735.000 495.600 736.800 496.200 ;
        RECT 738.000 485.700 739.200 496.200 ;
        RECT 741.000 496.200 745.200 497.400 ;
        RECT 741.000 495.600 742.800 496.200 ;
        RECT 744.000 485.700 745.200 496.200 ;
        RECT 752.700 496.800 753.900 500.400 ;
        RECT 763.800 499.500 765.300 500.400 ;
        RECT 772.800 499.800 774.600 500.400 ;
        RECT 776.700 499.800 777.600 500.400 ;
        RECT 756.900 498.300 765.300 499.500 ;
        RECT 770.400 498.600 777.600 499.800 ;
        RECT 792.300 498.600 798.900 500.400 ;
        RECT 756.900 497.700 758.700 498.300 ;
        RECT 767.400 496.800 769.500 497.700 ;
        RECT 752.700 495.600 769.500 496.800 ;
        RECT 770.400 495.600 771.300 498.600 ;
        RECT 775.800 495.900 777.600 496.800 ;
        RECT 785.100 496.500 786.900 498.300 ;
        RECT 803.100 497.100 804.600 500.400 ;
        RECT 778.800 495.900 780.900 496.050 ;
        RECT 746.400 493.050 748.200 494.850 ;
        RECT 746.100 490.950 748.200 493.050 ;
        RECT 727.050 484.500 729.900 485.700 ;
        RECT 732.000 484.500 735.900 485.700 ;
        RECT 738.000 484.500 741.900 485.700 ;
        RECT 744.000 484.500 747.900 485.700 ;
        RECT 673.200 471.000 675.000 477.600 ;
        RECT 676.200 471.600 678.000 477.600 ;
        RECT 679.200 474.600 681.300 476.700 ;
        RECT 682.200 474.600 684.300 476.700 ;
        RECT 685.200 474.600 687.300 476.700 ;
        RECT 679.200 471.600 681.000 474.600 ;
        RECT 682.200 471.600 684.000 474.600 ;
        RECT 685.200 471.600 687.000 474.600 ;
        RECT 688.200 471.000 690.000 477.600 ;
        RECT 691.200 471.600 693.000 477.600 ;
        RECT 694.200 471.000 696.000 477.600 ;
        RECT 697.200 471.600 699.000 477.600 ;
        RECT 700.200 471.000 702.000 477.600 ;
        RECT 703.500 471.600 705.300 477.600 ;
        RECT 706.500 471.000 708.300 477.600 ;
        RECT 725.100 471.000 726.900 483.600 ;
        RECT 728.100 471.600 729.900 484.500 ;
        RECT 731.100 471.000 732.900 483.600 ;
        RECT 734.100 471.600 735.900 484.500 ;
        RECT 737.100 471.000 738.900 483.600 ;
        RECT 740.100 471.600 741.900 484.500 ;
        RECT 743.100 471.000 744.900 483.600 ;
        RECT 746.100 471.600 747.900 484.500 ;
        RECT 749.100 471.000 750.900 483.600 ;
        RECT 752.700 479.400 753.900 495.600 ;
        RECT 770.400 493.800 772.200 495.600 ;
        RECT 775.800 495.000 780.900 495.900 ;
        RECT 778.800 493.950 780.900 495.000 ;
        RECT 785.100 495.900 787.200 496.500 ;
        RECT 785.100 494.400 802.200 495.900 ;
        RECT 803.100 495.300 810.900 497.100 ;
        RECT 800.700 492.900 807.300 494.400 ;
        RECT 755.100 491.700 799.500 492.900 ;
        RECT 755.100 490.050 756.900 491.700 ;
        RECT 754.800 487.950 756.900 490.050 ;
        RECT 760.800 489.750 762.900 490.050 ;
        RECT 773.400 489.900 775.200 490.500 ;
        RECT 782.400 489.900 795.900 490.800 ;
        RECT 760.800 487.950 764.700 489.750 ;
        RECT 773.400 488.700 784.500 489.900 ;
        RECT 762.900 487.200 764.700 487.950 ;
        RECT 782.400 487.800 784.500 488.700 ;
        RECT 786.000 487.200 789.900 489.000 ;
        RECT 795.000 488.700 795.900 489.900 ;
        RECT 762.900 486.300 776.400 487.200 ;
        RECT 787.800 486.900 789.900 487.200 ;
        RECT 794.100 486.900 795.900 488.700 ;
        RECT 798.600 490.200 799.500 491.700 ;
        RECT 798.600 488.400 803.700 490.200 ;
        RECT 805.800 490.050 807.300 492.900 ;
        RECT 805.800 487.950 807.900 490.050 ;
        RECT 775.200 485.700 776.400 486.300 ;
        RECT 809.100 485.700 810.900 486.300 ;
        RECT 770.400 484.500 772.500 484.800 ;
        RECT 775.200 484.500 810.900 485.700 ;
        RECT 760.500 483.300 772.500 484.500 ;
        RECT 811.800 483.600 812.700 500.400 ;
        RECT 760.500 482.700 762.300 483.300 ;
        RECT 770.400 482.700 772.500 483.300 ;
        RECT 775.200 482.400 792.900 483.600 ;
        RECT 757.200 481.800 759.000 482.100 ;
        RECT 775.200 481.800 776.400 482.400 ;
        RECT 757.200 480.600 776.400 481.800 ;
        RECT 790.800 481.500 792.900 482.400 ;
        RECT 796.200 482.700 812.700 483.600 ;
        RECT 796.200 481.500 798.300 482.700 ;
        RECT 757.200 480.300 759.000 480.600 ;
        RECT 752.700 478.500 756.300 479.400 ;
        RECT 755.400 477.600 756.300 478.500 ;
        RECT 752.700 471.000 754.500 477.600 ;
        RECT 755.400 476.700 757.500 477.600 ;
        RECT 755.700 471.600 757.500 476.700 ;
        RECT 758.700 471.000 760.500 477.600 ;
        RECT 761.700 471.600 763.500 480.600 ;
        RECT 773.700 477.600 775.800 479.700 ;
        RECT 781.200 479.100 784.500 481.200 ;
        RECT 764.700 471.000 766.500 477.600 ;
        RECT 768.300 474.600 770.400 476.700 ;
        RECT 771.300 474.600 773.400 476.700 ;
        RECT 768.300 471.600 770.100 474.600 ;
        RECT 771.300 471.600 773.100 474.600 ;
        RECT 774.300 471.600 776.100 477.600 ;
        RECT 777.300 471.000 779.100 477.600 ;
        RECT 781.200 471.600 783.000 479.100 ;
        RECT 787.200 477.600 789.900 481.500 ;
        RECT 802.200 480.600 807.900 481.800 ;
        RECT 799.500 479.700 801.300 480.300 ;
        RECT 793.200 478.500 801.300 479.700 ;
        RECT 793.200 477.600 795.300 478.500 ;
        RECT 802.200 477.600 803.400 480.600 ;
        RECT 806.100 480.000 807.900 480.600 ;
        RECT 811.800 479.400 812.700 482.700 ;
        RECT 808.800 478.500 812.700 479.400 ;
        RECT 814.500 503.400 816.300 506.400 ;
        RECT 817.500 503.400 819.300 507.000 ;
        RECT 836.100 503.400 837.900 507.000 ;
        RECT 839.100 503.400 840.900 506.400 ;
        RECT 857.100 503.400 858.900 507.000 ;
        RECT 860.100 503.400 861.900 506.400 ;
        RECT 863.100 503.400 864.900 507.000 ;
        RECT 814.500 490.050 816.000 503.400 ;
        RECT 820.950 498.450 823.050 499.050 ;
        RECT 835.950 498.450 838.050 498.900 ;
        RECT 820.950 497.550 838.050 498.450 ;
        RECT 820.950 496.950 823.050 497.550 ;
        RECT 835.950 496.800 838.050 497.550 ;
        RECT 817.800 493.950 819.900 496.050 ;
        RECT 820.950 495.450 823.050 495.900 ;
        RECT 832.950 495.450 835.050 496.050 ;
        RECT 820.950 494.550 835.050 495.450 ;
        RECT 814.500 487.950 816.900 490.050 ;
        RECT 818.550 489.450 819.450 493.950 ;
        RECT 820.950 493.800 823.050 494.550 ;
        RECT 832.950 493.950 835.050 494.550 ;
        RECT 839.100 493.050 840.300 503.400 ;
        RECT 860.400 493.050 861.300 503.400 ;
        RECT 866.700 500.400 868.500 506.400 ;
        RECT 872.100 500.400 873.900 507.000 ;
        RECT 877.500 500.400 879.300 506.400 ;
        RECT 881.700 503.400 883.500 506.400 ;
        RECT 884.700 503.400 886.500 506.400 ;
        RECT 887.700 503.400 889.500 506.400 ;
        RECT 890.700 503.400 892.500 507.000 ;
        RECT 881.700 501.300 883.800 503.400 ;
        RECT 884.700 501.300 886.800 503.400 ;
        RECT 887.700 501.300 889.800 503.400 ;
        RECT 895.200 502.500 897.000 506.400 ;
        RECT 898.200 503.400 900.000 507.000 ;
        RECT 901.200 503.400 903.000 506.400 ;
        RECT 904.200 503.400 906.000 506.400 ;
        RECT 907.200 503.400 909.000 506.400 ;
        RECT 910.200 503.400 912.000 506.400 ;
        RECT 891.600 501.600 893.400 502.500 ;
        RECT 890.700 500.400 893.400 501.600 ;
        RECT 895.200 500.400 897.900 502.500 ;
        RECT 901.200 501.300 903.300 503.400 ;
        RECT 904.200 501.300 906.300 503.400 ;
        RECT 907.200 501.300 909.300 503.400 ;
        RECT 910.200 501.300 912.300 503.400 ;
        RECT 914.400 501.600 916.200 506.400 ;
        RECT 914.400 500.400 918.600 501.600 ;
        RECT 919.500 500.400 921.300 507.000 ;
        RECT 924.900 500.400 926.700 506.400 ;
        RECT 866.700 496.800 867.900 500.400 ;
        RECT 877.800 499.500 879.300 500.400 ;
        RECT 886.800 499.800 888.600 500.400 ;
        RECT 890.700 499.800 891.600 500.400 ;
        RECT 870.900 498.300 879.300 499.500 ;
        RECT 884.400 498.600 891.600 499.800 ;
        RECT 906.300 498.600 912.900 500.400 ;
        RECT 870.900 497.700 872.700 498.300 ;
        RECT 881.400 496.800 883.500 497.700 ;
        RECT 866.700 495.600 883.500 496.800 ;
        RECT 884.400 495.600 885.300 498.600 ;
        RECT 889.800 495.900 891.600 496.800 ;
        RECT 899.100 496.500 900.900 498.300 ;
        RECT 917.100 497.100 918.600 500.400 ;
        RECT 892.800 495.900 894.900 496.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 832.950 489.450 835.050 490.050 ;
        RECT 818.550 488.550 835.050 489.450 ;
        RECT 836.100 489.150 837.900 490.950 ;
        RECT 832.950 487.950 835.050 488.550 ;
        RECT 808.800 477.600 810.000 478.500 ;
        RECT 814.500 477.600 816.000 487.950 ;
        RECT 839.100 477.600 840.300 490.950 ;
        RECT 857.250 489.150 859.050 490.950 ;
        RECT 850.950 486.450 853.050 487.050 ;
        RECT 856.950 486.450 859.050 487.050 ;
        RECT 850.950 485.550 859.050 486.450 ;
        RECT 850.950 484.950 853.050 485.550 ;
        RECT 856.950 484.950 859.050 485.550 ;
        RECT 860.400 483.600 861.300 490.950 ;
        RECT 863.100 489.150 864.900 490.950 ;
        RECT 784.200 471.000 786.000 477.600 ;
        RECT 787.200 471.600 789.000 477.600 ;
        RECT 790.200 474.600 792.300 476.700 ;
        RECT 793.200 474.600 795.300 476.700 ;
        RECT 796.200 474.600 798.300 476.700 ;
        RECT 790.200 471.600 792.000 474.600 ;
        RECT 793.200 471.600 795.000 474.600 ;
        RECT 796.200 471.600 798.000 474.600 ;
        RECT 799.200 471.000 801.000 477.600 ;
        RECT 802.200 471.600 804.000 477.600 ;
        RECT 805.200 471.000 807.000 477.600 ;
        RECT 808.200 471.600 810.000 477.600 ;
        RECT 811.200 471.000 813.000 477.600 ;
        RECT 814.500 471.600 816.300 477.600 ;
        RECT 817.500 471.000 819.300 477.600 ;
        RECT 836.100 471.000 837.900 477.600 ;
        RECT 839.100 471.600 840.900 477.600 ;
        RECT 857.100 471.000 858.900 483.600 ;
        RECT 860.400 482.400 864.000 483.600 ;
        RECT 862.200 471.600 864.000 482.400 ;
        RECT 866.700 479.400 867.900 495.600 ;
        RECT 884.400 493.800 886.200 495.600 ;
        RECT 889.800 495.000 894.900 495.900 ;
        RECT 892.800 493.950 894.900 495.000 ;
        RECT 899.100 495.900 901.200 496.500 ;
        RECT 899.100 494.400 916.200 495.900 ;
        RECT 917.100 495.300 924.900 497.100 ;
        RECT 914.700 492.900 921.300 494.400 ;
        RECT 869.100 491.700 913.500 492.900 ;
        RECT 869.100 490.050 870.900 491.700 ;
        RECT 868.800 487.950 870.900 490.050 ;
        RECT 874.800 489.750 876.900 490.050 ;
        RECT 887.400 489.900 889.200 490.500 ;
        RECT 896.400 489.900 909.900 490.800 ;
        RECT 874.800 487.950 878.700 489.750 ;
        RECT 887.400 488.700 898.500 489.900 ;
        RECT 876.900 487.200 878.700 487.950 ;
        RECT 896.400 487.800 898.500 488.700 ;
        RECT 900.000 487.200 903.900 489.000 ;
        RECT 909.000 488.700 909.900 489.900 ;
        RECT 876.900 486.300 890.400 487.200 ;
        RECT 901.800 486.900 903.900 487.200 ;
        RECT 908.100 486.900 909.900 488.700 ;
        RECT 912.600 490.200 913.500 491.700 ;
        RECT 912.600 488.400 917.700 490.200 ;
        RECT 919.800 490.050 921.300 492.900 ;
        RECT 919.800 487.950 921.900 490.050 ;
        RECT 889.200 485.700 890.400 486.300 ;
        RECT 923.100 485.700 924.900 486.300 ;
        RECT 884.400 484.500 886.500 484.800 ;
        RECT 889.200 484.500 924.900 485.700 ;
        RECT 874.500 483.300 886.500 484.500 ;
        RECT 925.800 483.600 926.700 500.400 ;
        RECT 874.500 482.700 876.300 483.300 ;
        RECT 884.400 482.700 886.500 483.300 ;
        RECT 889.200 482.400 906.900 483.600 ;
        RECT 871.200 481.800 873.000 482.100 ;
        RECT 889.200 481.800 890.400 482.400 ;
        RECT 871.200 480.600 890.400 481.800 ;
        RECT 904.800 481.500 906.900 482.400 ;
        RECT 910.200 482.700 926.700 483.600 ;
        RECT 910.200 481.500 912.300 482.700 ;
        RECT 871.200 480.300 873.000 480.600 ;
        RECT 866.700 478.500 870.300 479.400 ;
        RECT 869.400 477.600 870.300 478.500 ;
        RECT 866.700 471.000 868.500 477.600 ;
        RECT 869.400 476.700 871.500 477.600 ;
        RECT 869.700 471.600 871.500 476.700 ;
        RECT 872.700 471.000 874.500 477.600 ;
        RECT 875.700 471.600 877.500 480.600 ;
        RECT 887.700 477.600 889.800 479.700 ;
        RECT 895.200 479.100 898.500 481.200 ;
        RECT 878.700 471.000 880.500 477.600 ;
        RECT 882.300 474.600 884.400 476.700 ;
        RECT 885.300 474.600 887.400 476.700 ;
        RECT 882.300 471.600 884.100 474.600 ;
        RECT 885.300 471.600 887.100 474.600 ;
        RECT 888.300 471.600 890.100 477.600 ;
        RECT 891.300 471.000 893.100 477.600 ;
        RECT 895.200 471.600 897.000 479.100 ;
        RECT 901.200 477.600 903.900 481.500 ;
        RECT 916.200 480.600 921.900 481.800 ;
        RECT 913.500 479.700 915.300 480.300 ;
        RECT 907.200 478.500 915.300 479.700 ;
        RECT 907.200 477.600 909.300 478.500 ;
        RECT 916.200 477.600 917.400 480.600 ;
        RECT 920.100 480.000 921.900 480.600 ;
        RECT 925.800 479.400 926.700 482.700 ;
        RECT 922.800 478.500 926.700 479.400 ;
        RECT 928.500 503.400 930.300 506.400 ;
        RECT 931.500 503.400 933.300 507.000 ;
        RECT 928.500 490.050 930.000 503.400 ;
        RECT 950.100 500.400 951.900 507.000 ;
        RECT 953.100 500.400 954.900 506.400 ;
        RECT 971.100 503.400 972.900 507.000 ;
        RECT 974.100 503.400 975.900 506.400 ;
        RECT 977.100 503.400 978.900 507.000 ;
        RECT 982.950 504.450 985.050 505.050 ;
        RECT 991.950 504.450 994.050 505.050 ;
        RECT 982.950 503.550 994.050 504.450 ;
        RECT 961.950 501.450 964.050 502.050 ;
        RECT 961.950 501.000 972.450 501.450 ;
        RECT 961.950 500.550 973.050 501.000 ;
        RECT 950.100 493.050 951.900 494.850 ;
        RECT 953.100 493.050 954.300 500.400 ;
        RECT 961.950 499.950 964.050 500.550 ;
        RECT 970.950 496.800 973.050 500.550 ;
        RECT 955.950 495.450 960.000 496.050 ;
        RECT 961.950 495.450 964.050 496.050 ;
        RECT 967.950 495.450 970.050 496.050 ;
        RECT 955.950 493.950 960.450 495.450 ;
        RECT 961.950 494.550 970.050 495.450 ;
        RECT 961.950 493.950 964.050 494.550 ;
        RECT 967.950 493.950 970.050 494.550 ;
        RECT 949.950 490.950 952.050 493.050 ;
        RECT 952.950 490.950 955.050 493.050 ;
        RECT 959.550 492.450 960.450 493.950 ;
        RECT 974.700 493.050 975.600 503.400 ;
        RECT 982.950 502.950 985.050 503.550 ;
        RECT 991.950 502.950 994.050 503.550 ;
        RECT 995.100 500.400 996.900 506.400 ;
        RECT 995.700 498.300 996.900 500.400 ;
        RECT 998.100 501.300 999.900 506.400 ;
        RECT 1001.100 502.200 1002.900 507.000 ;
        RECT 1004.100 501.300 1005.900 506.400 ;
        RECT 998.100 499.950 1005.900 501.300 ;
        RECT 1022.100 500.400 1023.900 506.400 ;
        RECT 1025.100 500.400 1026.900 507.000 ;
        RECT 995.700 497.400 999.300 498.300 ;
        RECT 995.100 493.050 996.900 494.850 ;
        RECT 998.100 493.050 999.300 497.400 ;
        RECT 1001.100 493.050 1002.900 494.850 ;
        RECT 1022.700 493.050 1023.900 500.400 ;
        RECT 1025.100 493.050 1026.900 494.850 ;
        RECT 959.550 491.550 966.450 492.450 ;
        RECT 928.500 487.950 930.900 490.050 ;
        RECT 922.800 477.600 924.000 478.500 ;
        RECT 928.500 477.600 930.000 487.950 ;
        RECT 934.950 486.450 937.050 487.050 ;
        RECT 940.950 486.450 943.050 487.050 ;
        RECT 934.950 485.550 943.050 486.450 ;
        RECT 934.950 484.950 937.050 485.550 ;
        RECT 940.950 484.950 943.050 485.550 ;
        RECT 953.100 483.600 954.300 490.950 ;
        RECT 965.550 490.050 966.450 491.550 ;
        RECT 970.950 490.950 973.050 493.050 ;
        RECT 973.950 490.950 976.050 493.050 ;
        RECT 976.950 490.950 979.050 493.050 ;
        RECT 994.950 490.950 997.050 493.050 ;
        RECT 997.950 490.950 1000.050 493.050 ;
        RECT 1000.950 490.950 1003.050 493.050 ;
        RECT 1003.950 490.950 1006.050 493.050 ;
        RECT 1021.950 490.950 1024.050 493.050 ;
        RECT 1024.950 490.950 1027.050 493.050 ;
        RECT 965.550 488.550 970.050 490.050 ;
        RECT 971.100 489.150 972.900 490.950 ;
        RECT 966.000 487.950 970.050 488.550 ;
        RECT 974.700 483.600 975.600 490.950 ;
        RECT 976.950 489.150 978.750 490.950 ;
        RECT 998.100 483.600 999.300 490.950 ;
        RECT 1004.100 489.150 1005.900 490.950 ;
        RECT 1022.700 483.600 1023.900 490.950 ;
        RECT 898.200 471.000 900.000 477.600 ;
        RECT 901.200 471.600 903.000 477.600 ;
        RECT 904.200 474.600 906.300 476.700 ;
        RECT 907.200 474.600 909.300 476.700 ;
        RECT 910.200 474.600 912.300 476.700 ;
        RECT 904.200 471.600 906.000 474.600 ;
        RECT 907.200 471.600 909.000 474.600 ;
        RECT 910.200 471.600 912.000 474.600 ;
        RECT 913.200 471.000 915.000 477.600 ;
        RECT 916.200 471.600 918.000 477.600 ;
        RECT 919.200 471.000 921.000 477.600 ;
        RECT 922.200 471.600 924.000 477.600 ;
        RECT 925.200 471.000 927.000 477.600 ;
        RECT 928.500 471.600 930.300 477.600 ;
        RECT 931.500 471.000 933.300 477.600 ;
        RECT 950.100 471.000 951.900 483.600 ;
        RECT 953.100 471.600 954.900 483.600 ;
        RECT 972.000 482.400 975.600 483.600 ;
        RECT 972.000 471.600 973.800 482.400 ;
        RECT 977.100 471.000 978.900 483.600 ;
        RECT 998.100 482.100 1000.500 483.600 ;
        RECT 996.000 479.100 997.800 480.900 ;
        RECT 995.700 471.000 997.500 477.600 ;
        RECT 998.700 471.600 1000.500 482.100 ;
        RECT 1003.800 471.000 1005.600 483.600 ;
        RECT 1022.100 471.600 1023.900 483.600 ;
        RECT 1025.100 471.000 1026.900 483.600 ;
        RECT 2.700 461.400 4.500 468.000 ;
        RECT 5.700 462.300 7.500 467.400 ;
        RECT 5.400 461.400 7.500 462.300 ;
        RECT 8.700 461.400 10.500 468.000 ;
        RECT 5.400 460.500 6.300 461.400 ;
        RECT 2.700 459.600 6.300 460.500 ;
        RECT 2.700 443.400 3.900 459.600 ;
        RECT 7.200 458.400 9.000 458.700 ;
        RECT 11.700 458.400 13.500 467.400 ;
        RECT 14.700 461.400 16.500 468.000 ;
        RECT 18.300 464.400 20.100 467.400 ;
        RECT 21.300 464.400 23.100 467.400 ;
        RECT 18.300 462.300 20.400 464.400 ;
        RECT 21.300 462.300 23.400 464.400 ;
        RECT 24.300 461.400 26.100 467.400 ;
        RECT 27.300 461.400 29.100 468.000 ;
        RECT 23.700 459.300 25.800 461.400 ;
        RECT 31.200 459.900 33.000 467.400 ;
        RECT 34.200 461.400 36.000 468.000 ;
        RECT 37.200 461.400 39.000 467.400 ;
        RECT 40.200 464.400 42.000 467.400 ;
        RECT 43.200 464.400 45.000 467.400 ;
        RECT 46.200 464.400 48.000 467.400 ;
        RECT 40.200 462.300 42.300 464.400 ;
        RECT 43.200 462.300 45.300 464.400 ;
        RECT 46.200 462.300 48.300 464.400 ;
        RECT 49.200 461.400 51.000 468.000 ;
        RECT 52.200 461.400 54.000 467.400 ;
        RECT 55.200 461.400 57.000 468.000 ;
        RECT 58.200 461.400 60.000 467.400 ;
        RECT 61.200 461.400 63.000 468.000 ;
        RECT 64.500 461.400 66.300 467.400 ;
        RECT 67.500 461.400 69.300 468.000 ;
        RECT 86.100 461.400 87.900 468.000 ;
        RECT 89.100 461.400 90.900 467.400 ;
        RECT 107.100 461.400 108.900 467.400 ;
        RECT 110.100 462.000 111.900 468.000 ;
        RECT 7.200 457.200 26.400 458.400 ;
        RECT 31.200 457.800 34.500 459.900 ;
        RECT 37.200 457.500 39.900 461.400 ;
        RECT 43.200 460.500 45.300 461.400 ;
        RECT 43.200 459.300 51.300 460.500 ;
        RECT 49.500 458.700 51.300 459.300 ;
        RECT 52.200 458.400 53.400 461.400 ;
        RECT 58.800 460.500 60.000 461.400 ;
        RECT 58.800 459.600 62.700 460.500 ;
        RECT 56.100 458.400 57.900 459.000 ;
        RECT 7.200 456.900 9.000 457.200 ;
        RECT 25.200 456.600 26.400 457.200 ;
        RECT 40.800 456.600 42.900 457.500 ;
        RECT 10.500 455.700 12.300 456.300 ;
        RECT 20.400 455.700 22.500 456.300 ;
        RECT 10.500 454.500 22.500 455.700 ;
        RECT 25.200 455.400 42.900 456.600 ;
        RECT 46.200 456.300 48.300 457.500 ;
        RECT 52.200 457.200 57.900 458.400 ;
        RECT 61.800 456.300 62.700 459.600 ;
        RECT 46.200 455.400 62.700 456.300 ;
        RECT 20.400 454.200 22.500 454.500 ;
        RECT 25.200 453.300 60.900 454.500 ;
        RECT 25.200 452.700 26.400 453.300 ;
        RECT 59.100 452.700 60.900 453.300 ;
        RECT 12.900 451.800 26.400 452.700 ;
        RECT 37.800 451.800 39.900 452.100 ;
        RECT 12.900 451.050 14.700 451.800 ;
        RECT 4.800 448.950 6.900 451.050 ;
        RECT 10.800 449.250 14.700 451.050 ;
        RECT 32.400 450.300 34.500 451.200 ;
        RECT 10.800 448.950 12.900 449.250 ;
        RECT 23.400 449.100 34.500 450.300 ;
        RECT 36.000 450.000 39.900 451.800 ;
        RECT 44.100 450.300 45.900 452.100 ;
        RECT 45.000 449.100 45.900 450.300 ;
        RECT 5.100 447.300 6.900 448.950 ;
        RECT 23.400 448.500 25.200 449.100 ;
        RECT 32.400 448.200 45.900 449.100 ;
        RECT 48.600 448.800 53.700 450.600 ;
        RECT 55.800 448.950 57.900 451.050 ;
        RECT 48.600 447.300 49.500 448.800 ;
        RECT 5.100 446.100 49.500 447.300 ;
        RECT 55.800 446.100 57.300 448.950 ;
        RECT 20.400 443.400 22.200 445.200 ;
        RECT 28.800 444.000 30.900 445.050 ;
        RECT 50.700 444.600 57.300 446.100 ;
        RECT 2.700 442.200 19.500 443.400 ;
        RECT 2.700 438.600 3.900 442.200 ;
        RECT 17.400 441.300 19.500 442.200 ;
        RECT 6.900 440.700 8.700 441.300 ;
        RECT 6.900 439.500 15.300 440.700 ;
        RECT 13.800 438.600 15.300 439.500 ;
        RECT 20.400 440.400 21.300 443.400 ;
        RECT 25.800 443.100 30.900 444.000 ;
        RECT 25.800 442.200 27.600 443.100 ;
        RECT 28.800 442.950 30.900 443.100 ;
        RECT 35.100 443.100 52.200 444.600 ;
        RECT 35.100 442.500 37.200 443.100 ;
        RECT 35.100 440.700 36.900 442.500 ;
        RECT 53.100 441.900 60.900 443.700 ;
        RECT 20.400 439.200 27.600 440.400 ;
        RECT 22.800 438.600 24.600 439.200 ;
        RECT 26.700 438.600 27.600 439.200 ;
        RECT 42.300 438.600 48.900 440.400 ;
        RECT 53.100 438.600 54.600 441.900 ;
        RECT 61.800 438.600 62.700 455.400 ;
        RECT 2.700 432.600 4.500 438.600 ;
        RECT 8.100 432.000 9.900 438.600 ;
        RECT 13.500 432.600 15.300 438.600 ;
        RECT 17.700 435.600 19.800 437.700 ;
        RECT 20.700 435.600 22.800 437.700 ;
        RECT 23.700 435.600 25.800 437.700 ;
        RECT 26.700 437.400 29.400 438.600 ;
        RECT 27.600 436.500 29.400 437.400 ;
        RECT 31.200 436.500 33.900 438.600 ;
        RECT 17.700 432.600 19.500 435.600 ;
        RECT 20.700 432.600 22.500 435.600 ;
        RECT 23.700 432.600 25.500 435.600 ;
        RECT 26.700 432.000 28.500 435.600 ;
        RECT 31.200 432.600 33.000 436.500 ;
        RECT 37.200 435.600 39.300 437.700 ;
        RECT 40.200 435.600 42.300 437.700 ;
        RECT 43.200 435.600 45.300 437.700 ;
        RECT 46.200 435.600 48.300 437.700 ;
        RECT 50.400 437.400 54.600 438.600 ;
        RECT 34.200 432.000 36.000 435.600 ;
        RECT 37.200 432.600 39.000 435.600 ;
        RECT 40.200 432.600 42.000 435.600 ;
        RECT 43.200 432.600 45.000 435.600 ;
        RECT 46.200 432.600 48.000 435.600 ;
        RECT 50.400 432.600 52.200 437.400 ;
        RECT 55.500 432.000 57.300 438.600 ;
        RECT 60.900 432.600 62.700 438.600 ;
        RECT 64.500 451.050 66.000 461.400 ;
        RECT 64.500 448.950 66.900 451.050 ;
        RECT 64.500 435.600 66.000 448.950 ;
        RECT 86.100 448.050 87.900 449.850 ;
        RECT 89.100 448.050 90.300 461.400 ;
        RECT 108.000 461.100 108.900 461.400 ;
        RECT 113.100 461.400 114.900 467.400 ;
        RECT 116.100 461.400 117.900 468.000 ;
        RECT 113.100 461.100 114.600 461.400 ;
        RECT 108.000 460.200 114.600 461.100 ;
        RECT 108.000 448.050 108.900 460.200 ;
        RECT 135.000 456.600 136.800 467.400 ;
        RECT 135.000 455.400 138.600 456.600 ;
        RECT 140.100 455.400 141.900 468.000 ;
        RECT 158.700 461.400 160.500 468.000 ;
        RECT 159.000 458.100 160.800 459.900 ;
        RECT 161.700 456.900 163.500 467.400 ;
        RECT 161.100 455.400 163.500 456.900 ;
        RECT 166.800 455.400 168.600 468.000 ;
        RECT 185.100 461.400 186.900 468.000 ;
        RECT 188.100 461.400 189.900 467.400 ;
        RECT 191.100 461.400 192.900 468.000 ;
        RECT 113.100 448.050 114.900 449.850 ;
        RECT 134.100 448.050 135.900 449.850 ;
        RECT 137.700 448.050 138.600 455.400 ;
        RECT 139.950 448.050 141.750 449.850 ;
        RECT 161.100 448.050 162.300 455.400 ;
        RECT 167.100 448.050 168.900 449.850 ;
        RECT 188.100 448.050 189.300 461.400 ;
        RECT 209.100 455.400 210.900 468.000 ;
        RECT 212.100 454.500 213.900 467.400 ;
        RECT 215.100 455.400 216.900 468.000 ;
        RECT 218.100 455.400 219.900 467.400 ;
        RECT 221.100 455.400 222.900 468.000 ;
        RECT 239.400 455.400 241.200 468.000 ;
        RECT 244.500 456.900 246.300 467.400 ;
        RECT 247.500 461.400 249.300 468.000 ;
        RECT 247.200 458.100 249.000 459.900 ;
        RECT 244.500 455.400 246.900 456.900 ;
        RECT 266.100 455.400 267.900 468.000 ;
        RECT 271.200 456.600 273.000 467.400 ;
        RECT 269.400 455.400 273.000 456.600 ;
        RECT 290.100 455.400 291.900 468.000 ;
        RECT 295.200 456.600 297.000 467.400 ;
        RECT 293.400 455.400 297.000 456.600 ;
        RECT 315.000 456.600 316.800 467.400 ;
        RECT 315.000 455.400 318.600 456.600 ;
        RECT 320.100 455.400 321.900 468.000 ;
        RECT 338.100 461.400 339.900 468.000 ;
        RECT 341.100 461.400 342.900 467.400 ;
        RECT 359.100 461.400 360.900 468.000 ;
        RECT 362.100 461.400 363.900 467.400 ;
        RECT 365.100 461.400 366.900 468.000 ;
        RECT 383.100 461.400 384.900 468.000 ;
        RECT 386.100 461.400 387.900 467.400 ;
        RECT 389.100 462.000 390.900 468.000 ;
        RECT 218.100 454.500 219.300 455.400 ;
        RECT 212.100 453.600 219.300 454.500 ;
        RECT 212.100 448.050 213.900 449.850 ;
        RECT 218.100 448.050 219.300 453.600 ;
        RECT 239.100 448.050 240.900 449.850 ;
        RECT 245.700 448.050 246.900 455.400 ;
        RECT 266.250 448.050 268.050 449.850 ;
        RECT 269.400 448.050 270.300 455.400 ;
        RECT 272.100 448.050 273.900 449.850 ;
        RECT 290.250 448.050 292.050 449.850 ;
        RECT 293.400 448.050 294.300 455.400 ;
        RECT 296.100 448.050 297.900 449.850 ;
        RECT 314.100 448.050 315.900 449.850 ;
        RECT 317.700 448.050 318.600 455.400 ;
        RECT 319.950 453.450 322.050 454.050 ;
        RECT 325.950 453.450 328.050 454.050 ;
        RECT 319.950 452.550 328.050 453.450 ;
        RECT 319.950 451.950 322.050 452.550 ;
        RECT 325.950 451.950 328.050 452.550 ;
        RECT 319.950 448.050 321.750 449.850 ;
        RECT 338.100 448.050 339.900 449.850 ;
        RECT 341.100 448.050 342.300 461.400 ;
        RECT 362.700 448.050 363.900 461.400 ;
        RECT 386.400 461.100 387.900 461.400 ;
        RECT 392.100 461.400 393.900 467.400 ;
        RECT 410.100 461.400 411.900 468.000 ;
        RECT 413.100 461.400 414.900 467.400 ;
        RECT 416.100 461.400 417.900 468.000 ;
        RECT 392.100 461.100 393.000 461.400 ;
        RECT 386.400 460.200 393.000 461.100 ;
        RECT 373.950 456.450 376.050 457.050 ;
        RECT 379.950 456.450 382.050 457.050 ;
        RECT 373.950 455.550 382.050 456.450 ;
        RECT 373.950 454.950 376.050 455.550 ;
        RECT 379.950 454.950 382.050 455.550 ;
        RECT 386.100 448.050 387.900 449.850 ;
        RECT 392.100 448.050 393.000 460.200 ;
        RECT 413.100 448.050 414.300 461.400 ;
        RECT 435.000 456.600 436.800 467.400 ;
        RECT 435.000 455.400 438.600 456.600 ;
        RECT 440.100 455.400 441.900 468.000 ;
        RECT 458.400 455.400 460.200 468.000 ;
        RECT 463.500 456.900 465.300 467.400 ;
        RECT 466.500 461.400 468.300 468.000 ;
        RECT 485.100 461.400 486.900 468.000 ;
        RECT 488.100 461.400 489.900 467.400 ;
        RECT 491.100 461.400 492.900 468.000 ;
        RECT 509.100 461.400 510.900 468.000 ;
        RECT 512.100 461.400 513.900 467.400 ;
        RECT 515.100 461.400 516.900 468.000 ;
        RECT 533.100 461.400 534.900 468.000 ;
        RECT 536.100 461.400 537.900 467.400 ;
        RECT 539.100 462.000 540.900 468.000 ;
        RECT 466.200 458.100 468.000 459.900 ;
        RECT 463.500 455.400 465.900 456.900 ;
        RECT 421.950 453.450 424.050 454.050 ;
        RECT 427.950 453.450 430.050 454.050 ;
        RECT 421.950 452.550 430.050 453.450 ;
        RECT 421.950 451.950 424.050 452.550 ;
        RECT 427.950 451.950 430.050 452.550 ;
        RECT 434.100 448.050 435.900 449.850 ;
        RECT 437.700 448.050 438.600 455.400 ;
        RECT 451.950 453.450 454.050 454.050 ;
        RECT 460.950 453.450 463.050 454.050 ;
        RECT 451.950 452.550 463.050 453.450 ;
        RECT 451.950 451.950 454.050 452.550 ;
        RECT 460.950 451.950 463.050 452.550 ;
        RECT 439.950 448.050 441.750 449.850 ;
        RECT 458.100 448.050 459.900 449.850 ;
        RECT 464.700 448.050 465.900 455.400 ;
        RECT 488.700 448.050 489.900 461.400 ;
        RECT 496.950 453.450 499.050 454.050 ;
        RECT 508.950 453.450 511.050 454.050 ;
        RECT 496.950 452.550 511.050 453.450 ;
        RECT 496.950 451.950 499.050 452.550 ;
        RECT 508.950 451.950 511.050 452.550 ;
        RECT 512.700 448.050 513.900 461.400 ;
        RECT 536.400 461.100 537.900 461.400 ;
        RECT 542.100 461.400 543.900 467.400 ;
        RECT 560.700 461.400 562.500 468.000 ;
        RECT 542.100 461.100 543.000 461.400 ;
        RECT 536.400 460.200 543.000 461.100 ;
        RECT 536.100 448.050 537.900 449.850 ;
        RECT 542.100 448.050 543.000 460.200 ;
        RECT 561.000 458.100 562.800 459.900 ;
        RECT 563.700 456.900 565.500 467.400 ;
        RECT 563.100 455.400 565.500 456.900 ;
        RECT 568.800 455.400 570.600 468.000 ;
        RECT 587.100 455.400 588.900 468.000 ;
        RECT 592.200 456.600 594.000 467.400 ;
        RECT 611.700 461.400 613.500 468.000 ;
        RECT 612.000 458.100 613.800 459.900 ;
        RECT 614.700 456.900 616.500 467.400 ;
        RECT 590.400 455.400 594.000 456.600 ;
        RECT 614.100 455.400 616.500 456.900 ;
        RECT 619.800 455.400 621.600 468.000 ;
        RECT 638.100 461.400 639.900 468.000 ;
        RECT 641.100 461.400 642.900 467.400 ;
        RECT 563.100 448.050 564.300 455.400 ;
        RECT 569.100 448.050 570.900 449.850 ;
        RECT 587.250 448.050 589.050 449.850 ;
        RECT 590.400 448.050 591.300 455.400 ;
        RECT 593.100 448.050 594.900 449.850 ;
        RECT 614.100 448.050 615.300 455.400 ;
        RECT 620.100 448.050 621.900 449.850 ;
        RECT 638.100 448.050 639.900 449.850 ;
        RECT 641.100 448.050 642.300 461.400 ;
        RECT 659.100 456.300 660.900 467.400 ;
        RECT 662.100 457.200 663.900 468.000 ;
        RECT 665.100 456.300 666.900 467.400 ;
        RECT 659.100 455.400 666.900 456.300 ;
        RECT 668.100 455.400 669.900 467.400 ;
        RECT 686.100 461.400 687.900 468.000 ;
        RECT 689.100 461.400 690.900 467.400 ;
        RECT 692.100 461.400 693.900 468.000 ;
        RECT 646.950 453.450 649.050 454.050 ;
        RECT 658.950 453.450 661.050 454.050 ;
        RECT 646.950 452.550 661.050 453.450 ;
        RECT 646.950 451.950 649.050 452.550 ;
        RECT 658.950 451.950 661.050 452.550 ;
        RECT 662.250 448.050 664.050 449.850 ;
        RECT 668.700 448.050 669.600 455.400 ;
        RECT 681.000 450.450 685.050 451.050 ;
        RECT 680.550 450.000 685.050 450.450 ;
        RECT 679.950 448.950 685.050 450.000 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 190.950 445.950 193.050 448.050 ;
        RECT 212.100 445.950 214.200 448.050 ;
        RECT 218.100 445.950 220.200 448.050 ;
        RECT 238.950 445.950 241.050 448.050 ;
        RECT 241.950 445.950 244.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 295.950 445.950 298.050 448.050 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 535.950 445.950 538.050 448.050 ;
        RECT 538.950 445.950 541.050 448.050 ;
        RECT 541.950 445.950 544.050 448.050 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 562.950 445.950 565.050 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 679.950 445.950 682.050 448.950 ;
        RECT 689.700 448.050 690.900 461.400 ;
        RECT 710.100 455.400 711.900 467.400 ;
        RECT 713.100 456.300 714.900 467.400 ;
        RECT 716.100 457.200 717.900 468.000 ;
        RECT 719.100 456.300 720.900 467.400 ;
        RECT 722.700 461.400 724.500 468.000 ;
        RECT 725.700 461.400 727.500 467.400 ;
        RECT 729.000 461.400 730.800 468.000 ;
        RECT 732.000 461.400 733.800 467.400 ;
        RECT 735.000 461.400 736.800 468.000 ;
        RECT 738.000 461.400 739.800 467.400 ;
        RECT 741.000 461.400 742.800 468.000 ;
        RECT 744.000 464.400 745.800 467.400 ;
        RECT 747.000 464.400 748.800 467.400 ;
        RECT 750.000 464.400 751.800 467.400 ;
        RECT 743.700 462.300 745.800 464.400 ;
        RECT 746.700 462.300 748.800 464.400 ;
        RECT 749.700 462.300 751.800 464.400 ;
        RECT 753.000 461.400 754.800 467.400 ;
        RECT 756.000 461.400 757.800 468.000 ;
        RECT 713.100 455.400 720.900 456.300 ;
        RECT 705.000 450.450 709.050 451.050 ;
        RECT 704.550 448.950 709.050 450.450 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 89.100 435.600 90.300 445.950 ;
        RECT 108.000 442.200 108.900 445.950 ;
        RECT 110.100 444.150 111.900 445.950 ;
        RECT 116.100 444.150 117.900 445.950 ;
        RECT 108.000 441.000 111.300 442.200 ;
        RECT 64.500 432.600 66.300 435.600 ;
        RECT 67.500 432.000 69.300 435.600 ;
        RECT 86.100 432.000 87.900 435.600 ;
        RECT 89.100 432.600 90.900 435.600 ;
        RECT 109.500 432.600 111.300 441.000 ;
        RECT 116.100 432.000 117.900 441.600 ;
        RECT 137.700 435.600 138.600 445.950 ;
        RECT 158.100 444.150 159.900 445.950 ;
        RECT 161.100 441.600 162.300 445.950 ;
        RECT 164.100 444.150 165.900 445.950 ;
        RECT 185.250 444.150 187.050 445.950 ;
        RECT 158.700 440.700 162.300 441.600 ;
        RECT 188.100 440.700 189.300 445.950 ;
        RECT 191.100 444.150 192.900 445.950 ;
        RECT 218.100 440.700 219.300 445.950 ;
        RECT 242.100 444.150 243.900 445.950 ;
        RECT 245.700 441.600 246.900 445.950 ;
        RECT 248.100 444.150 249.900 445.950 ;
        RECT 245.700 440.700 249.300 441.600 ;
        RECT 158.700 438.600 159.900 440.700 ;
        RECT 188.100 439.800 192.300 440.700 ;
        RECT 134.100 432.000 135.900 435.600 ;
        RECT 137.100 432.600 138.900 435.600 ;
        RECT 140.100 432.000 141.900 435.600 ;
        RECT 158.100 432.600 159.900 438.600 ;
        RECT 161.100 437.700 168.900 439.050 ;
        RECT 161.100 432.600 162.900 437.700 ;
        RECT 164.100 432.000 165.900 436.800 ;
        RECT 167.100 432.600 168.900 437.700 ;
        RECT 185.400 432.000 187.200 438.600 ;
        RECT 190.500 432.600 192.300 439.800 ;
        RECT 212.100 439.500 219.300 440.700 ;
        RECT 212.100 438.600 213.300 439.500 ;
        RECT 218.100 438.600 219.300 439.500 ;
        RECT 209.100 432.000 210.900 438.600 ;
        RECT 212.100 432.600 213.900 438.600 ;
        RECT 215.100 432.000 216.900 438.600 ;
        RECT 218.100 432.600 219.900 438.600 ;
        RECT 221.100 432.000 222.900 438.600 ;
        RECT 239.100 437.700 246.900 439.050 ;
        RECT 239.100 432.600 240.900 437.700 ;
        RECT 242.100 432.000 243.900 436.800 ;
        RECT 245.100 432.600 246.900 437.700 ;
        RECT 248.100 438.600 249.300 440.700 ;
        RECT 248.100 432.600 249.900 438.600 ;
        RECT 269.400 435.600 270.300 445.950 ;
        RECT 277.950 441.450 280.050 442.050 ;
        RECT 289.950 441.450 292.050 442.050 ;
        RECT 277.950 440.550 292.050 441.450 ;
        RECT 277.950 439.950 280.050 440.550 ;
        RECT 289.950 439.950 292.050 440.550 ;
        RECT 293.400 435.600 294.300 445.950 ;
        RECT 317.700 435.600 318.600 445.950 ;
        RECT 341.100 435.600 342.300 445.950 ;
        RECT 359.100 444.150 360.900 445.950 ;
        RECT 362.700 440.700 363.900 445.950 ;
        RECT 364.950 444.150 366.750 445.950 ;
        RECT 383.100 444.150 384.900 445.950 ;
        RECT 389.100 444.150 390.900 445.950 ;
        RECT 392.100 442.200 393.000 445.950 ;
        RECT 410.250 444.150 412.050 445.950 ;
        RECT 359.700 439.800 363.900 440.700 ;
        RECT 266.100 432.000 267.900 435.600 ;
        RECT 269.100 432.600 270.900 435.600 ;
        RECT 272.100 432.000 273.900 435.600 ;
        RECT 290.100 432.000 291.900 435.600 ;
        RECT 293.100 432.600 294.900 435.600 ;
        RECT 296.100 432.000 297.900 435.600 ;
        RECT 314.100 432.000 315.900 435.600 ;
        RECT 317.100 432.600 318.900 435.600 ;
        RECT 320.100 432.000 321.900 435.600 ;
        RECT 338.100 432.000 339.900 435.600 ;
        RECT 341.100 432.600 342.900 435.600 ;
        RECT 359.700 432.600 361.500 439.800 ;
        RECT 364.800 432.000 366.600 438.600 ;
        RECT 383.100 432.000 384.900 441.600 ;
        RECT 389.700 441.000 393.000 442.200 ;
        RECT 389.700 432.600 391.500 441.000 ;
        RECT 413.100 440.700 414.300 445.950 ;
        RECT 416.100 444.150 417.900 445.950 ;
        RECT 413.100 439.800 417.300 440.700 ;
        RECT 410.400 432.000 412.200 438.600 ;
        RECT 415.500 432.600 417.300 439.800 ;
        RECT 437.700 435.600 438.600 445.950 ;
        RECT 461.100 444.150 462.900 445.950 ;
        RECT 464.700 441.600 465.900 445.950 ;
        RECT 467.100 444.150 468.900 445.950 ;
        RECT 485.100 444.150 486.900 445.950 ;
        RECT 464.700 440.700 468.300 441.600 ;
        RECT 458.100 437.700 465.900 439.050 ;
        RECT 434.100 432.000 435.900 435.600 ;
        RECT 437.100 432.600 438.900 435.600 ;
        RECT 440.100 432.000 441.900 435.600 ;
        RECT 458.100 432.600 459.900 437.700 ;
        RECT 461.100 432.000 462.900 436.800 ;
        RECT 464.100 432.600 465.900 437.700 ;
        RECT 467.100 438.600 468.300 440.700 ;
        RECT 472.950 441.450 475.050 442.050 ;
        RECT 481.950 441.450 484.050 442.050 ;
        RECT 472.950 440.550 484.050 441.450 ;
        RECT 488.700 440.700 489.900 445.950 ;
        RECT 490.950 444.150 492.750 445.950 ;
        RECT 509.100 444.150 510.900 445.950 ;
        RECT 512.700 440.700 513.900 445.950 ;
        RECT 514.950 444.150 516.750 445.950 ;
        RECT 533.100 444.150 534.900 445.950 ;
        RECT 539.100 444.150 540.900 445.950 ;
        RECT 542.100 442.200 543.000 445.950 ;
        RECT 560.100 444.150 561.900 445.950 ;
        RECT 472.950 439.950 475.050 440.550 ;
        RECT 481.950 439.950 484.050 440.550 ;
        RECT 485.700 439.800 489.900 440.700 ;
        RECT 509.700 439.800 513.900 440.700 ;
        RECT 467.100 432.600 468.900 438.600 ;
        RECT 485.700 432.600 487.500 439.800 ;
        RECT 490.800 432.000 492.600 438.600 ;
        RECT 509.700 432.600 511.500 439.800 ;
        RECT 514.800 432.000 516.600 438.600 ;
        RECT 533.100 432.000 534.900 441.600 ;
        RECT 539.700 441.000 543.000 442.200 ;
        RECT 563.100 441.600 564.300 445.950 ;
        RECT 566.100 444.150 567.900 445.950 ;
        RECT 539.700 432.600 541.500 441.000 ;
        RECT 560.700 440.700 564.300 441.600 ;
        RECT 574.950 441.450 577.050 442.050 ;
        RECT 586.950 441.450 589.050 441.750 ;
        RECT 560.700 438.600 561.900 440.700 ;
        RECT 574.950 440.550 589.050 441.450 ;
        RECT 574.950 439.950 577.050 440.550 ;
        RECT 586.950 439.650 589.050 440.550 ;
        RECT 560.100 432.600 561.900 438.600 ;
        RECT 563.100 437.700 570.900 439.050 ;
        RECT 563.100 432.600 564.900 437.700 ;
        RECT 566.100 432.000 567.900 436.800 ;
        RECT 569.100 432.600 570.900 437.700 ;
        RECT 590.400 435.600 591.300 445.950 ;
        RECT 611.100 444.150 612.900 445.950 ;
        RECT 614.100 441.600 615.300 445.950 ;
        RECT 617.100 444.150 618.900 445.950 ;
        RECT 611.700 440.700 615.300 441.600 ;
        RECT 611.700 438.600 612.900 440.700 ;
        RECT 587.100 432.000 588.900 435.600 ;
        RECT 590.100 432.600 591.900 435.600 ;
        RECT 593.100 432.000 594.900 435.600 ;
        RECT 611.100 432.600 612.900 438.600 ;
        RECT 614.100 437.700 621.900 439.050 ;
        RECT 614.100 432.600 615.900 437.700 ;
        RECT 617.100 432.000 618.900 436.800 ;
        RECT 620.100 432.600 621.900 437.700 ;
        RECT 641.100 435.600 642.300 445.950 ;
        RECT 659.100 444.150 660.900 445.950 ;
        RECT 665.250 444.150 667.050 445.950 ;
        RECT 668.700 438.600 669.600 445.950 ;
        RECT 686.100 444.150 687.900 445.950 ;
        RECT 689.700 440.700 690.900 445.950 ;
        RECT 691.950 444.150 693.750 445.950 ;
        RECT 704.550 442.050 705.450 448.950 ;
        RECT 710.400 448.050 711.300 455.400 ;
        RECT 726.000 451.050 727.500 461.400 ;
        RECT 732.000 460.500 733.200 461.400 ;
        RECT 715.950 448.050 717.750 449.850 ;
        RECT 725.100 448.950 727.500 451.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 712.950 445.950 715.050 448.050 ;
        RECT 715.950 445.950 718.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 638.100 432.000 639.900 435.600 ;
        RECT 641.100 432.600 642.900 435.600 ;
        RECT 660.000 432.000 661.800 438.600 ;
        RECT 664.500 437.400 669.600 438.600 ;
        RECT 686.700 439.800 690.900 440.700 ;
        RECT 703.950 439.950 706.050 442.050 ;
        RECT 664.500 432.600 666.300 437.400 ;
        RECT 667.500 432.000 669.300 435.600 ;
        RECT 686.700 432.600 688.500 439.800 ;
        RECT 710.400 438.600 711.300 445.950 ;
        RECT 712.950 444.150 714.750 445.950 ;
        RECT 719.100 444.150 720.900 445.950 ;
        RECT 691.800 432.000 693.600 438.600 ;
        RECT 710.400 437.400 715.500 438.600 ;
        RECT 710.700 432.000 712.500 435.600 ;
        RECT 713.700 432.600 715.500 437.400 ;
        RECT 718.200 432.000 720.000 438.600 ;
        RECT 726.000 435.600 727.500 448.950 ;
        RECT 722.700 432.000 724.500 435.600 ;
        RECT 725.700 432.600 727.500 435.600 ;
        RECT 729.300 459.600 733.200 460.500 ;
        RECT 729.300 456.300 730.200 459.600 ;
        RECT 734.100 458.400 735.900 459.000 ;
        RECT 738.600 458.400 739.800 461.400 ;
        RECT 746.700 460.500 748.800 461.400 ;
        RECT 740.700 459.300 748.800 460.500 ;
        RECT 740.700 458.700 742.500 459.300 ;
        RECT 734.100 457.200 739.800 458.400 ;
        RECT 752.100 457.500 754.800 461.400 ;
        RECT 759.000 459.900 760.800 467.400 ;
        RECT 762.900 461.400 764.700 468.000 ;
        RECT 765.900 461.400 767.700 467.400 ;
        RECT 768.900 464.400 770.700 467.400 ;
        RECT 771.900 464.400 773.700 467.400 ;
        RECT 768.600 462.300 770.700 464.400 ;
        RECT 771.600 462.300 773.700 464.400 ;
        RECT 775.500 461.400 777.300 468.000 ;
        RECT 757.500 457.800 760.800 459.900 ;
        RECT 766.200 459.300 768.300 461.400 ;
        RECT 778.500 458.400 780.300 467.400 ;
        RECT 781.500 461.400 783.300 468.000 ;
        RECT 784.500 462.300 786.300 467.400 ;
        RECT 784.500 461.400 786.600 462.300 ;
        RECT 787.500 461.400 789.300 468.000 ;
        RECT 806.100 461.400 807.900 467.400 ;
        RECT 809.100 461.400 810.900 468.000 ;
        RECT 827.700 461.400 829.500 468.000 ;
        RECT 785.700 460.500 786.600 461.400 ;
        RECT 785.700 459.600 789.300 460.500 ;
        RECT 783.000 458.400 784.800 458.700 ;
        RECT 743.700 456.300 745.800 457.500 ;
        RECT 729.300 455.400 745.800 456.300 ;
        RECT 749.100 456.600 751.200 457.500 ;
        RECT 765.600 457.200 784.800 458.400 ;
        RECT 765.600 456.600 766.800 457.200 ;
        RECT 783.000 456.900 784.800 457.200 ;
        RECT 749.100 455.400 766.800 456.600 ;
        RECT 769.500 455.700 771.600 456.300 ;
        RECT 779.700 455.700 781.500 456.300 ;
        RECT 729.300 438.600 730.200 455.400 ;
        RECT 769.500 454.500 781.500 455.700 ;
        RECT 731.100 453.300 766.800 454.500 ;
        RECT 769.500 454.200 771.600 454.500 ;
        RECT 731.100 452.700 732.900 453.300 ;
        RECT 765.600 452.700 766.800 453.300 ;
        RECT 734.100 448.950 736.200 451.050 ;
        RECT 734.700 446.100 736.200 448.950 ;
        RECT 738.300 448.800 743.400 450.600 ;
        RECT 742.500 447.300 743.400 448.800 ;
        RECT 746.100 450.300 747.900 452.100 ;
        RECT 752.100 451.800 754.200 452.100 ;
        RECT 765.600 451.800 779.100 452.700 ;
        RECT 746.100 449.100 747.000 450.300 ;
        RECT 752.100 450.000 756.000 451.800 ;
        RECT 757.500 450.300 759.600 451.200 ;
        RECT 777.300 451.050 779.100 451.800 ;
        RECT 757.500 449.100 768.600 450.300 ;
        RECT 777.300 449.250 781.200 451.050 ;
        RECT 746.100 448.200 759.600 449.100 ;
        RECT 766.800 448.500 768.600 449.100 ;
        RECT 779.100 448.950 781.200 449.250 ;
        RECT 785.100 448.950 787.200 451.050 ;
        RECT 785.100 447.300 786.900 448.950 ;
        RECT 742.500 446.100 786.900 447.300 ;
        RECT 734.700 444.600 741.300 446.100 ;
        RECT 731.100 441.900 738.900 443.700 ;
        RECT 739.800 443.100 756.900 444.600 ;
        RECT 754.800 442.500 756.900 443.100 ;
        RECT 761.100 444.000 763.200 445.050 ;
        RECT 761.100 443.100 766.200 444.000 ;
        RECT 769.800 443.400 771.600 445.200 ;
        RECT 788.100 443.400 789.300 459.600 ;
        RECT 802.950 450.450 805.050 451.050 ;
        RECT 791.550 449.550 805.050 450.450 ;
        RECT 791.550 444.900 792.450 449.550 ;
        RECT 802.950 448.950 805.050 449.550 ;
        RECT 806.700 448.050 807.900 461.400 ;
        RECT 808.950 459.450 811.050 460.050 ;
        RECT 820.950 459.450 823.050 460.050 ;
        RECT 808.950 458.550 823.050 459.450 ;
        RECT 808.950 457.950 811.050 458.550 ;
        RECT 820.950 457.950 823.050 458.550 ;
        RECT 828.000 458.100 829.800 459.900 ;
        RECT 830.700 456.900 832.500 467.400 ;
        RECT 830.100 455.400 832.500 456.900 ;
        RECT 835.800 455.400 837.600 468.000 ;
        RECT 854.100 461.400 855.900 467.400 ;
        RECT 811.950 450.450 816.000 451.050 ;
        RECT 809.100 448.050 810.900 449.850 ;
        RECT 811.950 448.950 816.450 450.450 ;
        RECT 805.950 445.950 808.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 761.100 442.950 763.200 443.100 ;
        RECT 737.400 438.600 738.900 441.900 ;
        RECT 755.100 440.700 756.900 442.500 ;
        RECT 764.400 442.200 766.200 443.100 ;
        RECT 770.700 440.400 771.600 443.400 ;
        RECT 772.500 442.200 789.300 443.400 ;
        RECT 790.950 442.800 793.050 444.900 ;
        RECT 772.500 441.300 774.600 442.200 ;
        RECT 783.300 440.700 785.100 441.300 ;
        RECT 743.100 438.600 749.700 440.400 ;
        RECT 764.400 439.200 771.600 440.400 ;
        RECT 776.700 439.500 785.100 440.700 ;
        RECT 764.400 438.600 765.300 439.200 ;
        RECT 767.400 438.600 769.200 439.200 ;
        RECT 776.700 438.600 778.200 439.500 ;
        RECT 788.100 438.600 789.300 442.200 ;
        RECT 729.300 432.600 731.100 438.600 ;
        RECT 734.700 432.000 736.500 438.600 ;
        RECT 737.400 437.400 741.600 438.600 ;
        RECT 739.800 432.600 741.600 437.400 ;
        RECT 743.700 435.600 745.800 437.700 ;
        RECT 746.700 435.600 748.800 437.700 ;
        RECT 749.700 435.600 751.800 437.700 ;
        RECT 752.700 435.600 754.800 437.700 ;
        RECT 758.100 436.500 760.800 438.600 ;
        RECT 762.600 437.400 765.300 438.600 ;
        RECT 762.600 436.500 764.400 437.400 ;
        RECT 744.000 432.600 745.800 435.600 ;
        RECT 747.000 432.600 748.800 435.600 ;
        RECT 750.000 432.600 751.800 435.600 ;
        RECT 753.000 432.600 754.800 435.600 ;
        RECT 756.000 432.000 757.800 435.600 ;
        RECT 759.000 432.600 760.800 436.500 ;
        RECT 766.200 435.600 768.300 437.700 ;
        RECT 769.200 435.600 771.300 437.700 ;
        RECT 772.200 435.600 774.300 437.700 ;
        RECT 763.500 432.000 765.300 435.600 ;
        RECT 766.500 432.600 768.300 435.600 ;
        RECT 769.500 432.600 771.300 435.600 ;
        RECT 772.500 432.600 774.300 435.600 ;
        RECT 776.700 432.600 778.500 438.600 ;
        RECT 782.100 432.000 783.900 438.600 ;
        RECT 787.500 432.600 789.300 438.600 ;
        RECT 806.700 435.600 807.900 445.950 ;
        RECT 815.550 441.900 816.450 448.950 ;
        RECT 830.100 448.050 831.300 455.400 ;
        RECT 854.100 454.500 855.300 461.400 ;
        RECT 857.100 457.200 858.900 468.000 ;
        RECT 860.100 455.400 861.900 467.400 ;
        RECT 863.700 461.400 865.500 468.000 ;
        RECT 866.700 462.300 868.500 467.400 ;
        RECT 866.400 461.400 868.500 462.300 ;
        RECT 869.700 461.400 871.500 468.000 ;
        RECT 866.400 460.500 867.300 461.400 ;
        RECT 854.100 453.600 859.800 454.500 ;
        RECT 858.000 452.700 859.800 453.600 ;
        RECT 838.950 450.450 843.000 451.050 ;
        RECT 836.100 448.050 837.900 449.850 ;
        RECT 838.950 448.950 843.450 450.450 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 827.100 444.150 828.900 445.950 ;
        RECT 814.950 439.800 817.050 441.900 ;
        RECT 830.100 441.600 831.300 445.950 ;
        RECT 833.100 444.150 834.900 445.950 ;
        RECT 842.550 445.050 843.450 448.950 ;
        RECT 854.400 448.050 856.200 449.850 ;
        RECT 854.400 445.950 856.500 448.050 ;
        RECT 838.950 443.550 843.450 445.050 ;
        RECT 838.950 442.950 843.000 443.550 ;
        RECT 827.700 440.700 831.300 441.600 ;
        RECT 858.000 441.300 858.900 452.700 ;
        RECT 860.700 448.050 861.900 455.400 ;
        RECT 859.800 445.950 861.900 448.050 ;
        RECT 827.700 438.600 828.900 440.700 ;
        RECT 858.000 440.400 859.800 441.300 ;
        RECT 854.100 439.500 859.800 440.400 ;
        RECT 806.100 432.600 807.900 435.600 ;
        RECT 809.100 432.000 810.900 435.600 ;
        RECT 827.100 432.600 828.900 438.600 ;
        RECT 830.100 437.700 837.900 439.050 ;
        RECT 830.100 432.600 831.900 437.700 ;
        RECT 833.100 432.000 834.900 436.800 ;
        RECT 836.100 432.600 837.900 437.700 ;
        RECT 854.100 435.600 855.300 439.500 ;
        RECT 860.700 438.600 861.900 445.950 ;
        RECT 854.100 432.600 855.900 435.600 ;
        RECT 857.100 432.000 858.900 438.600 ;
        RECT 860.100 432.600 861.900 438.600 ;
        RECT 863.700 459.600 867.300 460.500 ;
        RECT 863.700 443.400 864.900 459.600 ;
        RECT 868.200 458.400 870.000 458.700 ;
        RECT 872.700 458.400 874.500 467.400 ;
        RECT 875.700 461.400 877.500 468.000 ;
        RECT 879.300 464.400 881.100 467.400 ;
        RECT 882.300 464.400 884.100 467.400 ;
        RECT 879.300 462.300 881.400 464.400 ;
        RECT 882.300 462.300 884.400 464.400 ;
        RECT 885.300 461.400 887.100 467.400 ;
        RECT 888.300 461.400 890.100 468.000 ;
        RECT 884.700 459.300 886.800 461.400 ;
        RECT 892.200 459.900 894.000 467.400 ;
        RECT 895.200 461.400 897.000 468.000 ;
        RECT 898.200 461.400 900.000 467.400 ;
        RECT 901.200 464.400 903.000 467.400 ;
        RECT 904.200 464.400 906.000 467.400 ;
        RECT 907.200 464.400 909.000 467.400 ;
        RECT 901.200 462.300 903.300 464.400 ;
        RECT 904.200 462.300 906.300 464.400 ;
        RECT 907.200 462.300 909.300 464.400 ;
        RECT 910.200 461.400 912.000 468.000 ;
        RECT 913.200 461.400 915.000 467.400 ;
        RECT 916.200 461.400 918.000 468.000 ;
        RECT 919.200 461.400 921.000 467.400 ;
        RECT 922.200 461.400 924.000 468.000 ;
        RECT 925.500 461.400 927.300 467.400 ;
        RECT 928.500 461.400 930.300 468.000 ;
        RECT 868.200 457.200 887.400 458.400 ;
        RECT 892.200 457.800 895.500 459.900 ;
        RECT 898.200 457.500 900.900 461.400 ;
        RECT 904.200 460.500 906.300 461.400 ;
        RECT 904.200 459.300 912.300 460.500 ;
        RECT 910.500 458.700 912.300 459.300 ;
        RECT 913.200 458.400 914.400 461.400 ;
        RECT 919.800 460.500 921.000 461.400 ;
        RECT 919.800 459.600 923.700 460.500 ;
        RECT 917.100 458.400 918.900 459.000 ;
        RECT 868.200 456.900 870.000 457.200 ;
        RECT 886.200 456.600 887.400 457.200 ;
        RECT 901.800 456.600 903.900 457.500 ;
        RECT 871.500 455.700 873.300 456.300 ;
        RECT 881.400 455.700 883.500 456.300 ;
        RECT 871.500 454.500 883.500 455.700 ;
        RECT 886.200 455.400 903.900 456.600 ;
        RECT 907.200 456.300 909.300 457.500 ;
        RECT 913.200 457.200 918.900 458.400 ;
        RECT 922.800 456.300 923.700 459.600 ;
        RECT 907.200 455.400 923.700 456.300 ;
        RECT 881.400 454.200 883.500 454.500 ;
        RECT 886.200 453.300 921.900 454.500 ;
        RECT 886.200 452.700 887.400 453.300 ;
        RECT 920.100 452.700 921.900 453.300 ;
        RECT 873.900 451.800 887.400 452.700 ;
        RECT 898.800 451.800 900.900 452.100 ;
        RECT 873.900 451.050 875.700 451.800 ;
        RECT 865.800 448.950 867.900 451.050 ;
        RECT 871.800 449.250 875.700 451.050 ;
        RECT 893.400 450.300 895.500 451.200 ;
        RECT 871.800 448.950 873.900 449.250 ;
        RECT 884.400 449.100 895.500 450.300 ;
        RECT 897.000 450.000 900.900 451.800 ;
        RECT 905.100 450.300 906.900 452.100 ;
        RECT 906.000 449.100 906.900 450.300 ;
        RECT 866.100 447.300 867.900 448.950 ;
        RECT 884.400 448.500 886.200 449.100 ;
        RECT 893.400 448.200 906.900 449.100 ;
        RECT 909.600 448.800 914.700 450.600 ;
        RECT 916.800 448.950 918.900 451.050 ;
        RECT 909.600 447.300 910.500 448.800 ;
        RECT 866.100 446.100 910.500 447.300 ;
        RECT 916.800 446.100 918.300 448.950 ;
        RECT 881.400 443.400 883.200 445.200 ;
        RECT 889.800 444.000 891.900 445.050 ;
        RECT 911.700 444.600 918.300 446.100 ;
        RECT 863.700 442.200 880.500 443.400 ;
        RECT 863.700 438.600 864.900 442.200 ;
        RECT 878.400 441.300 880.500 442.200 ;
        RECT 867.900 440.700 869.700 441.300 ;
        RECT 867.900 439.500 876.300 440.700 ;
        RECT 874.800 438.600 876.300 439.500 ;
        RECT 881.400 440.400 882.300 443.400 ;
        RECT 886.800 443.100 891.900 444.000 ;
        RECT 886.800 442.200 888.600 443.100 ;
        RECT 889.800 442.950 891.900 443.100 ;
        RECT 896.100 443.100 913.200 444.600 ;
        RECT 896.100 442.500 898.200 443.100 ;
        RECT 896.100 440.700 897.900 442.500 ;
        RECT 914.100 441.900 921.900 443.700 ;
        RECT 881.400 439.200 888.600 440.400 ;
        RECT 883.800 438.600 885.600 439.200 ;
        RECT 887.700 438.600 888.600 439.200 ;
        RECT 903.300 438.600 909.900 440.400 ;
        RECT 914.100 438.600 915.600 441.900 ;
        RECT 922.800 438.600 923.700 455.400 ;
        RECT 863.700 432.600 865.500 438.600 ;
        RECT 869.100 432.000 870.900 438.600 ;
        RECT 874.500 432.600 876.300 438.600 ;
        RECT 878.700 435.600 880.800 437.700 ;
        RECT 881.700 435.600 883.800 437.700 ;
        RECT 884.700 435.600 886.800 437.700 ;
        RECT 887.700 437.400 890.400 438.600 ;
        RECT 888.600 436.500 890.400 437.400 ;
        RECT 892.200 436.500 894.900 438.600 ;
        RECT 878.700 432.600 880.500 435.600 ;
        RECT 881.700 432.600 883.500 435.600 ;
        RECT 884.700 432.600 886.500 435.600 ;
        RECT 887.700 432.000 889.500 435.600 ;
        RECT 892.200 432.600 894.000 436.500 ;
        RECT 898.200 435.600 900.300 437.700 ;
        RECT 901.200 435.600 903.300 437.700 ;
        RECT 904.200 435.600 906.300 437.700 ;
        RECT 907.200 435.600 909.300 437.700 ;
        RECT 911.400 437.400 915.600 438.600 ;
        RECT 895.200 432.000 897.000 435.600 ;
        RECT 898.200 432.600 900.000 435.600 ;
        RECT 901.200 432.600 903.000 435.600 ;
        RECT 904.200 432.600 906.000 435.600 ;
        RECT 907.200 432.600 909.000 435.600 ;
        RECT 911.400 432.600 913.200 437.400 ;
        RECT 916.500 432.000 918.300 438.600 ;
        RECT 921.900 432.600 923.700 438.600 ;
        RECT 925.500 451.050 927.000 461.400 ;
        RECT 947.100 456.600 948.900 467.400 ;
        RECT 950.100 457.500 951.900 468.000 ;
        RECT 947.100 455.400 951.900 456.600 ;
        RECT 949.800 454.500 951.900 455.400 ;
        RECT 954.600 455.400 956.400 467.400 ;
        RECT 959.100 457.500 960.900 468.000 ;
        RECT 962.100 456.300 963.900 467.400 ;
        RECT 959.400 455.400 963.900 456.300 ;
        RECT 980.100 456.600 981.900 467.400 ;
        RECT 983.100 457.500 984.900 468.000 ;
        RECT 980.100 455.400 984.900 456.600 ;
        RECT 954.600 454.050 955.800 455.400 ;
        RECT 954.300 453.000 955.800 454.050 ;
        RECT 959.400 453.300 961.500 455.400 ;
        RECT 982.800 454.500 984.900 455.400 ;
        RECT 987.600 455.400 989.400 467.400 ;
        RECT 992.100 457.500 993.900 468.000 ;
        RECT 995.100 456.300 996.900 467.400 ;
        RECT 1013.700 461.400 1015.500 468.000 ;
        RECT 1014.000 458.100 1015.800 459.900 ;
        RECT 1016.700 456.900 1018.500 467.400 ;
        RECT 992.400 455.400 996.900 456.300 ;
        RECT 1016.100 455.400 1018.500 456.900 ;
        RECT 1021.800 455.400 1023.600 468.000 ;
        RECT 1024.950 462.450 1027.050 463.050 ;
        RECT 1036.950 462.450 1039.050 463.050 ;
        RECT 1024.950 461.550 1039.050 462.450 ;
        RECT 1024.950 460.950 1027.050 461.550 ;
        RECT 1036.950 460.950 1039.050 461.550 ;
        RECT 987.600 454.050 988.800 455.400 ;
        RECT 987.300 453.000 988.800 454.050 ;
        RECT 992.400 453.300 994.500 455.400 ;
        RECT 954.300 451.050 955.200 453.000 ;
        RECT 925.500 448.950 927.900 451.050 ;
        RECT 925.500 435.600 927.000 448.950 ;
        RECT 947.400 448.050 949.200 449.850 ;
        RECT 953.100 448.950 955.200 451.050 ;
        RECT 956.100 451.500 958.200 451.800 ;
        RECT 956.100 449.700 960.000 451.500 ;
        RECT 987.300 451.050 988.200 453.000 ;
        RECT 947.100 445.950 949.200 448.050 ;
        RECT 953.700 448.800 955.200 448.950 ;
        RECT 953.700 447.900 956.100 448.800 ;
        RECT 951.900 445.200 953.700 447.000 ;
        RECT 951.900 443.100 954.000 445.200 ;
        RECT 954.900 442.200 956.100 447.900 ;
        RECT 957.000 448.050 958.800 448.500 ;
        RECT 980.400 448.050 982.200 449.850 ;
        RECT 986.100 448.950 988.200 451.050 ;
        RECT 989.100 451.500 991.200 451.800 ;
        RECT 989.100 449.700 993.000 451.500 ;
        RECT 957.000 446.700 963.900 448.050 ;
        RECT 961.800 445.950 963.900 446.700 ;
        RECT 980.100 445.950 982.200 448.050 ;
        RECT 986.700 448.800 988.200 448.950 ;
        RECT 986.700 447.900 989.100 448.800 ;
        RECT 949.800 439.500 951.900 440.700 ;
        RECT 953.100 440.100 956.100 442.200 ;
        RECT 957.000 443.400 958.800 445.200 ;
        RECT 961.800 444.150 963.600 445.950 ;
        RECT 984.900 445.200 986.700 447.000 ;
        RECT 957.000 441.300 959.100 443.400 ;
        RECT 984.900 443.100 987.000 445.200 ;
        RECT 987.900 442.200 989.100 447.900 ;
        RECT 990.000 448.050 991.800 448.500 ;
        RECT 1016.100 448.050 1017.300 455.400 ;
        RECT 1018.950 453.450 1021.050 454.050 ;
        RECT 1036.950 453.450 1039.050 454.050 ;
        RECT 1018.950 452.550 1039.050 453.450 ;
        RECT 1018.950 451.950 1021.050 452.550 ;
        RECT 1036.950 451.950 1039.050 452.550 ;
        RECT 1024.950 450.450 1029.000 451.050 ;
        RECT 1022.100 448.050 1023.900 449.850 ;
        RECT 1024.950 448.950 1029.450 450.450 ;
        RECT 990.000 446.700 996.900 448.050 ;
        RECT 994.800 445.950 996.900 446.700 ;
        RECT 1012.950 445.950 1015.050 448.050 ;
        RECT 1015.950 445.950 1018.050 448.050 ;
        RECT 1018.950 445.950 1021.050 448.050 ;
        RECT 1021.950 445.950 1024.050 448.050 ;
        RECT 957.000 440.400 963.300 441.300 ;
        RECT 947.100 438.600 951.900 439.500 ;
        RECT 954.900 438.600 956.100 440.100 ;
        RECT 962.100 438.600 963.300 440.400 ;
        RECT 982.800 439.500 984.900 440.700 ;
        RECT 986.100 440.100 989.100 442.200 ;
        RECT 990.000 443.400 991.800 445.200 ;
        RECT 994.800 444.150 996.600 445.950 ;
        RECT 1013.100 444.150 1014.900 445.950 ;
        RECT 990.000 441.300 992.100 443.400 ;
        RECT 1016.100 441.600 1017.300 445.950 ;
        RECT 1019.100 444.150 1020.900 445.950 ;
        RECT 1028.550 445.050 1029.450 448.950 ;
        RECT 1024.950 443.550 1029.450 445.050 ;
        RECT 1024.950 442.950 1029.000 443.550 ;
        RECT 990.000 440.400 996.300 441.300 ;
        RECT 980.100 438.600 984.900 439.500 ;
        RECT 987.900 438.600 989.100 440.100 ;
        RECT 995.100 438.600 996.300 440.400 ;
        RECT 1013.700 440.700 1017.300 441.600 ;
        RECT 1013.700 438.600 1014.900 440.700 ;
        RECT 925.500 432.600 927.300 435.600 ;
        RECT 928.500 432.000 930.300 435.600 ;
        RECT 947.100 432.600 948.900 438.600 ;
        RECT 950.100 432.000 951.900 437.700 ;
        RECT 954.600 432.600 956.400 438.600 ;
        RECT 959.100 432.000 960.900 437.700 ;
        RECT 962.100 432.600 963.900 438.600 ;
        RECT 967.950 435.450 970.050 436.050 ;
        RECT 976.950 435.450 979.050 436.050 ;
        RECT 967.950 434.550 979.050 435.450 ;
        RECT 967.950 433.950 970.050 434.550 ;
        RECT 976.950 433.950 979.050 434.550 ;
        RECT 980.100 432.600 981.900 438.600 ;
        RECT 983.100 432.000 984.900 437.700 ;
        RECT 987.600 432.600 989.400 438.600 ;
        RECT 992.100 432.000 993.900 437.700 ;
        RECT 995.100 432.600 996.900 438.600 ;
        RECT 1013.100 432.600 1014.900 438.600 ;
        RECT 1016.100 437.700 1023.900 439.050 ;
        RECT 1016.100 432.600 1017.900 437.700 ;
        RECT 1019.100 432.000 1020.900 436.800 ;
        RECT 1022.100 432.600 1023.900 437.700 ;
        RECT 17.100 425.400 18.900 429.000 ;
        RECT 20.100 425.400 21.900 428.400 ;
        RECT 23.100 425.400 24.900 429.000 ;
        RECT 20.700 415.050 21.600 425.400 ;
        RECT 41.100 423.300 42.900 428.400 ;
        RECT 44.100 424.200 45.900 429.000 ;
        RECT 47.100 423.300 48.900 428.400 ;
        RECT 41.100 421.950 48.900 423.300 ;
        RECT 50.100 422.400 51.900 428.400 ;
        RECT 53.700 422.400 55.500 428.400 ;
        RECT 59.100 422.400 60.900 429.000 ;
        RECT 64.500 422.400 66.300 428.400 ;
        RECT 68.700 425.400 70.500 428.400 ;
        RECT 71.700 425.400 73.500 428.400 ;
        RECT 74.700 425.400 76.500 428.400 ;
        RECT 77.700 425.400 79.500 429.000 ;
        RECT 68.700 423.300 70.800 425.400 ;
        RECT 71.700 423.300 73.800 425.400 ;
        RECT 74.700 423.300 76.800 425.400 ;
        RECT 82.200 424.500 84.000 428.400 ;
        RECT 85.200 425.400 87.000 429.000 ;
        RECT 88.200 425.400 90.000 428.400 ;
        RECT 91.200 425.400 93.000 428.400 ;
        RECT 94.200 425.400 96.000 428.400 ;
        RECT 97.200 425.400 99.000 428.400 ;
        RECT 78.600 423.600 80.400 424.500 ;
        RECT 77.700 422.400 80.400 423.600 ;
        RECT 82.200 422.400 84.900 424.500 ;
        RECT 88.200 423.300 90.300 425.400 ;
        RECT 91.200 423.300 93.300 425.400 ;
        RECT 94.200 423.300 96.300 425.400 ;
        RECT 97.200 423.300 99.300 425.400 ;
        RECT 101.400 423.600 103.200 428.400 ;
        RECT 101.400 422.400 105.600 423.600 ;
        RECT 106.500 422.400 108.300 429.000 ;
        RECT 111.900 422.400 113.700 428.400 ;
        RECT 50.100 420.300 51.300 422.400 ;
        RECT 47.700 419.400 51.300 420.300 ;
        RECT 44.100 415.050 45.900 416.850 ;
        RECT 47.700 415.050 48.900 419.400 ;
        RECT 53.700 418.800 54.900 422.400 ;
        RECT 64.800 421.500 66.300 422.400 ;
        RECT 73.800 421.800 75.600 422.400 ;
        RECT 77.700 421.800 78.600 422.400 ;
        RECT 57.900 420.300 66.300 421.500 ;
        RECT 71.400 420.600 78.600 421.800 ;
        RECT 93.300 420.600 99.900 422.400 ;
        RECT 57.900 419.700 59.700 420.300 ;
        RECT 68.400 418.800 70.500 419.700 ;
        RECT 53.700 417.600 70.500 418.800 ;
        RECT 71.400 417.600 72.300 420.600 ;
        RECT 76.800 417.900 78.600 418.800 ;
        RECT 86.100 418.500 87.900 420.300 ;
        RECT 104.100 419.100 105.600 422.400 ;
        RECT 79.800 417.900 81.900 418.050 ;
        RECT 50.100 415.050 51.900 416.850 ;
        RECT 16.950 412.950 19.050 415.050 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 22.950 412.950 25.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 17.100 411.150 18.900 412.950 ;
        RECT 20.700 405.600 21.600 412.950 ;
        RECT 22.950 411.150 24.750 412.950 ;
        RECT 41.100 411.150 42.900 412.950 ;
        RECT 47.700 405.600 48.900 412.950 ;
        RECT 18.000 404.400 21.600 405.600 ;
        RECT 18.000 393.600 19.800 404.400 ;
        RECT 23.100 393.000 24.900 405.600 ;
        RECT 41.400 393.000 43.200 405.600 ;
        RECT 46.500 404.100 48.900 405.600 ;
        RECT 46.500 393.600 48.300 404.100 ;
        RECT 49.200 401.100 51.000 402.900 ;
        RECT 53.700 401.400 54.900 417.600 ;
        RECT 71.400 415.800 73.200 417.600 ;
        RECT 76.800 417.000 81.900 417.900 ;
        RECT 79.800 415.950 81.900 417.000 ;
        RECT 86.100 417.900 88.200 418.500 ;
        RECT 86.100 416.400 103.200 417.900 ;
        RECT 104.100 417.300 111.900 419.100 ;
        RECT 101.700 414.900 108.300 416.400 ;
        RECT 56.100 413.700 100.500 414.900 ;
        RECT 56.100 412.050 57.900 413.700 ;
        RECT 55.800 409.950 57.900 412.050 ;
        RECT 61.800 411.750 63.900 412.050 ;
        RECT 74.400 411.900 76.200 412.500 ;
        RECT 83.400 411.900 96.900 412.800 ;
        RECT 61.800 409.950 65.700 411.750 ;
        RECT 74.400 410.700 85.500 411.900 ;
        RECT 63.900 409.200 65.700 409.950 ;
        RECT 83.400 409.800 85.500 410.700 ;
        RECT 87.000 409.200 90.900 411.000 ;
        RECT 96.000 410.700 96.900 411.900 ;
        RECT 63.900 408.300 77.400 409.200 ;
        RECT 88.800 408.900 90.900 409.200 ;
        RECT 95.100 408.900 96.900 410.700 ;
        RECT 99.600 412.200 100.500 413.700 ;
        RECT 99.600 410.400 104.700 412.200 ;
        RECT 106.800 412.050 108.300 414.900 ;
        RECT 106.800 409.950 108.900 412.050 ;
        RECT 76.200 407.700 77.400 408.300 ;
        RECT 110.100 407.700 111.900 408.300 ;
        RECT 71.400 406.500 73.500 406.800 ;
        RECT 76.200 406.500 111.900 407.700 ;
        RECT 61.500 405.300 73.500 406.500 ;
        RECT 112.800 405.600 113.700 422.400 ;
        RECT 61.500 404.700 63.300 405.300 ;
        RECT 71.400 404.700 73.500 405.300 ;
        RECT 76.200 404.400 93.900 405.600 ;
        RECT 58.200 403.800 60.000 404.100 ;
        RECT 76.200 403.800 77.400 404.400 ;
        RECT 58.200 402.600 77.400 403.800 ;
        RECT 91.800 403.500 93.900 404.400 ;
        RECT 97.200 404.700 113.700 405.600 ;
        RECT 97.200 403.500 99.300 404.700 ;
        RECT 58.200 402.300 60.000 402.600 ;
        RECT 53.700 400.500 57.300 401.400 ;
        RECT 56.400 399.600 57.300 400.500 ;
        RECT 49.500 393.000 51.300 399.600 ;
        RECT 53.700 393.000 55.500 399.600 ;
        RECT 56.400 398.700 58.500 399.600 ;
        RECT 56.700 393.600 58.500 398.700 ;
        RECT 59.700 393.000 61.500 399.600 ;
        RECT 62.700 393.600 64.500 402.600 ;
        RECT 74.700 399.600 76.800 401.700 ;
        RECT 82.200 401.100 85.500 403.200 ;
        RECT 65.700 393.000 67.500 399.600 ;
        RECT 69.300 396.600 71.400 398.700 ;
        RECT 72.300 396.600 74.400 398.700 ;
        RECT 69.300 393.600 71.100 396.600 ;
        RECT 72.300 393.600 74.100 396.600 ;
        RECT 75.300 393.600 77.100 399.600 ;
        RECT 78.300 393.000 80.100 399.600 ;
        RECT 82.200 393.600 84.000 401.100 ;
        RECT 88.200 399.600 90.900 403.500 ;
        RECT 103.200 402.600 108.900 403.800 ;
        RECT 100.500 401.700 102.300 402.300 ;
        RECT 94.200 400.500 102.300 401.700 ;
        RECT 94.200 399.600 96.300 400.500 ;
        RECT 103.200 399.600 104.400 402.600 ;
        RECT 107.100 402.000 108.900 402.600 ;
        RECT 112.800 401.400 113.700 404.700 ;
        RECT 109.800 400.500 113.700 401.400 ;
        RECT 115.500 425.400 117.300 428.400 ;
        RECT 118.500 425.400 120.300 429.000 ;
        RECT 137.100 425.400 138.900 429.000 ;
        RECT 140.100 425.400 141.900 428.400 ;
        RECT 158.100 425.400 159.900 429.000 ;
        RECT 161.100 425.400 162.900 428.400 ;
        RECT 164.100 425.400 165.900 429.000 ;
        RECT 115.500 412.050 117.000 425.400 ;
        RECT 140.100 415.050 141.300 425.400 ;
        RECT 161.400 415.050 162.300 425.400 ;
        RECT 182.700 421.200 184.500 428.400 ;
        RECT 187.800 422.400 189.600 429.000 ;
        RECT 206.100 422.400 207.900 428.400 ;
        RECT 182.700 420.300 186.900 421.200 ;
        RECT 182.100 415.050 183.900 416.850 ;
        RECT 185.700 415.050 186.900 420.300 ;
        RECT 206.700 420.300 207.900 422.400 ;
        RECT 209.100 423.300 210.900 428.400 ;
        RECT 212.100 424.200 213.900 429.000 ;
        RECT 215.100 423.300 216.900 428.400 ;
        RECT 209.100 421.950 216.900 423.300 ;
        RECT 206.700 419.400 210.300 420.300 ;
        RECT 187.950 415.050 189.750 416.850 ;
        RECT 206.100 415.050 207.900 416.850 ;
        RECT 209.100 415.050 210.300 419.400 ;
        RECT 223.950 418.950 226.050 421.050 ;
        RECT 233.100 419.400 234.900 429.000 ;
        RECT 239.700 420.000 241.500 428.400 ;
        RECT 244.950 426.450 247.050 427.050 ;
        RECT 256.950 426.450 259.050 427.050 ;
        RECT 244.950 425.550 259.050 426.450 ;
        RECT 244.950 424.950 247.050 425.550 ;
        RECT 256.950 424.950 259.050 425.550 ;
        RECT 260.100 425.400 261.900 429.000 ;
        RECT 263.100 425.400 264.900 428.400 ;
        RECT 266.100 425.400 267.900 429.000 ;
        RECT 284.100 425.400 285.900 429.000 ;
        RECT 287.100 425.400 288.900 428.400 ;
        RECT 212.100 415.050 213.900 416.850 ;
        RECT 136.950 412.950 139.050 415.050 ;
        RECT 139.950 412.950 142.050 415.050 ;
        RECT 157.950 412.950 160.050 415.050 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 211.950 412.950 214.050 415.050 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 115.500 409.950 117.900 412.050 ;
        RECT 137.100 411.150 138.900 412.950 ;
        RECT 109.800 399.600 111.000 400.500 ;
        RECT 115.500 399.600 117.000 409.950 ;
        RECT 140.100 399.600 141.300 412.950 ;
        RECT 158.250 411.150 160.050 412.950 ;
        RECT 161.400 405.600 162.300 412.950 ;
        RECT 164.100 411.150 165.900 412.950 ;
        RECT 85.200 393.000 87.000 399.600 ;
        RECT 88.200 393.600 90.000 399.600 ;
        RECT 91.200 396.600 93.300 398.700 ;
        RECT 94.200 396.600 96.300 398.700 ;
        RECT 97.200 396.600 99.300 398.700 ;
        RECT 91.200 393.600 93.000 396.600 ;
        RECT 94.200 393.600 96.000 396.600 ;
        RECT 97.200 393.600 99.000 396.600 ;
        RECT 100.200 393.000 102.000 399.600 ;
        RECT 103.200 393.600 105.000 399.600 ;
        RECT 106.200 393.000 108.000 399.600 ;
        RECT 109.200 393.600 111.000 399.600 ;
        RECT 112.200 393.000 114.000 399.600 ;
        RECT 115.500 393.600 117.300 399.600 ;
        RECT 118.500 393.000 120.300 399.600 ;
        RECT 137.100 393.000 138.900 399.600 ;
        RECT 140.100 393.600 141.900 399.600 ;
        RECT 158.100 393.000 159.900 405.600 ;
        RECT 161.400 404.400 165.000 405.600 ;
        RECT 163.200 393.600 165.000 404.400 ;
        RECT 185.700 399.600 186.900 412.950 ;
        RECT 187.950 405.450 190.050 406.050 ;
        RECT 205.950 405.450 208.050 406.050 ;
        RECT 187.950 404.550 208.050 405.450 ;
        RECT 187.950 403.950 190.050 404.550 ;
        RECT 205.950 403.950 208.050 404.550 ;
        RECT 209.100 405.600 210.300 412.950 ;
        RECT 215.100 411.150 216.900 412.950 ;
        RECT 224.550 411.450 225.450 418.950 ;
        RECT 239.700 418.800 243.000 420.000 ;
        RECT 233.100 415.050 234.900 416.850 ;
        RECT 239.100 415.050 240.900 416.850 ;
        RECT 242.100 415.050 243.000 418.800 ;
        RECT 263.700 415.050 264.600 425.400 ;
        RECT 271.950 420.450 274.050 421.050 ;
        RECT 283.950 420.450 286.050 421.050 ;
        RECT 271.950 419.550 286.050 420.450 ;
        RECT 271.950 418.950 274.050 419.550 ;
        RECT 283.950 418.950 286.050 419.550 ;
        RECT 287.100 415.050 288.300 425.400 ;
        RECT 305.100 422.400 306.900 428.400 ;
        RECT 308.100 423.300 309.900 429.000 ;
        RECT 312.600 422.400 314.400 428.400 ;
        RECT 317.100 423.300 318.900 429.000 ;
        RECT 320.100 422.400 321.900 428.400 ;
        RECT 305.700 420.600 306.900 422.400 ;
        RECT 312.900 420.900 314.100 422.400 ;
        RECT 317.100 421.500 321.900 422.400 ;
        RECT 338.100 422.400 339.900 428.400 ;
        RECT 341.100 423.300 342.900 429.000 ;
        RECT 345.600 422.400 347.400 428.400 ;
        RECT 350.100 423.300 351.900 429.000 ;
        RECT 353.100 422.400 354.900 428.400 ;
        RECT 372.000 422.400 373.800 429.000 ;
        RECT 376.500 423.600 378.300 428.400 ;
        RECT 379.500 425.400 381.300 429.000 ;
        RECT 376.500 422.400 381.600 423.600 ;
        RECT 400.500 422.400 402.300 429.000 ;
        RECT 405.000 422.400 406.800 428.400 ;
        RECT 409.500 422.400 411.300 429.000 ;
        RECT 338.100 421.500 342.900 422.400 ;
        RECT 305.700 419.700 312.000 420.600 ;
        RECT 309.900 417.600 312.000 419.700 ;
        RECT 305.400 415.050 307.200 416.850 ;
        RECT 310.200 415.800 312.000 417.600 ;
        RECT 312.900 418.800 315.900 420.900 ;
        RECT 317.100 420.300 319.200 421.500 ;
        RECT 325.950 420.450 328.050 421.050 ;
        RECT 331.950 420.450 334.050 421.050 ;
        RECT 325.950 419.550 334.050 420.450 ;
        RECT 340.800 420.300 342.900 421.500 ;
        RECT 345.900 420.900 347.100 422.400 ;
        RECT 325.950 418.950 328.050 419.550 ;
        RECT 331.950 418.950 334.050 419.550 ;
        RECT 344.100 418.800 347.100 420.900 ;
        RECT 353.100 420.600 354.300 422.400 ;
        RECT 232.950 412.950 235.050 415.050 ;
        RECT 235.950 412.950 238.050 415.050 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 305.100 414.300 307.200 415.050 ;
        RECT 305.100 412.950 312.000 414.300 ;
        RECT 229.950 411.450 232.050 412.050 ;
        RECT 224.550 410.550 232.050 411.450 ;
        RECT 236.100 411.150 237.900 412.950 ;
        RECT 229.950 409.950 232.050 410.550 ;
        RECT 209.100 404.100 211.500 405.600 ;
        RECT 207.000 401.100 208.800 402.900 ;
        RECT 182.100 393.000 183.900 399.600 ;
        RECT 185.100 393.600 186.900 399.600 ;
        RECT 188.100 393.000 189.900 399.600 ;
        RECT 206.700 393.000 208.500 399.600 ;
        RECT 209.700 393.600 211.500 404.100 ;
        RECT 214.800 393.000 216.600 405.600 ;
        RECT 242.100 400.800 243.000 412.950 ;
        RECT 260.100 411.150 261.900 412.950 ;
        RECT 263.700 405.600 264.600 412.950 ;
        RECT 265.950 411.150 267.750 412.950 ;
        RECT 284.100 411.150 285.900 412.950 ;
        RECT 236.400 399.900 243.000 400.800 ;
        RECT 236.400 399.600 237.900 399.900 ;
        RECT 233.100 393.000 234.900 399.600 ;
        RECT 236.100 393.600 237.900 399.600 ;
        RECT 242.100 399.600 243.000 399.900 ;
        RECT 261.000 404.400 264.600 405.600 ;
        RECT 239.100 393.000 240.900 399.000 ;
        RECT 242.100 393.600 243.900 399.600 ;
        RECT 261.000 393.600 262.800 404.400 ;
        RECT 266.100 393.000 267.900 405.600 ;
        RECT 287.100 399.600 288.300 412.950 ;
        RECT 310.200 412.500 312.000 412.950 ;
        RECT 312.900 413.100 314.100 418.800 ;
        RECT 315.000 415.800 317.100 417.900 ;
        RECT 315.300 414.000 317.100 415.800 ;
        RECT 342.900 415.800 345.000 417.900 ;
        RECT 312.900 412.200 315.300 413.100 ;
        RECT 313.800 412.050 315.300 412.200 ;
        RECT 319.800 412.950 321.900 415.050 ;
        RECT 338.100 412.950 340.200 415.050 ;
        RECT 342.900 414.000 344.700 415.800 ;
        RECT 345.900 413.100 347.100 418.800 ;
        RECT 348.000 419.700 354.300 420.600 ;
        RECT 348.000 417.600 350.100 419.700 ;
        RECT 348.000 415.800 349.800 417.600 ;
        RECT 352.800 415.050 354.600 416.850 ;
        RECT 371.100 415.050 372.900 416.850 ;
        RECT 377.250 415.050 379.050 416.850 ;
        RECT 380.700 415.050 381.600 422.400 ;
        RECT 398.100 415.050 399.900 416.850 ;
        RECT 404.700 415.050 405.900 422.400 ;
        RECT 428.100 419.400 429.900 429.000 ;
        RECT 434.700 420.000 436.500 428.400 ;
        RECT 455.100 425.400 456.900 428.400 ;
        RECT 458.100 425.400 459.900 429.000 ;
        RECT 460.950 426.450 463.050 427.050 ;
        RECT 472.950 426.450 475.050 427.050 ;
        RECT 460.950 425.550 475.050 426.450 ;
        RECT 434.700 418.800 438.000 420.000 ;
        RECT 409.950 415.050 411.750 416.850 ;
        RECT 428.100 415.050 429.900 416.850 ;
        RECT 434.100 415.050 435.900 416.850 ;
        RECT 437.100 415.050 438.000 418.800 ;
        RECT 455.700 415.050 456.900 425.400 ;
        RECT 460.950 424.950 463.050 425.550 ;
        RECT 472.950 424.950 475.050 425.550 ;
        RECT 476.100 425.400 477.900 428.400 ;
        RECT 479.100 425.400 480.900 429.000 ;
        RECT 476.700 415.050 477.900 425.400 ;
        RECT 497.100 422.400 498.900 428.400 ;
        RECT 500.100 423.300 501.900 429.000 ;
        RECT 504.600 422.400 506.400 428.400 ;
        RECT 509.100 423.300 510.900 429.000 ;
        RECT 512.100 422.400 513.900 428.400 ;
        RECT 530.100 425.400 531.900 429.000 ;
        RECT 533.100 425.400 534.900 428.400 ;
        RECT 536.100 425.400 537.900 429.000 ;
        RECT 554.100 425.400 555.900 429.000 ;
        RECT 557.100 425.400 558.900 428.400 ;
        RECT 560.100 425.400 561.900 429.000 ;
        RECT 497.100 421.500 501.900 422.400 ;
        RECT 499.800 420.300 501.900 421.500 ;
        RECT 504.900 420.900 506.100 422.400 ;
        RECT 503.100 418.800 506.100 420.900 ;
        RECT 512.100 420.600 513.300 422.400 ;
        RECT 501.900 415.800 504.000 417.900 ;
        RECT 352.800 414.300 354.900 415.050 ;
        RECT 309.000 409.500 312.900 411.300 ;
        RECT 310.800 409.200 312.900 409.500 ;
        RECT 313.800 409.950 315.900 412.050 ;
        RECT 319.800 411.150 321.600 412.950 ;
        RECT 338.400 411.150 340.200 412.950 ;
        RECT 344.700 412.200 347.100 413.100 ;
        RECT 348.000 412.950 354.900 414.300 ;
        RECT 370.950 412.950 373.050 415.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 376.950 412.950 379.050 415.050 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 433.950 412.950 436.050 415.050 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 497.100 412.950 499.200 415.050 ;
        RECT 501.900 414.000 503.700 415.800 ;
        RECT 504.900 413.100 506.100 418.800 ;
        RECT 507.000 419.700 513.300 420.600 ;
        RECT 507.000 417.600 509.100 419.700 ;
        RECT 507.000 415.800 508.800 417.600 ;
        RECT 511.800 415.050 513.600 416.850 ;
        RECT 533.400 415.050 534.300 425.400 ;
        RECT 557.400 415.050 558.300 425.400 ;
        RECT 575.100 422.400 576.900 428.400 ;
        RECT 578.100 422.400 579.900 429.000 ;
        RECT 597.000 422.400 598.800 429.000 ;
        RECT 601.500 423.600 603.300 428.400 ;
        RECT 604.500 425.400 606.300 429.000 ;
        RECT 601.500 422.400 606.600 423.600 ;
        RECT 624.000 422.400 625.800 429.000 ;
        RECT 628.500 423.600 630.300 428.400 ;
        RECT 631.500 425.400 633.300 429.000 ;
        RECT 650.100 425.400 651.900 428.400 ;
        RECT 653.100 425.400 654.900 429.000 ;
        RECT 628.500 422.400 633.600 423.600 ;
        RECT 575.700 415.050 576.900 422.400 ;
        RECT 583.950 420.450 586.050 421.050 ;
        RECT 598.950 420.450 601.050 421.050 ;
        RECT 583.950 419.550 601.050 420.450 ;
        RECT 583.950 418.950 586.050 419.550 ;
        RECT 598.950 418.950 601.050 419.550 ;
        RECT 578.100 415.050 579.900 416.850 ;
        RECT 596.100 415.050 597.900 416.850 ;
        RECT 602.250 415.050 604.050 416.850 ;
        RECT 605.700 415.050 606.600 422.400 ;
        RECT 607.950 420.450 610.050 421.050 ;
        RECT 628.950 420.450 631.050 421.050 ;
        RECT 607.950 419.550 631.050 420.450 ;
        RECT 607.950 418.950 610.050 419.550 ;
        RECT 628.950 418.950 631.050 419.550 ;
        RECT 623.100 415.050 624.900 416.850 ;
        RECT 629.250 415.050 631.050 416.850 ;
        RECT 632.700 415.050 633.600 422.400 ;
        RECT 650.700 415.050 651.900 425.400 ;
        RECT 671.100 422.400 672.900 428.400 ;
        RECT 671.700 420.300 672.900 422.400 ;
        RECT 674.100 423.300 675.900 428.400 ;
        RECT 677.100 424.200 678.900 429.000 ;
        RECT 680.100 423.300 681.900 428.400 ;
        RECT 674.100 421.950 681.900 423.300 ;
        RECT 698.100 422.400 699.900 428.400 ;
        RECT 701.100 422.400 702.900 429.000 ;
        RECT 719.100 422.400 720.900 428.400 ;
        RECT 722.100 423.300 723.900 429.000 ;
        RECT 726.600 422.400 728.400 428.400 ;
        RECT 731.100 423.300 732.900 429.000 ;
        RECT 734.100 422.400 735.900 428.400 ;
        RECT 752.100 425.400 753.900 429.000 ;
        RECT 755.100 425.400 756.900 428.400 ;
        RECT 758.100 425.400 759.900 429.000 ;
        RECT 671.700 419.400 675.300 420.300 ;
        RECT 671.100 415.050 672.900 416.850 ;
        RECT 674.100 415.050 675.300 419.400 ;
        RECT 677.100 415.050 678.900 416.850 ;
        RECT 698.700 415.050 699.900 422.400 ;
        RECT 719.700 420.600 720.900 422.400 ;
        RECT 726.900 420.900 728.100 422.400 ;
        RECT 731.100 421.500 735.900 422.400 ;
        RECT 719.700 419.700 726.000 420.600 ;
        RECT 723.900 417.600 726.000 419.700 ;
        RECT 701.100 415.050 702.900 416.850 ;
        RECT 719.400 415.050 721.200 416.850 ;
        RECT 724.200 415.800 726.000 417.600 ;
        RECT 726.900 418.800 729.900 420.900 ;
        RECT 731.100 420.300 733.200 421.500 ;
        RECT 511.800 414.300 513.900 415.050 ;
        RECT 348.000 412.500 349.800 412.950 ;
        RECT 344.700 412.050 346.200 412.200 ;
        RECT 344.100 409.950 346.200 412.050 ;
        RECT 313.800 408.000 314.700 409.950 ;
        RECT 307.500 405.600 309.600 407.700 ;
        RECT 313.200 406.950 314.700 408.000 ;
        RECT 345.300 408.000 346.200 409.950 ;
        RECT 347.100 409.500 351.000 411.300 ;
        RECT 374.250 411.150 376.050 412.950 ;
        RECT 347.100 409.200 349.200 409.500 ;
        RECT 345.300 406.950 346.800 408.000 ;
        RECT 313.200 405.600 314.400 406.950 ;
        RECT 305.100 404.700 309.600 405.600 ;
        RECT 284.100 393.000 285.900 399.600 ;
        RECT 287.100 393.600 288.900 399.600 ;
        RECT 305.100 393.600 306.900 404.700 ;
        RECT 308.100 393.000 309.900 403.500 ;
        RECT 312.600 393.600 314.400 405.600 ;
        RECT 317.100 405.600 319.200 406.500 ;
        RECT 340.800 405.600 342.900 406.500 ;
        RECT 317.100 404.400 321.900 405.600 ;
        RECT 317.100 393.000 318.900 403.500 ;
        RECT 320.100 393.600 321.900 404.400 ;
        RECT 338.100 404.400 342.900 405.600 ;
        RECT 345.600 405.600 346.800 406.950 ;
        RECT 350.400 405.600 352.500 407.700 ;
        RECT 380.700 405.600 381.600 412.950 ;
        RECT 401.100 411.150 402.900 412.950 ;
        RECT 405.000 407.400 405.900 412.950 ;
        RECT 406.950 411.150 408.750 412.950 ;
        RECT 431.100 411.150 432.900 412.950 ;
        RECT 401.100 406.500 405.900 407.400 ;
        RECT 409.950 408.450 412.050 409.050 ;
        RECT 415.950 408.450 418.050 409.050 ;
        RECT 409.950 407.550 418.050 408.450 ;
        RECT 409.950 406.950 412.050 407.550 ;
        RECT 415.950 406.950 418.050 407.550 ;
        RECT 427.950 408.450 430.050 409.050 ;
        RECT 433.950 408.450 436.050 408.750 ;
        RECT 427.950 407.550 436.050 408.450 ;
        RECT 427.950 406.950 430.050 407.550 ;
        RECT 433.950 406.650 436.050 407.550 ;
        RECT 338.100 393.600 339.900 404.400 ;
        RECT 341.100 393.000 342.900 403.500 ;
        RECT 345.600 393.600 347.400 405.600 ;
        RECT 350.400 404.700 354.900 405.600 ;
        RECT 350.100 393.000 351.900 403.500 ;
        RECT 353.100 393.600 354.900 404.700 ;
        RECT 371.100 404.700 378.900 405.600 ;
        RECT 371.100 393.600 372.900 404.700 ;
        RECT 374.100 393.000 375.900 403.800 ;
        RECT 377.100 393.600 378.900 404.700 ;
        RECT 380.100 393.600 381.900 405.600 ;
        RECT 382.950 399.450 385.050 400.050 ;
        RECT 388.950 399.450 391.050 400.050 ;
        RECT 382.950 398.550 391.050 399.450 ;
        RECT 382.950 397.950 385.050 398.550 ;
        RECT 388.950 397.950 391.050 398.550 ;
        RECT 398.100 394.500 399.900 405.600 ;
        RECT 401.100 395.400 402.900 406.500 ;
        RECT 404.100 404.400 411.900 405.300 ;
        RECT 404.100 394.500 405.900 404.400 ;
        RECT 398.100 393.600 405.900 394.500 ;
        RECT 407.100 393.000 408.900 403.500 ;
        RECT 410.100 393.600 411.900 404.400 ;
        RECT 437.100 400.800 438.000 412.950 ;
        RECT 439.950 408.450 442.050 408.750 ;
        RECT 451.950 408.450 454.050 409.050 ;
        RECT 439.950 407.550 454.050 408.450 ;
        RECT 439.950 406.650 442.050 407.550 ;
        RECT 451.950 406.950 454.050 407.550 ;
        RECT 431.400 399.900 438.000 400.800 ;
        RECT 431.400 399.600 432.900 399.900 ;
        RECT 428.100 393.000 429.900 399.600 ;
        RECT 431.100 393.600 432.900 399.600 ;
        RECT 437.100 399.600 438.000 399.900 ;
        RECT 455.700 399.600 456.900 412.950 ;
        RECT 458.100 411.150 459.900 412.950 ;
        RECT 476.700 399.600 477.900 412.950 ;
        RECT 479.100 411.150 480.900 412.950 ;
        RECT 497.400 411.150 499.200 412.950 ;
        RECT 503.700 412.200 506.100 413.100 ;
        RECT 507.000 412.950 513.900 414.300 ;
        RECT 529.950 412.950 532.050 415.050 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 553.950 412.950 556.050 415.050 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 574.950 412.950 577.050 415.050 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 649.950 412.950 652.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 712.950 414.450 715.050 415.050 ;
        RECT 707.550 413.550 715.050 414.450 ;
        RECT 507.000 412.500 508.800 412.950 ;
        RECT 503.700 412.050 505.200 412.200 ;
        RECT 503.100 409.950 505.200 412.050 ;
        RECT 504.300 408.000 505.200 409.950 ;
        RECT 506.100 409.500 510.000 411.300 ;
        RECT 530.250 411.150 532.050 412.950 ;
        RECT 506.100 409.200 508.200 409.500 ;
        RECT 504.300 406.950 505.800 408.000 ;
        RECT 499.800 405.600 501.900 406.500 ;
        RECT 497.100 404.400 501.900 405.600 ;
        RECT 504.600 405.600 505.800 406.950 ;
        RECT 509.400 405.600 511.500 407.700 ;
        RECT 533.400 405.600 534.300 412.950 ;
        RECT 536.100 411.150 537.900 412.950 ;
        RECT 554.250 411.150 556.050 412.950 ;
        RECT 557.400 405.600 558.300 412.950 ;
        RECT 560.100 411.150 561.900 412.950 ;
        RECT 575.700 405.600 576.900 412.950 ;
        RECT 599.250 411.150 601.050 412.950 ;
        RECT 605.700 405.600 606.600 412.950 ;
        RECT 626.250 411.150 628.050 412.950 ;
        RECT 632.700 405.600 633.600 412.950 ;
        RECT 434.100 393.000 435.900 399.000 ;
        RECT 437.100 393.600 438.900 399.600 ;
        RECT 455.100 393.600 456.900 399.600 ;
        RECT 458.100 393.000 459.900 399.600 ;
        RECT 476.100 393.600 477.900 399.600 ;
        RECT 479.100 393.000 480.900 399.600 ;
        RECT 497.100 393.600 498.900 404.400 ;
        RECT 500.100 393.000 501.900 403.500 ;
        RECT 504.600 393.600 506.400 405.600 ;
        RECT 509.400 404.700 513.900 405.600 ;
        RECT 509.100 393.000 510.900 403.500 ;
        RECT 512.100 393.600 513.900 404.700 ;
        RECT 530.100 393.000 531.900 405.600 ;
        RECT 533.400 404.400 537.000 405.600 ;
        RECT 535.200 393.600 537.000 404.400 ;
        RECT 554.100 393.000 555.900 405.600 ;
        RECT 557.400 404.400 561.000 405.600 ;
        RECT 559.200 393.600 561.000 404.400 ;
        RECT 575.100 393.600 576.900 405.600 ;
        RECT 578.100 393.000 579.900 405.600 ;
        RECT 596.100 404.700 603.900 405.600 ;
        RECT 596.100 393.600 597.900 404.700 ;
        RECT 599.100 393.000 600.900 403.800 ;
        RECT 602.100 393.600 603.900 404.700 ;
        RECT 605.100 393.600 606.900 405.600 ;
        RECT 623.100 404.700 630.900 405.600 ;
        RECT 623.100 393.600 624.900 404.700 ;
        RECT 626.100 393.000 627.900 403.800 ;
        RECT 629.100 393.600 630.900 404.700 ;
        RECT 632.100 393.600 633.900 405.600 ;
        RECT 650.700 399.600 651.900 412.950 ;
        RECT 653.100 411.150 654.900 412.950 ;
        RECT 674.100 405.600 675.300 412.950 ;
        RECT 680.100 411.150 681.900 412.950 ;
        RECT 698.700 405.600 699.900 412.950 ;
        RECT 707.550 412.050 708.450 413.550 ;
        RECT 712.950 412.950 715.050 413.550 ;
        RECT 719.100 414.300 721.200 415.050 ;
        RECT 719.100 412.950 726.000 414.300 ;
        RECT 724.200 412.500 726.000 412.950 ;
        RECT 726.900 413.100 728.100 418.800 ;
        RECT 729.000 415.800 731.100 417.900 ;
        RECT 729.300 414.000 731.100 415.800 ;
        RECT 755.400 415.050 756.300 425.400 ;
        RECT 776.100 423.300 777.900 428.400 ;
        RECT 779.100 424.200 780.900 429.000 ;
        RECT 782.100 423.300 783.900 428.400 ;
        RECT 776.100 421.950 783.900 423.300 ;
        RECT 785.100 422.400 786.900 428.400 ;
        RECT 803.100 422.400 804.900 428.400 ;
        RECT 806.100 422.400 807.900 429.000 ;
        RECT 824.700 425.400 826.500 429.000 ;
        RECT 827.700 423.600 829.500 428.400 ;
        RECT 824.400 422.400 829.500 423.600 ;
        RECT 832.200 422.400 834.000 429.000 ;
        RECT 851.100 424.200 852.900 427.200 ;
        RECT 854.100 426.600 855.300 429.000 ;
        RECT 863.100 427.200 864.300 429.000 ;
        RECT 757.950 420.450 760.050 421.050 ;
        RECT 772.950 420.450 775.050 421.050 ;
        RECT 757.950 419.550 775.050 420.450 ;
        RECT 785.100 420.300 786.300 422.400 ;
        RECT 757.950 418.950 760.050 419.550 ;
        RECT 772.950 418.950 775.050 419.550 ;
        RECT 782.700 419.400 786.300 420.300 ;
        RECT 779.100 415.050 780.900 416.850 ;
        RECT 782.700 415.050 783.900 419.400 ;
        RECT 785.100 415.050 786.900 416.850 ;
        RECT 803.700 415.050 804.900 422.400 ;
        RECT 806.100 415.050 807.900 416.850 ;
        RECT 824.400 415.050 825.300 422.400 ;
        RECT 851.100 420.900 852.000 424.200 ;
        RECT 854.100 421.800 855.900 426.600 ;
        RECT 858.600 422.700 860.400 427.200 ;
        RECT 858.600 421.800 860.700 422.700 ;
        RECT 851.100 420.000 858.300 420.900 ;
        RECT 826.950 415.050 828.750 416.850 ;
        RECT 833.100 415.050 834.900 416.850 ;
        RECT 851.100 415.050 852.900 416.850 ;
        RECT 726.900 412.200 729.300 413.100 ;
        RECT 703.950 410.550 708.450 412.050 ;
        RECT 727.800 412.050 729.300 412.200 ;
        RECT 733.800 412.950 735.900 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 757.950 412.950 760.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 802.950 412.950 805.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 851.100 412.950 853.200 415.050 ;
        RECT 854.100 412.950 856.200 415.050 ;
        RECT 857.100 412.950 858.300 420.000 ;
        RECT 859.800 415.050 860.700 421.800 ;
        RECT 863.100 421.200 864.900 427.200 ;
        RECT 881.100 424.200 882.900 427.200 ;
        RECT 884.100 426.600 885.300 429.000 ;
        RECT 893.100 427.200 894.300 429.000 ;
        RECT 881.100 420.900 882.000 424.200 ;
        RECT 884.100 421.800 885.900 426.600 ;
        RECT 888.600 422.700 890.400 427.200 ;
        RECT 888.600 421.800 890.700 422.700 ;
        RECT 881.100 420.000 888.300 420.900 ;
        RECT 881.100 415.050 882.900 416.850 ;
        RECT 859.800 412.950 861.900 415.050 ;
        RECT 862.800 412.950 864.900 415.050 ;
        RECT 881.100 412.950 883.200 415.050 ;
        RECT 884.100 412.950 886.200 415.050 ;
        RECT 887.100 412.950 888.300 420.000 ;
        RECT 889.800 415.050 890.700 421.800 ;
        RECT 893.100 421.200 894.900 427.200 ;
        RECT 911.100 422.400 912.900 428.400 ;
        RECT 914.100 423.300 915.900 429.000 ;
        RECT 918.600 422.400 920.400 428.400 ;
        RECT 923.100 423.300 924.900 429.000 ;
        RECT 926.100 422.400 927.900 428.400 ;
        RECT 911.100 421.500 915.900 422.400 ;
        RECT 913.800 420.300 915.900 421.500 ;
        RECT 918.900 420.900 920.100 422.400 ;
        RECT 917.100 418.800 920.100 420.900 ;
        RECT 926.100 420.600 927.300 422.400 ;
        RECT 915.900 415.800 918.000 417.900 ;
        RECT 889.800 412.950 891.900 415.050 ;
        RECT 892.800 412.950 894.900 415.050 ;
        RECT 911.100 412.950 913.200 415.050 ;
        RECT 915.900 414.000 917.700 415.800 ;
        RECT 918.900 413.100 920.100 418.800 ;
        RECT 921.000 419.700 927.300 420.600 ;
        RECT 944.700 421.200 946.500 428.400 ;
        RECT 949.800 422.400 951.600 429.000 ;
        RECT 965.100 425.400 966.900 429.000 ;
        RECT 968.100 425.400 969.900 428.400 ;
        RECT 971.100 425.400 972.900 429.000 ;
        RECT 944.700 420.300 948.900 421.200 ;
        RECT 921.000 417.600 923.100 419.700 ;
        RECT 921.000 415.800 922.800 417.600 ;
        RECT 925.800 415.050 927.600 416.850 ;
        RECT 944.100 415.050 945.900 416.850 ;
        RECT 947.700 415.050 948.900 420.300 ;
        RECT 952.950 420.450 955.050 421.050 ;
        RECT 964.950 420.450 967.050 421.050 ;
        RECT 952.950 419.550 967.050 420.450 ;
        RECT 952.950 418.950 955.050 419.550 ;
        RECT 964.950 418.950 967.050 419.550 ;
        RECT 949.950 415.050 951.750 416.850 ;
        RECT 968.400 415.050 969.300 425.400 ;
        RECT 989.700 421.200 991.500 428.400 ;
        RECT 994.800 422.400 996.600 429.000 ;
        RECT 989.700 420.300 993.900 421.200 ;
        RECT 973.950 417.450 976.050 418.050 ;
        RECT 979.950 417.450 982.050 418.050 ;
        RECT 973.950 416.550 982.050 417.450 ;
        RECT 973.950 415.950 976.050 416.550 ;
        RECT 979.950 415.950 982.050 416.550 ;
        RECT 989.100 415.050 990.900 416.850 ;
        RECT 992.700 415.050 993.900 420.300 ;
        RECT 1015.500 420.000 1017.300 428.400 ;
        RECT 1014.000 418.800 1017.300 420.000 ;
        RECT 1022.100 419.400 1023.900 429.000 ;
        RECT 994.950 415.050 996.750 416.850 ;
        RECT 1014.000 415.050 1014.900 418.800 ;
        RECT 1016.100 415.050 1017.900 416.850 ;
        RECT 1022.100 415.050 1023.900 416.850 ;
        RECT 925.800 414.300 927.900 415.050 ;
        RECT 703.950 409.950 708.000 410.550 ;
        RECT 723.000 409.500 726.900 411.300 ;
        RECT 724.800 409.200 726.900 409.500 ;
        RECT 727.800 409.950 729.900 412.050 ;
        RECT 733.800 411.150 735.600 412.950 ;
        RECT 752.250 411.150 754.050 412.950 ;
        RECT 727.800 408.000 728.700 409.950 ;
        RECT 721.500 405.600 723.600 407.700 ;
        RECT 727.200 406.950 728.700 408.000 ;
        RECT 727.200 405.600 728.400 406.950 ;
        RECT 674.100 404.100 676.500 405.600 ;
        RECT 672.000 401.100 673.800 402.900 ;
        RECT 650.100 393.600 651.900 399.600 ;
        RECT 653.100 393.000 654.900 399.600 ;
        RECT 671.700 393.000 673.500 399.600 ;
        RECT 674.700 393.600 676.500 404.100 ;
        RECT 679.800 393.000 681.600 405.600 ;
        RECT 698.100 393.600 699.900 405.600 ;
        RECT 701.100 393.000 702.900 405.600 ;
        RECT 719.100 404.700 723.600 405.600 ;
        RECT 719.100 393.600 720.900 404.700 ;
        RECT 722.100 393.000 723.900 403.500 ;
        RECT 726.600 393.600 728.400 405.600 ;
        RECT 731.100 405.600 733.200 406.500 ;
        RECT 755.400 405.600 756.300 412.950 ;
        RECT 758.100 411.150 759.900 412.950 ;
        RECT 776.100 411.150 777.900 412.950 ;
        RECT 782.700 405.600 783.900 412.950 ;
        RECT 803.700 405.600 804.900 412.950 ;
        RECT 824.400 405.600 825.300 412.950 ;
        RECT 829.950 411.150 831.750 412.950 ;
        RECT 854.100 411.150 855.900 412.950 ;
        RECT 857.100 411.150 858.900 412.950 ;
        RECT 829.950 408.450 832.050 409.050 ;
        RECT 847.950 408.450 850.050 409.050 ;
        RECT 829.950 407.550 850.050 408.450 ;
        RECT 829.950 406.950 832.050 407.550 ;
        RECT 847.950 406.950 850.050 407.550 ;
        RECT 857.700 406.800 858.900 411.150 ;
        RECT 851.100 405.900 858.900 406.800 ;
        RECT 731.100 404.400 735.900 405.600 ;
        RECT 731.100 393.000 732.900 403.500 ;
        RECT 734.100 393.600 735.900 404.400 ;
        RECT 752.100 393.000 753.900 405.600 ;
        RECT 755.400 404.400 759.000 405.600 ;
        RECT 757.200 393.600 759.000 404.400 ;
        RECT 776.400 393.000 778.200 405.600 ;
        RECT 781.500 404.100 783.900 405.600 ;
        RECT 781.500 393.600 783.300 404.100 ;
        RECT 784.200 401.100 786.000 402.900 ;
        RECT 784.500 393.000 786.300 399.600 ;
        RECT 803.100 393.600 804.900 405.600 ;
        RECT 806.100 393.000 807.900 405.600 ;
        RECT 824.100 393.600 825.900 405.600 ;
        RECT 827.100 404.700 834.900 405.600 ;
        RECT 827.100 393.600 828.900 404.700 ;
        RECT 830.100 393.000 831.900 403.800 ;
        RECT 833.100 393.600 834.900 404.700 ;
        RECT 851.100 400.800 852.000 405.900 ;
        RECT 859.800 405.000 860.700 412.950 ;
        RECT 862.800 411.150 864.600 412.950 ;
        RECT 884.100 411.150 885.900 412.950 ;
        RECT 887.100 411.150 888.900 412.950 ;
        RECT 887.700 406.800 888.900 411.150 ;
        RECT 881.100 405.900 888.900 406.800 ;
        RECT 851.100 394.800 852.900 400.800 ;
        RECT 854.100 393.000 855.900 405.000 ;
        RECT 858.600 404.100 860.700 405.000 ;
        RECT 858.600 393.600 860.400 404.100 ;
        RECT 863.100 393.000 864.900 405.600 ;
        RECT 881.100 400.800 882.000 405.900 ;
        RECT 889.800 405.000 890.700 412.950 ;
        RECT 892.800 411.150 894.600 412.950 ;
        RECT 911.400 411.150 913.200 412.950 ;
        RECT 917.700 412.200 920.100 413.100 ;
        RECT 921.000 412.950 927.900 414.300 ;
        RECT 943.950 412.950 946.050 415.050 ;
        RECT 946.950 412.950 949.050 415.050 ;
        RECT 949.950 412.950 952.050 415.050 ;
        RECT 964.950 412.950 967.050 415.050 ;
        RECT 967.950 412.950 970.050 415.050 ;
        RECT 970.950 412.950 973.050 415.050 ;
        RECT 988.950 412.950 991.050 415.050 ;
        RECT 991.950 412.950 994.050 415.050 ;
        RECT 994.950 412.950 997.050 415.050 ;
        RECT 1012.950 412.950 1015.050 415.050 ;
        RECT 1015.950 412.950 1018.050 415.050 ;
        RECT 1018.950 412.950 1021.050 415.050 ;
        RECT 1021.950 412.950 1024.050 415.050 ;
        RECT 921.000 412.500 922.800 412.950 ;
        RECT 917.700 412.050 919.200 412.200 ;
        RECT 917.100 409.950 919.200 412.050 ;
        RECT 918.300 408.000 919.200 409.950 ;
        RECT 920.100 409.500 924.000 411.300 ;
        RECT 920.100 409.200 922.200 409.500 ;
        RECT 918.300 406.950 919.800 408.000 ;
        RECT 913.800 405.600 915.900 406.500 ;
        RECT 881.100 394.800 882.900 400.800 ;
        RECT 884.100 393.000 885.900 405.000 ;
        RECT 888.600 404.100 890.700 405.000 ;
        RECT 888.600 393.600 890.400 404.100 ;
        RECT 893.100 393.000 894.900 405.600 ;
        RECT 911.100 404.400 915.900 405.600 ;
        RECT 918.600 405.600 919.800 406.950 ;
        RECT 923.400 405.600 925.500 407.700 ;
        RECT 911.100 393.600 912.900 404.400 ;
        RECT 914.100 393.000 915.900 403.500 ;
        RECT 918.600 393.600 920.400 405.600 ;
        RECT 923.400 404.700 927.900 405.600 ;
        RECT 923.100 393.000 924.900 403.500 ;
        RECT 926.100 393.600 927.900 404.700 ;
        RECT 947.700 399.600 948.900 412.950 ;
        RECT 952.950 411.450 955.050 412.050 ;
        RECT 958.950 411.450 961.050 412.050 ;
        RECT 952.950 410.550 961.050 411.450 ;
        RECT 965.250 411.150 967.050 412.950 ;
        RECT 952.950 409.950 955.050 410.550 ;
        RECT 958.950 409.950 961.050 410.550 ;
        RECT 968.400 405.600 969.300 412.950 ;
        RECT 971.100 411.150 972.900 412.950 ;
        RECT 944.100 393.000 945.900 399.600 ;
        RECT 947.100 393.600 948.900 399.600 ;
        RECT 950.100 393.000 951.900 399.600 ;
        RECT 965.100 393.000 966.900 405.600 ;
        RECT 968.400 404.400 972.000 405.600 ;
        RECT 970.200 393.600 972.000 404.400 ;
        RECT 992.700 399.600 993.900 412.950 ;
        RECT 1014.000 400.800 1014.900 412.950 ;
        RECT 1019.100 411.150 1020.900 412.950 ;
        RECT 1014.000 399.900 1020.600 400.800 ;
        RECT 1014.000 399.600 1014.900 399.900 ;
        RECT 989.100 393.000 990.900 399.600 ;
        RECT 992.100 393.600 993.900 399.600 ;
        RECT 995.100 393.000 996.900 399.600 ;
        RECT 1013.100 393.600 1014.900 399.600 ;
        RECT 1019.100 399.600 1020.600 399.900 ;
        RECT 1016.100 393.000 1017.900 399.000 ;
        RECT 1019.100 393.600 1020.900 399.600 ;
        RECT 1022.100 393.000 1023.900 399.600 ;
        RECT 17.100 383.400 18.900 389.400 ;
        RECT 20.100 383.400 21.900 390.000 ;
        RECT 17.700 370.050 18.900 383.400 ;
        RECT 38.100 377.400 39.900 389.400 ;
        RECT 41.100 378.300 42.900 389.400 ;
        RECT 44.100 379.200 45.900 390.000 ;
        RECT 47.100 378.300 48.900 389.400 ;
        RECT 41.100 377.400 48.900 378.300 ;
        RECT 66.000 378.600 67.800 389.400 ;
        RECT 66.000 377.400 69.600 378.600 ;
        RECT 71.100 377.400 72.900 390.000 ;
        RECT 89.100 377.400 90.900 390.000 ;
        RECT 94.200 378.600 96.000 389.400 ;
        RECT 113.100 383.400 114.900 390.000 ;
        RECT 116.100 383.400 117.900 389.400 ;
        RECT 119.100 384.000 120.900 390.000 ;
        RECT 116.400 383.100 117.900 383.400 ;
        RECT 122.100 383.400 123.900 389.400 ;
        RECT 122.100 383.100 123.000 383.400 ;
        RECT 116.400 382.200 123.000 383.100 ;
        RECT 92.400 377.400 96.000 378.600 ;
        RECT 20.100 370.050 21.900 371.850 ;
        RECT 38.400 370.050 39.300 377.400 ;
        RECT 43.950 375.450 46.050 376.050 ;
        RECT 52.950 375.450 55.050 376.050 ;
        RECT 43.950 374.550 55.050 375.450 ;
        RECT 43.950 373.950 46.050 374.550 ;
        RECT 52.950 373.950 55.050 374.550 ;
        RECT 43.950 370.050 45.750 371.850 ;
        RECT 65.100 370.050 66.900 371.850 ;
        RECT 68.700 370.050 69.600 377.400 ;
        RECT 70.950 370.050 72.750 371.850 ;
        RECT 89.250 370.050 91.050 371.850 ;
        RECT 92.400 370.050 93.300 377.400 ;
        RECT 94.950 375.450 97.050 376.050 ;
        RECT 118.950 375.450 121.050 376.050 ;
        RECT 94.950 374.550 121.050 375.450 ;
        RECT 94.950 373.950 97.050 374.550 ;
        RECT 118.950 373.950 121.050 374.550 ;
        RECT 95.100 370.050 96.900 371.850 ;
        RECT 116.100 370.050 117.900 371.850 ;
        RECT 122.100 370.050 123.000 382.200 ;
        RECT 141.000 378.600 142.800 389.400 ;
        RECT 141.000 377.400 144.600 378.600 ;
        RECT 146.100 377.400 147.900 390.000 ;
        RECT 164.700 383.400 166.500 390.000 ;
        RECT 165.000 380.100 166.800 381.900 ;
        RECT 167.700 378.900 169.500 389.400 ;
        RECT 167.100 377.400 169.500 378.900 ;
        RECT 172.800 377.400 174.600 390.000 ;
        RECT 191.100 383.400 192.900 389.400 ;
        RECT 194.100 383.400 195.900 390.000 ;
        RECT 212.100 383.400 213.900 389.400 ;
        RECT 215.100 383.400 216.900 390.000 ;
        RECT 140.100 370.050 141.900 371.850 ;
        RECT 143.700 370.050 144.600 377.400 ;
        RECT 145.950 370.050 147.750 371.850 ;
        RECT 167.100 370.050 168.300 377.400 ;
        RECT 173.100 370.050 174.900 371.850 ;
        RECT 191.700 370.050 192.900 383.400 ;
        RECT 196.950 372.450 199.050 373.050 ;
        RECT 205.950 372.450 208.050 373.050 ;
        RECT 194.100 370.050 195.900 371.850 ;
        RECT 196.950 371.550 208.050 372.450 ;
        RECT 196.950 370.950 199.050 371.550 ;
        RECT 205.950 370.950 208.050 371.550 ;
        RECT 212.700 370.050 213.900 383.400 ;
        RECT 233.400 377.400 235.200 390.000 ;
        RECT 238.500 378.900 240.300 389.400 ;
        RECT 241.500 383.400 243.300 390.000 ;
        RECT 260.100 383.400 261.900 390.000 ;
        RECT 263.100 383.400 264.900 389.400 ;
        RECT 266.100 383.400 267.900 390.000 ;
        RECT 241.200 380.100 243.000 381.900 ;
        RECT 238.500 377.400 240.900 378.900 ;
        RECT 217.950 372.450 222.000 373.050 ;
        RECT 215.100 370.050 216.900 371.850 ;
        RECT 217.950 370.950 222.450 372.450 ;
        RECT 221.550 370.050 222.450 370.950 ;
        RECT 233.100 370.050 234.900 371.850 ;
        RECT 239.700 370.050 240.900 377.400 ;
        RECT 263.700 370.050 264.900 383.400 ;
        RECT 284.400 377.400 286.200 390.000 ;
        RECT 289.500 378.900 291.300 389.400 ;
        RECT 292.500 383.400 294.300 390.000 ;
        RECT 311.100 383.400 312.900 390.000 ;
        RECT 314.100 383.400 315.900 389.400 ;
        RECT 317.100 383.400 318.900 390.000 ;
        RECT 335.100 383.400 336.900 390.000 ;
        RECT 338.100 383.400 339.900 389.400 ;
        RECT 341.100 384.000 342.900 390.000 ;
        RECT 292.200 380.100 294.000 381.900 ;
        RECT 289.500 377.400 291.900 378.900 ;
        RECT 284.100 370.050 285.900 371.850 ;
        RECT 290.700 370.050 291.900 377.400 ;
        RECT 292.950 375.450 295.050 376.050 ;
        RECT 301.950 375.450 304.050 376.050 ;
        RECT 292.950 374.550 304.050 375.450 ;
        RECT 292.950 373.950 295.050 374.550 ;
        RECT 301.950 373.950 304.050 374.550 ;
        RECT 314.100 370.050 315.300 383.400 ;
        RECT 338.400 383.100 339.900 383.400 ;
        RECT 344.100 383.400 345.900 389.400 ;
        RECT 344.100 383.100 345.000 383.400 ;
        RECT 338.400 382.200 345.000 383.100 ;
        RECT 338.100 370.050 339.900 371.850 ;
        RECT 344.100 370.050 345.000 382.200 ;
        RECT 362.100 379.500 363.900 389.400 ;
        RECT 365.100 380.400 366.900 390.000 ;
        RECT 368.100 388.500 375.900 389.400 ;
        RECT 368.100 379.500 369.900 388.500 ;
        RECT 362.100 378.600 369.900 379.500 ;
        RECT 371.100 379.800 372.900 387.600 ;
        RECT 374.100 380.700 375.900 388.500 ;
        RECT 377.100 388.500 384.900 389.400 ;
        RECT 377.100 379.800 378.900 388.500 ;
        RECT 371.100 378.900 378.900 379.800 ;
        RECT 380.100 379.800 381.900 387.600 ;
        RECT 365.100 370.050 366.900 371.850 ;
        RECT 374.250 370.050 376.050 371.850 ;
        RECT 380.100 370.050 381.300 379.800 ;
        RECT 383.100 379.200 384.900 388.500 ;
        RECT 401.100 383.400 402.900 390.000 ;
        RECT 404.100 383.400 405.900 389.400 ;
        RECT 16.950 367.950 19.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 67.950 367.950 70.050 370.050 ;
        RECT 70.950 367.950 73.050 370.050 ;
        RECT 88.950 367.950 91.050 370.050 ;
        RECT 91.950 367.950 94.050 370.050 ;
        RECT 94.950 367.950 97.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 221.550 369.900 225.000 370.050 ;
        RECT 221.550 368.550 226.050 369.900 ;
        RECT 222.000 367.950 226.050 368.550 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 364.800 367.950 366.900 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 373.950 367.950 376.050 370.050 ;
        RECT 379.500 367.950 381.600 370.050 ;
        RECT 401.100 367.950 403.200 370.050 ;
        RECT 17.700 357.600 18.900 367.950 ;
        RECT 38.400 360.600 39.300 367.950 ;
        RECT 40.950 366.150 42.750 367.950 ;
        RECT 47.100 366.150 48.900 367.950 ;
        RECT 38.400 359.400 43.500 360.600 ;
        RECT 17.100 354.600 18.900 357.600 ;
        RECT 20.100 354.000 21.900 357.600 ;
        RECT 38.700 354.000 40.500 357.600 ;
        RECT 41.700 354.600 43.500 359.400 ;
        RECT 46.200 354.000 48.000 360.600 ;
        RECT 68.700 357.600 69.600 367.950 ;
        RECT 92.400 357.600 93.300 367.950 ;
        RECT 113.100 366.150 114.900 367.950 ;
        RECT 119.100 366.150 120.900 367.950 ;
        RECT 122.100 364.200 123.000 367.950 ;
        RECT 65.100 354.000 66.900 357.600 ;
        RECT 68.100 354.600 69.900 357.600 ;
        RECT 71.100 354.000 72.900 357.600 ;
        RECT 89.100 354.000 90.900 357.600 ;
        RECT 92.100 354.600 93.900 357.600 ;
        RECT 95.100 354.000 96.900 357.600 ;
        RECT 113.100 354.000 114.900 363.600 ;
        RECT 119.700 363.000 123.000 364.200 ;
        RECT 119.700 354.600 121.500 363.000 ;
        RECT 143.700 357.600 144.600 367.950 ;
        RECT 164.100 366.150 165.900 367.950 ;
        RECT 167.100 363.600 168.300 367.950 ;
        RECT 170.100 366.150 171.900 367.950 ;
        RECT 164.700 362.700 168.300 363.600 ;
        RECT 164.700 360.600 165.900 362.700 ;
        RECT 140.100 354.000 141.900 357.600 ;
        RECT 143.100 354.600 144.900 357.600 ;
        RECT 146.100 354.000 147.900 357.600 ;
        RECT 164.100 354.600 165.900 360.600 ;
        RECT 167.100 359.700 174.900 361.050 ;
        RECT 167.100 354.600 168.900 359.700 ;
        RECT 170.100 354.000 171.900 358.800 ;
        RECT 173.100 354.600 174.900 359.700 ;
        RECT 191.700 357.600 192.900 367.950 ;
        RECT 193.950 363.450 196.050 364.050 ;
        RECT 199.950 363.450 202.050 364.050 ;
        RECT 193.950 362.550 202.050 363.450 ;
        RECT 193.950 361.950 196.050 362.550 ;
        RECT 199.950 361.950 202.050 362.550 ;
        RECT 212.700 357.600 213.900 367.950 ;
        RECT 223.950 367.800 226.050 367.950 ;
        RECT 236.100 366.150 237.900 367.950 ;
        RECT 239.700 363.600 240.900 367.950 ;
        RECT 242.100 366.150 243.900 367.950 ;
        RECT 260.100 366.150 261.900 367.950 ;
        RECT 239.700 362.700 243.300 363.600 ;
        RECT 263.700 362.700 264.900 367.950 ;
        RECT 265.950 366.150 267.750 367.950 ;
        RECT 287.100 366.150 288.900 367.950 ;
        RECT 290.700 363.600 291.900 367.950 ;
        RECT 293.100 366.150 294.900 367.950 ;
        RECT 311.250 366.150 313.050 367.950 ;
        RECT 290.700 362.700 294.300 363.600 ;
        RECT 233.100 359.700 240.900 361.050 ;
        RECT 191.100 354.600 192.900 357.600 ;
        RECT 194.100 354.000 195.900 357.600 ;
        RECT 212.100 354.600 213.900 357.600 ;
        RECT 215.100 354.000 216.900 357.600 ;
        RECT 233.100 354.600 234.900 359.700 ;
        RECT 236.100 354.000 237.900 358.800 ;
        RECT 239.100 354.600 240.900 359.700 ;
        RECT 242.100 360.600 243.300 362.700 ;
        RECT 260.700 361.800 264.900 362.700 ;
        RECT 242.100 354.600 243.900 360.600 ;
        RECT 260.700 354.600 262.500 361.800 ;
        RECT 265.800 354.000 267.600 360.600 ;
        RECT 284.100 359.700 291.900 361.050 ;
        RECT 284.100 354.600 285.900 359.700 ;
        RECT 287.100 354.000 288.900 358.800 ;
        RECT 290.100 354.600 291.900 359.700 ;
        RECT 293.100 360.600 294.300 362.700 ;
        RECT 314.100 362.700 315.300 367.950 ;
        RECT 317.100 366.150 318.900 367.950 ;
        RECT 335.100 366.150 336.900 367.950 ;
        RECT 341.100 366.150 342.900 367.950 ;
        RECT 344.100 364.200 345.000 367.950 ;
        RECT 370.950 366.150 372.750 367.950 ;
        RECT 314.100 361.800 318.300 362.700 ;
        RECT 293.100 354.600 294.900 360.600 ;
        RECT 311.400 354.000 313.200 360.600 ;
        RECT 316.500 354.600 318.300 361.800 ;
        RECT 335.100 354.000 336.900 363.600 ;
        RECT 341.700 363.000 345.000 364.200 ;
        RECT 355.950 363.450 358.050 364.050 ;
        RECT 373.950 363.450 376.050 364.050 ;
        RECT 341.700 354.600 343.500 363.000 ;
        RECT 355.950 362.550 376.050 363.450 ;
        RECT 355.950 361.950 358.050 362.550 ;
        RECT 373.950 361.950 376.050 362.550 ;
        RECT 380.100 359.400 381.300 367.950 ;
        RECT 401.250 366.150 403.050 367.950 ;
        RECT 404.100 363.300 405.000 383.400 ;
        RECT 407.100 378.000 408.900 390.000 ;
        RECT 410.100 377.400 411.900 389.400 ;
        RECT 428.400 377.400 430.200 390.000 ;
        RECT 433.500 378.900 435.300 389.400 ;
        RECT 436.500 383.400 438.300 390.000 ;
        RECT 455.100 383.400 456.900 389.400 ;
        RECT 458.100 383.400 459.900 390.000 ;
        RECT 476.100 383.400 477.900 390.000 ;
        RECT 479.100 383.400 480.900 389.400 ;
        RECT 482.100 383.400 483.900 390.000 ;
        RECT 500.100 383.400 501.900 389.400 ;
        RECT 503.100 383.400 504.900 390.000 ;
        RECT 521.700 383.400 523.500 390.000 ;
        RECT 436.200 380.100 438.000 381.900 ;
        RECT 433.500 377.400 435.900 378.900 ;
        RECT 406.200 370.050 408.000 371.850 ;
        RECT 410.400 370.050 411.300 377.400 ;
        RECT 428.100 370.050 429.900 371.850 ;
        RECT 434.700 370.050 435.900 377.400 ;
        RECT 455.700 370.050 456.900 383.400 ;
        RECT 458.100 370.050 459.900 371.850 ;
        RECT 479.100 370.050 480.300 383.400 ;
        RECT 500.700 370.050 501.900 383.400 ;
        RECT 522.000 380.100 523.800 381.900 ;
        RECT 524.700 378.900 526.500 389.400 ;
        RECT 524.100 377.400 526.500 378.900 ;
        RECT 529.800 377.400 531.600 390.000 ;
        RECT 548.100 377.400 549.900 389.400 ;
        RECT 552.600 377.400 554.400 390.000 ;
        RECT 555.600 378.900 557.400 389.400 ;
        RECT 575.100 383.400 576.900 390.000 ;
        RECT 578.100 383.400 579.900 389.400 ;
        RECT 581.100 383.400 582.900 390.000 ;
        RECT 555.600 377.400 558.000 378.900 ;
        RECT 503.100 370.050 504.900 371.850 ;
        RECT 524.100 370.050 525.300 377.400 ;
        RECT 548.100 375.900 549.300 377.400 ;
        RECT 548.100 374.700 555.900 375.900 ;
        RECT 554.100 374.100 555.900 374.700 ;
        RECT 530.100 370.050 531.900 371.850 ;
        RECT 552.000 370.050 553.800 371.850 ;
        RECT 406.500 367.950 408.600 370.050 ;
        RECT 409.800 367.950 411.900 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 548.100 367.950 550.200 370.050 ;
        RECT 551.400 367.950 553.500 370.050 ;
        RECT 368.700 358.500 381.300 359.400 ;
        RECT 401.100 362.400 409.500 363.300 ;
        RECT 368.700 357.600 369.600 358.500 ;
        RECT 375.900 357.600 376.800 358.500 ;
        RECT 364.800 354.000 366.900 357.600 ;
        RECT 368.100 354.600 369.900 357.600 ;
        RECT 371.100 354.000 372.900 357.600 ;
        RECT 374.100 354.600 376.800 357.600 ;
        RECT 401.100 354.600 402.900 362.400 ;
        RECT 407.700 361.500 409.500 362.400 ;
        RECT 410.400 360.600 411.300 367.950 ;
        RECT 431.100 366.150 432.900 367.950 ;
        RECT 434.700 363.600 435.900 367.950 ;
        RECT 437.100 366.150 438.900 367.950 ;
        RECT 434.700 362.700 438.300 363.600 ;
        RECT 405.600 354.000 407.400 360.600 ;
        RECT 408.600 358.800 411.300 360.600 ;
        RECT 428.100 359.700 435.900 361.050 ;
        RECT 408.600 354.600 410.400 358.800 ;
        RECT 428.100 354.600 429.900 359.700 ;
        RECT 431.100 354.000 432.900 358.800 ;
        RECT 434.100 354.600 435.900 359.700 ;
        RECT 437.100 360.600 438.300 362.700 ;
        RECT 437.100 354.600 438.900 360.600 ;
        RECT 455.700 357.600 456.900 367.950 ;
        RECT 476.250 366.150 478.050 367.950 ;
        RECT 479.100 362.700 480.300 367.950 ;
        RECT 482.100 366.150 483.900 367.950 ;
        RECT 479.100 361.800 483.300 362.700 ;
        RECT 455.100 354.600 456.900 357.600 ;
        RECT 458.100 354.000 459.900 357.600 ;
        RECT 476.400 354.000 478.200 360.600 ;
        RECT 481.500 354.600 483.300 361.800 ;
        RECT 500.700 357.600 501.900 367.950 ;
        RECT 521.100 366.150 522.900 367.950 ;
        RECT 524.100 363.600 525.300 367.950 ;
        RECT 527.100 366.150 528.900 367.950 ;
        RECT 548.400 366.150 550.200 367.950 ;
        RECT 521.700 362.700 525.300 363.600 ;
        RECT 554.700 363.600 555.600 374.100 ;
        RECT 556.800 370.050 558.000 377.400 ;
        RECT 578.700 370.050 579.900 383.400 ;
        RECT 600.000 378.600 601.800 389.400 ;
        RECT 600.000 377.400 603.600 378.600 ;
        RECT 605.100 377.400 606.900 390.000 ;
        RECT 624.000 378.600 625.800 389.400 ;
        RECT 624.000 377.400 627.600 378.600 ;
        RECT 629.100 377.400 630.900 390.000 ;
        RECT 647.100 383.400 648.900 390.000 ;
        RECT 650.100 383.400 651.900 389.400 ;
        RECT 599.100 370.050 600.900 371.850 ;
        RECT 602.700 370.050 603.600 377.400 ;
        RECT 604.950 370.050 606.750 371.850 ;
        RECT 623.100 370.050 624.900 371.850 ;
        RECT 626.700 370.050 627.600 377.400 ;
        RECT 628.950 370.050 630.750 371.850 ;
        RECT 556.800 367.950 558.900 370.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 647.100 367.950 649.200 370.050 ;
        RECT 554.700 362.700 556.800 363.600 ;
        RECT 521.700 360.600 522.900 362.700 ;
        RECT 551.400 361.800 556.800 362.700 ;
        RECT 500.100 354.600 501.900 357.600 ;
        RECT 503.100 354.000 504.900 357.600 ;
        RECT 521.100 354.600 522.900 360.600 ;
        RECT 524.100 359.700 531.900 361.050 ;
        RECT 524.100 354.600 525.900 359.700 ;
        RECT 527.100 354.000 528.900 358.800 ;
        RECT 530.100 354.600 531.900 359.700 ;
        RECT 551.400 357.600 552.300 361.800 ;
        RECT 558.000 360.600 558.900 367.950 ;
        RECT 575.100 366.150 576.900 367.950 ;
        RECT 578.700 362.700 579.900 367.950 ;
        RECT 580.950 366.150 582.750 367.950 ;
        RECT 548.100 354.600 549.900 357.600 ;
        RECT 551.100 354.600 552.900 357.600 ;
        RECT 548.100 354.000 549.300 354.600 ;
        RECT 554.100 354.000 555.900 360.000 ;
        RECT 557.100 354.600 558.900 360.600 ;
        RECT 575.700 361.800 579.900 362.700 ;
        RECT 575.700 354.600 577.500 361.800 ;
        RECT 580.800 354.000 582.600 360.600 ;
        RECT 602.700 357.600 603.600 367.950 ;
        RECT 626.700 357.600 627.600 367.950 ;
        RECT 647.250 366.150 649.050 367.950 ;
        RECT 628.950 363.450 631.050 363.750 ;
        RECT 643.950 363.450 646.050 364.050 ;
        RECT 628.950 362.550 646.050 363.450 ;
        RECT 650.100 363.300 651.000 383.400 ;
        RECT 653.100 378.000 654.900 390.000 ;
        RECT 656.100 377.400 657.900 389.400 ;
        RECT 675.000 378.600 676.800 389.400 ;
        RECT 675.000 377.400 678.600 378.600 ;
        RECT 680.100 377.400 681.900 390.000 ;
        RECT 698.100 378.600 699.900 389.400 ;
        RECT 701.100 379.500 702.900 390.000 ;
        RECT 698.100 377.400 702.900 378.600 ;
        RECT 652.200 370.050 654.000 371.850 ;
        RECT 656.400 370.050 657.300 377.400 ;
        RECT 658.950 375.450 661.050 376.050 ;
        RECT 673.950 375.450 676.050 376.050 ;
        RECT 658.950 374.550 676.050 375.450 ;
        RECT 658.950 373.950 661.050 374.550 ;
        RECT 673.950 373.950 676.050 374.550 ;
        RECT 674.100 370.050 675.900 371.850 ;
        RECT 677.700 370.050 678.600 377.400 ;
        RECT 700.800 376.500 702.900 377.400 ;
        RECT 705.600 377.400 707.400 389.400 ;
        RECT 710.100 379.500 711.900 390.000 ;
        RECT 713.100 378.300 714.900 389.400 ;
        RECT 710.400 377.400 714.900 378.300 ;
        RECT 732.000 378.600 733.800 389.400 ;
        RECT 732.000 377.400 735.600 378.600 ;
        RECT 737.100 377.400 738.900 390.000 ;
        RECT 756.000 378.600 757.800 389.400 ;
        RECT 756.000 377.400 759.600 378.600 ;
        RECT 761.100 377.400 762.900 390.000 ;
        RECT 764.700 383.400 766.500 390.000 ;
        RECT 767.700 383.400 769.500 389.400 ;
        RECT 771.000 383.400 772.800 390.000 ;
        RECT 774.000 383.400 775.800 389.400 ;
        RECT 777.000 383.400 778.800 390.000 ;
        RECT 780.000 383.400 781.800 389.400 ;
        RECT 783.000 383.400 784.800 390.000 ;
        RECT 786.000 386.400 787.800 389.400 ;
        RECT 789.000 386.400 790.800 389.400 ;
        RECT 792.000 386.400 793.800 389.400 ;
        RECT 785.700 384.300 787.800 386.400 ;
        RECT 788.700 384.300 790.800 386.400 ;
        RECT 791.700 384.300 793.800 386.400 ;
        RECT 795.000 383.400 796.800 389.400 ;
        RECT 798.000 383.400 799.800 390.000 ;
        RECT 705.600 376.050 706.800 377.400 ;
        RECT 705.300 375.000 706.800 376.050 ;
        RECT 710.400 375.300 712.500 377.400 ;
        RECT 705.300 373.050 706.200 375.000 ;
        RECT 679.950 370.050 681.750 371.850 ;
        RECT 698.400 370.050 700.200 371.850 ;
        RECT 704.100 370.950 706.200 373.050 ;
        RECT 707.100 373.500 709.200 373.800 ;
        RECT 707.100 371.700 711.000 373.500 ;
        RECT 727.950 372.450 730.050 373.050 ;
        RECT 652.500 367.950 654.600 370.050 ;
        RECT 655.800 367.950 657.900 370.050 ;
        RECT 673.950 367.950 676.050 370.050 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 698.100 367.950 700.200 370.050 ;
        RECT 704.700 370.800 706.200 370.950 ;
        RECT 716.550 371.550 730.050 372.450 ;
        RECT 704.700 369.900 707.100 370.800 ;
        RECT 628.950 361.650 631.050 362.550 ;
        RECT 643.950 361.950 646.050 362.550 ;
        RECT 647.100 362.400 655.500 363.300 ;
        RECT 599.100 354.000 600.900 357.600 ;
        RECT 602.100 354.600 603.900 357.600 ;
        RECT 605.100 354.000 606.900 357.600 ;
        RECT 623.100 354.000 624.900 357.600 ;
        RECT 626.100 354.600 627.900 357.600 ;
        RECT 629.100 354.000 630.900 357.600 ;
        RECT 647.100 354.600 648.900 362.400 ;
        RECT 653.700 361.500 655.500 362.400 ;
        RECT 656.400 360.600 657.300 367.950 ;
        RECT 651.600 354.000 653.400 360.600 ;
        RECT 654.600 358.800 657.300 360.600 ;
        RECT 654.600 354.600 656.400 358.800 ;
        RECT 677.700 357.600 678.600 367.950 ;
        RECT 702.900 367.200 704.700 369.000 ;
        RECT 688.950 364.950 691.050 367.050 ;
        RECT 702.900 365.100 705.000 367.200 ;
        RECT 689.550 361.050 690.450 364.950 ;
        RECT 705.900 364.200 707.100 369.900 ;
        RECT 708.000 370.050 709.800 370.500 ;
        RECT 708.000 368.700 714.900 370.050 ;
        RECT 712.800 367.950 714.900 368.700 ;
        RECT 700.800 361.500 702.900 362.700 ;
        RECT 704.100 362.100 707.100 364.200 ;
        RECT 708.000 365.400 709.800 367.200 ;
        RECT 712.800 366.150 714.600 367.950 ;
        RECT 708.000 363.300 710.100 365.400 ;
        RECT 708.000 362.400 714.300 363.300 ;
        RECT 688.950 358.950 691.050 361.050 ;
        RECT 698.100 360.600 702.900 361.500 ;
        RECT 705.900 360.600 707.100 362.100 ;
        RECT 713.100 360.600 714.300 362.400 ;
        RECT 674.100 354.000 675.900 357.600 ;
        RECT 677.100 354.600 678.900 357.600 ;
        RECT 680.100 354.000 681.900 357.600 ;
        RECT 698.100 354.600 699.900 360.600 ;
        RECT 701.100 354.000 702.900 359.700 ;
        RECT 705.600 354.600 707.400 360.600 ;
        RECT 710.100 354.000 711.900 359.700 ;
        RECT 713.100 354.600 714.900 360.600 ;
        RECT 716.550 357.450 717.450 371.550 ;
        RECT 727.950 370.950 730.050 371.550 ;
        RECT 731.100 370.050 732.900 371.850 ;
        RECT 734.700 370.050 735.600 377.400 ;
        RECT 748.950 375.450 751.050 376.050 ;
        RECT 754.950 375.450 757.050 376.050 ;
        RECT 748.950 374.550 757.050 375.450 ;
        RECT 748.950 373.950 751.050 374.550 ;
        RECT 754.950 373.950 757.050 374.550 ;
        RECT 751.950 372.450 754.050 373.050 ;
        RECT 736.950 370.050 738.750 371.850 ;
        RECT 743.550 371.550 754.050 372.450 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 718.950 360.450 721.050 361.050 ;
        RECT 730.950 360.450 733.050 361.050 ;
        RECT 718.950 359.550 733.050 360.450 ;
        RECT 718.950 358.950 721.050 359.550 ;
        RECT 730.950 358.950 733.050 359.550 ;
        RECT 727.950 357.450 730.050 358.050 ;
        RECT 734.700 357.600 735.600 367.950 ;
        RECT 743.550 367.050 744.450 371.550 ;
        RECT 751.950 370.950 754.050 371.550 ;
        RECT 755.100 370.050 756.900 371.850 ;
        RECT 758.700 370.050 759.600 377.400 ;
        RECT 768.000 373.050 769.500 383.400 ;
        RECT 774.000 382.500 775.200 383.400 ;
        RECT 760.950 370.050 762.750 371.850 ;
        RECT 767.100 370.950 769.500 373.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 739.950 365.550 744.450 367.050 ;
        RECT 739.950 364.950 744.000 365.550 ;
        RECT 758.700 357.600 759.600 367.950 ;
        RECT 768.000 357.600 769.500 370.950 ;
        RECT 716.550 356.550 730.050 357.450 ;
        RECT 727.950 355.950 730.050 356.550 ;
        RECT 731.100 354.000 732.900 357.600 ;
        RECT 734.100 354.600 735.900 357.600 ;
        RECT 737.100 354.000 738.900 357.600 ;
        RECT 755.100 354.000 756.900 357.600 ;
        RECT 758.100 354.600 759.900 357.600 ;
        RECT 761.100 354.000 762.900 357.600 ;
        RECT 764.700 354.000 766.500 357.600 ;
        RECT 767.700 354.600 769.500 357.600 ;
        RECT 771.300 381.600 775.200 382.500 ;
        RECT 771.300 378.300 772.200 381.600 ;
        RECT 776.100 380.400 777.900 381.000 ;
        RECT 780.600 380.400 781.800 383.400 ;
        RECT 788.700 382.500 790.800 383.400 ;
        RECT 782.700 381.300 790.800 382.500 ;
        RECT 782.700 380.700 784.500 381.300 ;
        RECT 776.100 379.200 781.800 380.400 ;
        RECT 794.100 379.500 796.800 383.400 ;
        RECT 801.000 381.900 802.800 389.400 ;
        RECT 804.900 383.400 806.700 390.000 ;
        RECT 807.900 383.400 809.700 389.400 ;
        RECT 810.900 386.400 812.700 389.400 ;
        RECT 813.900 386.400 815.700 389.400 ;
        RECT 810.600 384.300 812.700 386.400 ;
        RECT 813.600 384.300 815.700 386.400 ;
        RECT 817.500 383.400 819.300 390.000 ;
        RECT 799.500 379.800 802.800 381.900 ;
        RECT 808.200 381.300 810.300 383.400 ;
        RECT 820.500 380.400 822.300 389.400 ;
        RECT 823.500 383.400 825.300 390.000 ;
        RECT 826.500 384.300 828.300 389.400 ;
        RECT 826.500 383.400 828.600 384.300 ;
        RECT 829.500 383.400 831.300 390.000 ;
        RECT 833.700 383.400 835.500 390.000 ;
        RECT 836.700 384.300 838.500 389.400 ;
        RECT 836.400 383.400 838.500 384.300 ;
        RECT 839.700 383.400 841.500 390.000 ;
        RECT 827.700 382.500 828.600 383.400 ;
        RECT 836.400 382.500 837.300 383.400 ;
        RECT 827.700 381.600 831.300 382.500 ;
        RECT 825.000 380.400 826.800 380.700 ;
        RECT 785.700 378.300 787.800 379.500 ;
        RECT 771.300 377.400 787.800 378.300 ;
        RECT 791.100 378.600 793.200 379.500 ;
        RECT 807.600 379.200 826.800 380.400 ;
        RECT 807.600 378.600 808.800 379.200 ;
        RECT 825.000 378.900 826.800 379.200 ;
        RECT 791.100 377.400 808.800 378.600 ;
        RECT 811.500 377.700 813.600 378.300 ;
        RECT 821.700 377.700 823.500 378.300 ;
        RECT 771.300 360.600 772.200 377.400 ;
        RECT 811.500 376.500 823.500 377.700 ;
        RECT 773.100 375.300 808.800 376.500 ;
        RECT 811.500 376.200 813.600 376.500 ;
        RECT 773.100 374.700 774.900 375.300 ;
        RECT 807.600 374.700 808.800 375.300 ;
        RECT 776.100 370.950 778.200 373.050 ;
        RECT 776.700 368.100 778.200 370.950 ;
        RECT 780.300 370.800 785.400 372.600 ;
        RECT 784.500 369.300 785.400 370.800 ;
        RECT 788.100 372.300 789.900 374.100 ;
        RECT 794.100 373.800 796.200 374.100 ;
        RECT 807.600 373.800 821.100 374.700 ;
        RECT 788.100 371.100 789.000 372.300 ;
        RECT 794.100 372.000 798.000 373.800 ;
        RECT 799.500 372.300 801.600 373.200 ;
        RECT 819.300 373.050 821.100 373.800 ;
        RECT 799.500 371.100 810.600 372.300 ;
        RECT 819.300 371.250 823.200 373.050 ;
        RECT 788.100 370.200 801.600 371.100 ;
        RECT 808.800 370.500 810.600 371.100 ;
        RECT 821.100 370.950 823.200 371.250 ;
        RECT 827.100 370.950 829.200 373.050 ;
        RECT 827.100 369.300 828.900 370.950 ;
        RECT 784.500 368.100 828.900 369.300 ;
        RECT 776.700 366.600 783.300 368.100 ;
        RECT 773.100 363.900 780.900 365.700 ;
        RECT 781.800 365.100 798.900 366.600 ;
        RECT 796.800 364.500 798.900 365.100 ;
        RECT 803.100 366.000 805.200 367.050 ;
        RECT 803.100 365.100 808.200 366.000 ;
        RECT 811.800 365.400 813.600 367.200 ;
        RECT 830.100 365.400 831.300 381.600 ;
        RECT 803.100 364.950 805.200 365.100 ;
        RECT 779.400 360.600 780.900 363.900 ;
        RECT 797.100 362.700 798.900 364.500 ;
        RECT 806.400 364.200 808.200 365.100 ;
        RECT 812.700 362.400 813.600 365.400 ;
        RECT 814.500 364.200 831.300 365.400 ;
        RECT 814.500 363.300 816.600 364.200 ;
        RECT 825.300 362.700 827.100 363.300 ;
        RECT 785.100 360.600 791.700 362.400 ;
        RECT 806.400 361.200 813.600 362.400 ;
        RECT 818.700 361.500 827.100 362.700 ;
        RECT 806.400 360.600 807.300 361.200 ;
        RECT 809.400 360.600 811.200 361.200 ;
        RECT 818.700 360.600 820.200 361.500 ;
        RECT 830.100 360.600 831.300 364.200 ;
        RECT 771.300 354.600 773.100 360.600 ;
        RECT 776.700 354.000 778.500 360.600 ;
        RECT 779.400 359.400 783.600 360.600 ;
        RECT 781.800 354.600 783.600 359.400 ;
        RECT 785.700 357.600 787.800 359.700 ;
        RECT 788.700 357.600 790.800 359.700 ;
        RECT 791.700 357.600 793.800 359.700 ;
        RECT 794.700 357.600 796.800 359.700 ;
        RECT 800.100 358.500 802.800 360.600 ;
        RECT 804.600 359.400 807.300 360.600 ;
        RECT 804.600 358.500 806.400 359.400 ;
        RECT 786.000 354.600 787.800 357.600 ;
        RECT 789.000 354.600 790.800 357.600 ;
        RECT 792.000 354.600 793.800 357.600 ;
        RECT 795.000 354.600 796.800 357.600 ;
        RECT 798.000 354.000 799.800 357.600 ;
        RECT 801.000 354.600 802.800 358.500 ;
        RECT 808.200 357.600 810.300 359.700 ;
        RECT 811.200 357.600 813.300 359.700 ;
        RECT 814.200 357.600 816.300 359.700 ;
        RECT 805.500 354.000 807.300 357.600 ;
        RECT 808.500 354.600 810.300 357.600 ;
        RECT 811.500 354.600 813.300 357.600 ;
        RECT 814.500 354.600 816.300 357.600 ;
        RECT 818.700 354.600 820.500 360.600 ;
        RECT 824.100 354.000 825.900 360.600 ;
        RECT 829.500 354.600 831.300 360.600 ;
        RECT 833.700 381.600 837.300 382.500 ;
        RECT 833.700 365.400 834.900 381.600 ;
        RECT 838.200 380.400 840.000 380.700 ;
        RECT 842.700 380.400 844.500 389.400 ;
        RECT 845.700 383.400 847.500 390.000 ;
        RECT 849.300 386.400 851.100 389.400 ;
        RECT 852.300 386.400 854.100 389.400 ;
        RECT 849.300 384.300 851.400 386.400 ;
        RECT 852.300 384.300 854.400 386.400 ;
        RECT 855.300 383.400 857.100 389.400 ;
        RECT 858.300 383.400 860.100 390.000 ;
        RECT 854.700 381.300 856.800 383.400 ;
        RECT 862.200 381.900 864.000 389.400 ;
        RECT 865.200 383.400 867.000 390.000 ;
        RECT 868.200 383.400 870.000 389.400 ;
        RECT 871.200 386.400 873.000 389.400 ;
        RECT 874.200 386.400 876.000 389.400 ;
        RECT 877.200 386.400 879.000 389.400 ;
        RECT 871.200 384.300 873.300 386.400 ;
        RECT 874.200 384.300 876.300 386.400 ;
        RECT 877.200 384.300 879.300 386.400 ;
        RECT 880.200 383.400 882.000 390.000 ;
        RECT 883.200 383.400 885.000 389.400 ;
        RECT 886.200 383.400 888.000 390.000 ;
        RECT 889.200 383.400 891.000 389.400 ;
        RECT 892.200 383.400 894.000 390.000 ;
        RECT 895.500 383.400 897.300 389.400 ;
        RECT 898.500 383.400 900.300 390.000 ;
        RECT 838.200 379.200 857.400 380.400 ;
        RECT 862.200 379.800 865.500 381.900 ;
        RECT 868.200 379.500 870.900 383.400 ;
        RECT 874.200 382.500 876.300 383.400 ;
        RECT 874.200 381.300 882.300 382.500 ;
        RECT 880.500 380.700 882.300 381.300 ;
        RECT 883.200 380.400 884.400 383.400 ;
        RECT 889.800 382.500 891.000 383.400 ;
        RECT 889.800 381.600 893.700 382.500 ;
        RECT 887.100 380.400 888.900 381.000 ;
        RECT 838.200 378.900 840.000 379.200 ;
        RECT 856.200 378.600 857.400 379.200 ;
        RECT 871.800 378.600 873.900 379.500 ;
        RECT 841.500 377.700 843.300 378.300 ;
        RECT 851.400 377.700 853.500 378.300 ;
        RECT 841.500 376.500 853.500 377.700 ;
        RECT 856.200 377.400 873.900 378.600 ;
        RECT 877.200 378.300 879.300 379.500 ;
        RECT 883.200 379.200 888.900 380.400 ;
        RECT 892.800 378.300 893.700 381.600 ;
        RECT 877.200 377.400 893.700 378.300 ;
        RECT 851.400 376.200 853.500 376.500 ;
        RECT 856.200 375.300 891.900 376.500 ;
        RECT 856.200 374.700 857.400 375.300 ;
        RECT 890.100 374.700 891.900 375.300 ;
        RECT 843.900 373.800 857.400 374.700 ;
        RECT 868.800 373.800 870.900 374.100 ;
        RECT 843.900 373.050 845.700 373.800 ;
        RECT 835.800 370.950 837.900 373.050 ;
        RECT 841.800 371.250 845.700 373.050 ;
        RECT 863.400 372.300 865.500 373.200 ;
        RECT 841.800 370.950 843.900 371.250 ;
        RECT 854.400 371.100 865.500 372.300 ;
        RECT 867.000 372.000 870.900 373.800 ;
        RECT 875.100 372.300 876.900 374.100 ;
        RECT 876.000 371.100 876.900 372.300 ;
        RECT 836.100 369.300 837.900 370.950 ;
        RECT 854.400 370.500 856.200 371.100 ;
        RECT 863.400 370.200 876.900 371.100 ;
        RECT 879.600 370.800 884.700 372.600 ;
        RECT 886.800 370.950 888.900 373.050 ;
        RECT 879.600 369.300 880.500 370.800 ;
        RECT 836.100 368.100 880.500 369.300 ;
        RECT 886.800 368.100 888.300 370.950 ;
        RECT 851.400 365.400 853.200 367.200 ;
        RECT 859.800 366.000 861.900 367.050 ;
        RECT 881.700 366.600 888.300 368.100 ;
        RECT 833.700 364.200 850.500 365.400 ;
        RECT 833.700 360.600 834.900 364.200 ;
        RECT 848.400 363.300 850.500 364.200 ;
        RECT 837.900 362.700 839.700 363.300 ;
        RECT 837.900 361.500 846.300 362.700 ;
        RECT 844.800 360.600 846.300 361.500 ;
        RECT 851.400 362.400 852.300 365.400 ;
        RECT 856.800 365.100 861.900 366.000 ;
        RECT 856.800 364.200 858.600 365.100 ;
        RECT 859.800 364.950 861.900 365.100 ;
        RECT 866.100 365.100 883.200 366.600 ;
        RECT 866.100 364.500 868.200 365.100 ;
        RECT 866.100 362.700 867.900 364.500 ;
        RECT 884.100 363.900 891.900 365.700 ;
        RECT 851.400 361.200 858.600 362.400 ;
        RECT 853.800 360.600 855.600 361.200 ;
        RECT 857.700 360.600 858.600 361.200 ;
        RECT 873.300 360.600 879.900 362.400 ;
        RECT 884.100 360.600 885.600 363.900 ;
        RECT 892.800 360.600 893.700 377.400 ;
        RECT 833.700 354.600 835.500 360.600 ;
        RECT 839.100 354.000 840.900 360.600 ;
        RECT 844.500 354.600 846.300 360.600 ;
        RECT 848.700 357.600 850.800 359.700 ;
        RECT 851.700 357.600 853.800 359.700 ;
        RECT 854.700 357.600 856.800 359.700 ;
        RECT 857.700 359.400 860.400 360.600 ;
        RECT 858.600 358.500 860.400 359.400 ;
        RECT 862.200 358.500 864.900 360.600 ;
        RECT 848.700 354.600 850.500 357.600 ;
        RECT 851.700 354.600 853.500 357.600 ;
        RECT 854.700 354.600 856.500 357.600 ;
        RECT 857.700 354.000 859.500 357.600 ;
        RECT 862.200 354.600 864.000 358.500 ;
        RECT 868.200 357.600 870.300 359.700 ;
        RECT 871.200 357.600 873.300 359.700 ;
        RECT 874.200 357.600 876.300 359.700 ;
        RECT 877.200 357.600 879.300 359.700 ;
        RECT 881.400 359.400 885.600 360.600 ;
        RECT 865.200 354.000 867.000 357.600 ;
        RECT 868.200 354.600 870.000 357.600 ;
        RECT 871.200 354.600 873.000 357.600 ;
        RECT 874.200 354.600 876.000 357.600 ;
        RECT 877.200 354.600 879.000 357.600 ;
        RECT 881.400 354.600 883.200 359.400 ;
        RECT 886.500 354.000 888.300 360.600 ;
        RECT 891.900 354.600 893.700 360.600 ;
        RECT 895.500 373.050 897.000 383.400 ;
        RECT 917.100 377.400 918.900 390.000 ;
        RECT 920.100 377.400 921.900 389.400 ;
        RECT 938.100 383.400 939.900 390.000 ;
        RECT 941.100 383.400 942.900 389.400 ;
        RECT 944.100 384.000 945.900 390.000 ;
        RECT 941.400 383.100 942.900 383.400 ;
        RECT 947.100 383.400 948.900 389.400 ;
        RECT 947.100 383.100 948.000 383.400 ;
        RECT 941.400 382.200 948.000 383.100 ;
        RECT 895.500 370.950 897.900 373.050 ;
        RECT 898.950 372.450 901.050 373.050 ;
        RECT 913.950 372.450 916.050 373.050 ;
        RECT 898.950 371.550 916.050 372.450 ;
        RECT 898.950 370.950 901.050 371.550 ;
        RECT 913.950 370.950 916.050 371.550 ;
        RECT 895.500 357.600 897.000 370.950 ;
        RECT 920.100 370.050 921.300 377.400 ;
        RECT 925.950 372.450 928.050 373.050 ;
        RECT 934.950 372.450 937.050 373.050 ;
        RECT 925.950 371.550 937.050 372.450 ;
        RECT 925.950 370.950 928.050 371.550 ;
        RECT 934.950 370.950 937.050 371.550 ;
        RECT 941.100 370.050 942.900 371.850 ;
        RECT 947.100 370.050 948.000 382.200 ;
        RECT 965.400 377.400 967.200 390.000 ;
        RECT 970.500 378.900 972.300 389.400 ;
        RECT 973.500 383.400 975.300 390.000 ;
        RECT 973.200 380.100 975.000 381.900 ;
        RECT 970.500 377.400 972.900 378.900 ;
        RECT 992.100 378.300 993.900 389.400 ;
        RECT 995.100 379.200 996.900 390.000 ;
        RECT 998.100 378.300 999.900 389.400 ;
        RECT 992.100 377.400 999.900 378.300 ;
        RECT 1001.100 377.400 1002.900 389.400 ;
        RECT 1019.700 383.400 1021.500 390.000 ;
        RECT 1020.000 380.100 1021.800 381.900 ;
        RECT 1022.700 378.900 1024.500 389.400 ;
        RECT 1022.100 377.400 1024.500 378.900 ;
        RECT 1027.800 377.400 1029.600 390.000 ;
        RECT 952.950 372.450 955.050 373.050 ;
        RECT 961.950 372.450 964.050 373.050 ;
        RECT 952.950 371.550 964.050 372.450 ;
        RECT 952.950 370.950 955.050 371.550 ;
        RECT 961.950 370.950 964.050 371.550 ;
        RECT 965.100 370.050 966.900 371.850 ;
        RECT 971.700 370.050 972.900 377.400 ;
        RECT 979.950 375.450 982.050 376.050 ;
        RECT 997.950 375.450 1000.050 376.050 ;
        RECT 979.950 374.550 1000.050 375.450 ;
        RECT 979.950 373.950 982.050 374.550 ;
        RECT 997.950 373.950 1000.050 374.550 ;
        RECT 982.950 372.450 985.050 373.050 ;
        RECT 988.950 372.450 991.050 373.050 ;
        RECT 982.950 371.550 991.050 372.450 ;
        RECT 982.950 370.950 985.050 371.550 ;
        RECT 988.950 370.950 991.050 371.550 ;
        RECT 995.250 370.050 997.050 371.850 ;
        RECT 1001.700 370.050 1002.600 377.400 ;
        RECT 1022.100 370.050 1023.300 377.400 ;
        RECT 1028.100 370.050 1029.900 371.850 ;
        RECT 916.950 367.950 919.050 370.050 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 937.950 367.950 940.050 370.050 ;
        RECT 940.950 367.950 943.050 370.050 ;
        RECT 943.950 367.950 946.050 370.050 ;
        RECT 946.950 367.950 949.050 370.050 ;
        RECT 964.950 367.950 967.050 370.050 ;
        RECT 967.950 367.950 970.050 370.050 ;
        RECT 970.950 367.950 973.050 370.050 ;
        RECT 973.950 367.950 976.050 370.050 ;
        RECT 991.950 367.950 994.050 370.050 ;
        RECT 994.950 367.950 997.050 370.050 ;
        RECT 997.950 367.950 1000.050 370.050 ;
        RECT 1000.950 367.950 1003.050 370.050 ;
        RECT 1018.950 367.950 1021.050 370.050 ;
        RECT 1021.950 367.950 1024.050 370.050 ;
        RECT 1024.950 367.950 1027.050 370.050 ;
        RECT 1027.950 367.950 1030.050 370.050 ;
        RECT 1033.950 369.450 1036.050 370.050 ;
        RECT 1039.950 369.450 1042.050 370.050 ;
        RECT 1033.950 368.550 1042.050 369.450 ;
        RECT 1033.950 367.950 1036.050 368.550 ;
        RECT 1039.950 367.950 1042.050 368.550 ;
        RECT 917.100 366.150 918.900 367.950 ;
        RECT 898.950 363.450 901.050 364.050 ;
        RECT 910.950 363.450 913.050 364.050 ;
        RECT 898.950 362.550 913.050 363.450 ;
        RECT 898.950 361.950 901.050 362.550 ;
        RECT 910.950 361.950 913.050 362.550 ;
        RECT 920.100 360.600 921.300 367.950 ;
        RECT 938.100 366.150 939.900 367.950 ;
        RECT 944.100 366.150 945.900 367.950 ;
        RECT 947.100 364.200 948.000 367.950 ;
        RECT 968.100 366.150 969.900 367.950 ;
        RECT 895.500 354.600 897.300 357.600 ;
        RECT 898.500 354.000 900.300 357.600 ;
        RECT 917.100 354.000 918.900 360.600 ;
        RECT 920.100 354.600 921.900 360.600 ;
        RECT 938.100 354.000 939.900 363.600 ;
        RECT 944.700 363.000 948.000 364.200 ;
        RECT 971.700 363.600 972.900 367.950 ;
        RECT 974.100 366.150 975.900 367.950 ;
        RECT 992.100 366.150 993.900 367.950 ;
        RECT 998.250 366.150 1000.050 367.950 ;
        RECT 944.700 354.600 946.500 363.000 ;
        RECT 971.700 362.700 975.300 363.600 ;
        RECT 965.100 359.700 972.900 361.050 ;
        RECT 965.100 354.600 966.900 359.700 ;
        RECT 968.100 354.000 969.900 358.800 ;
        RECT 971.100 354.600 972.900 359.700 ;
        RECT 974.100 360.600 975.300 362.700 ;
        RECT 1001.700 360.600 1002.600 367.950 ;
        RECT 1019.100 366.150 1020.900 367.950 ;
        RECT 1022.100 363.600 1023.300 367.950 ;
        RECT 1025.100 366.150 1026.900 367.950 ;
        RECT 1019.700 362.700 1023.300 363.600 ;
        RECT 1019.700 360.600 1020.900 362.700 ;
        RECT 974.100 354.600 975.900 360.600 ;
        RECT 993.000 354.000 994.800 360.600 ;
        RECT 997.500 359.400 1002.600 360.600 ;
        RECT 997.500 354.600 999.300 359.400 ;
        RECT 1000.500 354.000 1002.300 357.600 ;
        RECT 1019.100 354.600 1020.900 360.600 ;
        RECT 1022.100 359.700 1029.900 361.050 ;
        RECT 1022.100 354.600 1023.900 359.700 ;
        RECT 1025.100 354.000 1026.900 358.800 ;
        RECT 1028.100 354.600 1029.900 359.700 ;
        RECT 2.700 344.400 4.500 350.400 ;
        RECT 8.100 344.400 9.900 351.000 ;
        RECT 13.500 344.400 15.300 350.400 ;
        RECT 17.700 347.400 19.500 350.400 ;
        RECT 20.700 347.400 22.500 350.400 ;
        RECT 23.700 347.400 25.500 350.400 ;
        RECT 26.700 347.400 28.500 351.000 ;
        RECT 17.700 345.300 19.800 347.400 ;
        RECT 20.700 345.300 22.800 347.400 ;
        RECT 23.700 345.300 25.800 347.400 ;
        RECT 31.200 346.500 33.000 350.400 ;
        RECT 34.200 347.400 36.000 351.000 ;
        RECT 37.200 347.400 39.000 350.400 ;
        RECT 40.200 347.400 42.000 350.400 ;
        RECT 43.200 347.400 45.000 350.400 ;
        RECT 46.200 347.400 48.000 350.400 ;
        RECT 27.600 345.600 29.400 346.500 ;
        RECT 26.700 344.400 29.400 345.600 ;
        RECT 31.200 344.400 33.900 346.500 ;
        RECT 37.200 345.300 39.300 347.400 ;
        RECT 40.200 345.300 42.300 347.400 ;
        RECT 43.200 345.300 45.300 347.400 ;
        RECT 46.200 345.300 48.300 347.400 ;
        RECT 50.400 345.600 52.200 350.400 ;
        RECT 50.400 344.400 54.600 345.600 ;
        RECT 55.500 344.400 57.300 351.000 ;
        RECT 60.900 344.400 62.700 350.400 ;
        RECT 2.700 340.800 3.900 344.400 ;
        RECT 13.800 343.500 15.300 344.400 ;
        RECT 22.800 343.800 24.600 344.400 ;
        RECT 26.700 343.800 27.600 344.400 ;
        RECT 6.900 342.300 15.300 343.500 ;
        RECT 20.400 342.600 27.600 343.800 ;
        RECT 42.300 342.600 48.900 344.400 ;
        RECT 6.900 341.700 8.700 342.300 ;
        RECT 17.400 340.800 19.500 341.700 ;
        RECT 2.700 339.600 19.500 340.800 ;
        RECT 20.400 339.600 21.300 342.600 ;
        RECT 25.800 339.900 27.600 340.800 ;
        RECT 35.100 340.500 36.900 342.300 ;
        RECT 53.100 341.100 54.600 344.400 ;
        RECT 28.800 339.900 30.900 340.050 ;
        RECT 2.700 323.400 3.900 339.600 ;
        RECT 20.400 337.800 22.200 339.600 ;
        RECT 25.800 339.000 30.900 339.900 ;
        RECT 28.800 337.950 30.900 339.000 ;
        RECT 35.100 339.900 37.200 340.500 ;
        RECT 35.100 338.400 52.200 339.900 ;
        RECT 53.100 339.300 60.900 341.100 ;
        RECT 50.700 336.900 57.300 338.400 ;
        RECT 5.100 335.700 49.500 336.900 ;
        RECT 5.100 334.050 6.900 335.700 ;
        RECT 4.800 331.950 6.900 334.050 ;
        RECT 10.800 333.750 12.900 334.050 ;
        RECT 23.400 333.900 25.200 334.500 ;
        RECT 32.400 333.900 45.900 334.800 ;
        RECT 10.800 331.950 14.700 333.750 ;
        RECT 23.400 332.700 34.500 333.900 ;
        RECT 12.900 331.200 14.700 331.950 ;
        RECT 32.400 331.800 34.500 332.700 ;
        RECT 36.000 331.200 39.900 333.000 ;
        RECT 45.000 332.700 45.900 333.900 ;
        RECT 12.900 330.300 26.400 331.200 ;
        RECT 37.800 330.900 39.900 331.200 ;
        RECT 44.100 330.900 45.900 332.700 ;
        RECT 48.600 334.200 49.500 335.700 ;
        RECT 48.600 332.400 53.700 334.200 ;
        RECT 55.800 334.050 57.300 336.900 ;
        RECT 55.800 331.950 57.900 334.050 ;
        RECT 25.200 329.700 26.400 330.300 ;
        RECT 59.100 329.700 60.900 330.300 ;
        RECT 20.400 328.500 22.500 328.800 ;
        RECT 25.200 328.500 60.900 329.700 ;
        RECT 10.500 327.300 22.500 328.500 ;
        RECT 61.800 327.600 62.700 344.400 ;
        RECT 10.500 326.700 12.300 327.300 ;
        RECT 20.400 326.700 22.500 327.300 ;
        RECT 25.200 326.400 42.900 327.600 ;
        RECT 7.200 325.800 9.000 326.100 ;
        RECT 25.200 325.800 26.400 326.400 ;
        RECT 7.200 324.600 26.400 325.800 ;
        RECT 40.800 325.500 42.900 326.400 ;
        RECT 46.200 326.700 62.700 327.600 ;
        RECT 46.200 325.500 48.300 326.700 ;
        RECT 7.200 324.300 9.000 324.600 ;
        RECT 2.700 322.500 6.300 323.400 ;
        RECT 5.400 321.600 6.300 322.500 ;
        RECT 2.700 315.000 4.500 321.600 ;
        RECT 5.400 320.700 7.500 321.600 ;
        RECT 5.700 315.600 7.500 320.700 ;
        RECT 8.700 315.000 10.500 321.600 ;
        RECT 11.700 315.600 13.500 324.600 ;
        RECT 23.700 321.600 25.800 323.700 ;
        RECT 31.200 323.100 34.500 325.200 ;
        RECT 14.700 315.000 16.500 321.600 ;
        RECT 18.300 318.600 20.400 320.700 ;
        RECT 21.300 318.600 23.400 320.700 ;
        RECT 18.300 315.600 20.100 318.600 ;
        RECT 21.300 315.600 23.100 318.600 ;
        RECT 24.300 315.600 26.100 321.600 ;
        RECT 27.300 315.000 29.100 321.600 ;
        RECT 31.200 315.600 33.000 323.100 ;
        RECT 37.200 321.600 39.900 325.500 ;
        RECT 52.200 324.600 57.900 325.800 ;
        RECT 49.500 323.700 51.300 324.300 ;
        RECT 43.200 322.500 51.300 323.700 ;
        RECT 43.200 321.600 45.300 322.500 ;
        RECT 52.200 321.600 53.400 324.600 ;
        RECT 56.100 324.000 57.900 324.600 ;
        RECT 61.800 323.400 62.700 326.700 ;
        RECT 58.800 322.500 62.700 323.400 ;
        RECT 64.500 347.400 66.300 350.400 ;
        RECT 67.500 347.400 69.300 351.000 ;
        RECT 64.500 334.050 66.000 347.400 ;
        RECT 86.100 344.400 87.900 351.000 ;
        RECT 89.100 343.500 90.900 350.400 ;
        RECT 92.100 344.400 93.900 351.000 ;
        RECT 95.100 343.500 96.900 350.400 ;
        RECT 98.100 344.400 99.900 351.000 ;
        RECT 101.100 343.500 102.900 350.400 ;
        RECT 104.100 344.400 105.900 351.000 ;
        RECT 107.100 343.500 108.900 350.400 ;
        RECT 110.100 344.400 111.900 351.000 ;
        RECT 128.100 347.400 129.900 351.000 ;
        RECT 131.100 347.400 132.900 350.400 ;
        RECT 149.100 347.400 150.900 351.000 ;
        RECT 152.100 347.400 153.900 350.400 ;
        RECT 155.100 347.400 156.900 351.000 ;
        RECT 173.100 347.400 174.900 351.000 ;
        RECT 176.100 347.400 177.900 350.400 ;
        RECT 194.100 347.400 195.900 351.000 ;
        RECT 197.100 347.400 198.900 350.400 ;
        RECT 200.100 347.400 201.900 351.000 ;
        RECT 89.100 342.300 93.000 343.500 ;
        RECT 95.100 342.300 99.000 343.500 ;
        RECT 101.100 342.300 105.000 343.500 ;
        RECT 107.100 342.300 109.950 343.500 ;
        RECT 91.800 341.400 93.000 342.300 ;
        RECT 97.800 341.400 99.000 342.300 ;
        RECT 103.800 341.400 105.000 342.300 ;
        RECT 91.800 340.200 96.000 341.400 ;
        RECT 88.800 337.050 90.600 338.850 ;
        RECT 88.800 334.950 90.900 337.050 ;
        RECT 64.500 331.950 66.900 334.050 ;
        RECT 58.800 321.600 60.000 322.500 ;
        RECT 64.500 321.600 66.000 331.950 ;
        RECT 91.800 329.700 93.000 340.200 ;
        RECT 94.200 339.600 96.000 340.200 ;
        RECT 97.800 340.200 102.000 341.400 ;
        RECT 97.800 329.700 99.000 340.200 ;
        RECT 100.200 339.600 102.000 340.200 ;
        RECT 103.800 340.200 108.000 341.400 ;
        RECT 103.800 329.700 105.000 340.200 ;
        RECT 106.200 339.600 108.000 340.200 ;
        RECT 108.900 337.050 109.950 342.300 ;
        RECT 131.100 337.050 132.300 347.400 ;
        RECT 152.700 337.050 153.600 347.400 ;
        RECT 157.950 339.450 160.050 340.050 ;
        RECT 166.950 339.450 169.050 340.050 ;
        RECT 157.950 338.550 169.050 339.450 ;
        RECT 157.950 337.950 160.050 338.550 ;
        RECT 166.950 337.950 169.050 338.550 ;
        RECT 176.100 337.050 177.300 347.400 ;
        RECT 197.700 337.050 198.600 347.400 ;
        RECT 218.100 341.400 219.900 351.000 ;
        RECT 224.700 342.000 226.500 350.400 ;
        RECT 242.100 345.300 243.900 350.400 ;
        RECT 245.100 346.200 246.900 351.000 ;
        RECT 248.100 345.300 249.900 350.400 ;
        RECT 242.100 343.950 249.900 345.300 ;
        RECT 251.100 344.400 252.900 350.400 ;
        RECT 269.100 347.400 270.900 351.000 ;
        RECT 272.100 347.400 273.900 350.400 ;
        RECT 275.100 347.400 276.900 351.000 ;
        RECT 251.100 342.300 252.300 344.400 ;
        RECT 224.700 340.800 228.000 342.000 ;
        RECT 218.100 337.050 219.900 338.850 ;
        RECT 224.100 337.050 225.900 338.850 ;
        RECT 227.100 337.050 228.000 340.800 ;
        RECT 248.700 341.400 252.300 342.300 ;
        RECT 245.100 337.050 246.900 338.850 ;
        RECT 248.700 337.050 249.900 341.400 ;
        RECT 251.100 337.050 252.900 338.850 ;
        RECT 272.400 337.050 273.300 347.400 ;
        RECT 293.100 345.300 294.900 350.400 ;
        RECT 296.100 346.200 297.900 351.000 ;
        RECT 299.100 345.300 300.900 350.400 ;
        RECT 293.100 343.950 300.900 345.300 ;
        RECT 302.100 344.400 303.900 350.400 ;
        RECT 320.400 344.400 322.200 351.000 ;
        RECT 302.100 342.300 303.300 344.400 ;
        RECT 325.500 343.200 327.300 350.400 ;
        RECT 344.400 344.400 346.200 351.000 ;
        RECT 349.500 343.200 351.300 350.400 ;
        RECT 365.100 347.400 366.900 351.000 ;
        RECT 368.100 347.400 369.900 350.400 ;
        RECT 371.700 347.400 373.500 351.000 ;
        RECT 374.700 347.400 376.500 350.400 ;
        RECT 299.700 341.400 303.300 342.300 ;
        RECT 323.100 342.300 327.300 343.200 ;
        RECT 347.100 342.300 351.300 343.200 ;
        RECT 296.100 337.050 297.900 338.850 ;
        RECT 299.700 337.050 300.900 341.400 ;
        RECT 302.100 337.050 303.900 338.850 ;
        RECT 320.250 337.050 322.050 338.850 ;
        RECT 323.100 337.050 324.300 342.300 ;
        RECT 326.100 337.050 327.900 338.850 ;
        RECT 344.250 337.050 346.050 338.850 ;
        RECT 347.100 337.050 348.300 342.300 ;
        RECT 350.100 337.050 351.900 338.850 ;
        RECT 368.100 337.050 369.300 347.400 ;
        RECT 106.800 334.950 109.950 337.050 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 217.950 334.950 220.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 268.950 334.950 271.050 337.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 292.950 334.950 295.050 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 108.900 329.700 109.950 334.950 ;
        RECT 128.100 333.150 129.900 334.950 ;
        RECT 89.100 328.500 93.000 329.700 ;
        RECT 95.100 328.500 99.000 329.700 ;
        RECT 101.100 328.500 105.000 329.700 ;
        RECT 107.100 328.500 109.950 329.700 ;
        RECT 34.200 315.000 36.000 321.600 ;
        RECT 37.200 315.600 39.000 321.600 ;
        RECT 40.200 318.600 42.300 320.700 ;
        RECT 43.200 318.600 45.300 320.700 ;
        RECT 46.200 318.600 48.300 320.700 ;
        RECT 40.200 315.600 42.000 318.600 ;
        RECT 43.200 315.600 45.000 318.600 ;
        RECT 46.200 315.600 48.000 318.600 ;
        RECT 49.200 315.000 51.000 321.600 ;
        RECT 52.200 315.600 54.000 321.600 ;
        RECT 55.200 315.000 57.000 321.600 ;
        RECT 58.200 315.600 60.000 321.600 ;
        RECT 61.200 315.000 63.000 321.600 ;
        RECT 64.500 315.600 66.300 321.600 ;
        RECT 67.500 315.000 69.300 321.600 ;
        RECT 86.100 315.000 87.900 327.600 ;
        RECT 89.100 315.600 90.900 328.500 ;
        RECT 92.100 315.000 93.900 327.600 ;
        RECT 95.100 315.600 96.900 328.500 ;
        RECT 98.100 315.000 99.900 327.600 ;
        RECT 101.100 315.600 102.900 328.500 ;
        RECT 104.100 315.000 105.900 327.600 ;
        RECT 107.100 315.600 108.900 328.500 ;
        RECT 110.100 315.000 111.900 327.600 ;
        RECT 131.100 321.600 132.300 334.950 ;
        RECT 149.100 333.150 150.900 334.950 ;
        RECT 152.700 327.600 153.600 334.950 ;
        RECT 154.950 333.150 156.750 334.950 ;
        RECT 173.100 333.150 174.900 334.950 ;
        RECT 150.000 326.400 153.600 327.600 ;
        RECT 128.100 315.000 129.900 321.600 ;
        RECT 131.100 315.600 132.900 321.600 ;
        RECT 150.000 315.600 151.800 326.400 ;
        RECT 155.100 315.000 156.900 327.600 ;
        RECT 176.100 321.600 177.300 334.950 ;
        RECT 194.100 333.150 195.900 334.950 ;
        RECT 197.700 327.600 198.600 334.950 ;
        RECT 199.950 333.150 201.750 334.950 ;
        RECT 205.950 333.450 210.000 334.050 ;
        RECT 205.950 331.950 210.450 333.450 ;
        RECT 195.000 326.400 198.600 327.600 ;
        RECT 173.100 315.000 174.900 321.600 ;
        RECT 176.100 315.600 177.900 321.600 ;
        RECT 195.000 315.600 196.800 326.400 ;
        RECT 200.100 315.000 201.900 327.600 ;
        RECT 209.550 327.450 210.450 331.950 ;
        RECT 211.950 330.450 214.050 334.050 ;
        RECT 221.100 333.150 222.900 334.950 ;
        RECT 217.950 330.450 220.050 331.050 ;
        RECT 211.950 330.000 220.050 330.450 ;
        RECT 212.550 329.550 220.050 330.000 ;
        RECT 217.950 328.950 220.050 329.550 ;
        RECT 214.950 327.450 217.050 328.050 ;
        RECT 209.550 326.550 217.050 327.450 ;
        RECT 214.950 325.950 217.050 326.550 ;
        RECT 227.100 322.800 228.000 334.950 ;
        RECT 242.100 333.150 243.900 334.950 ;
        RECT 248.700 327.600 249.900 334.950 ;
        RECT 269.250 333.150 271.050 334.950 ;
        RECT 272.400 327.600 273.300 334.950 ;
        RECT 275.100 333.150 276.900 334.950 ;
        RECT 277.950 333.450 280.050 334.050 ;
        RECT 286.950 333.450 289.050 334.050 ;
        RECT 277.950 332.550 289.050 333.450 ;
        RECT 293.100 333.150 294.900 334.950 ;
        RECT 277.950 331.950 280.050 332.550 ;
        RECT 286.950 331.950 289.050 332.550 ;
        RECT 283.950 330.450 286.050 331.050 ;
        RECT 295.950 330.450 298.050 330.750 ;
        RECT 283.950 329.550 298.050 330.450 ;
        RECT 283.950 328.950 286.050 329.550 ;
        RECT 295.950 328.650 298.050 329.550 ;
        RECT 299.700 327.600 300.900 334.950 ;
        RECT 221.400 321.900 228.000 322.800 ;
        RECT 221.400 321.600 222.900 321.900 ;
        RECT 218.100 315.000 219.900 321.600 ;
        RECT 221.100 315.600 222.900 321.600 ;
        RECT 227.100 321.600 228.000 321.900 ;
        RECT 224.100 315.000 225.900 321.000 ;
        RECT 227.100 315.600 228.900 321.600 ;
        RECT 242.400 315.000 244.200 327.600 ;
        RECT 247.500 326.100 249.900 327.600 ;
        RECT 247.500 315.600 249.300 326.100 ;
        RECT 250.200 323.100 252.000 324.900 ;
        RECT 250.500 315.000 252.300 321.600 ;
        RECT 269.100 315.000 270.900 327.600 ;
        RECT 272.400 326.400 276.000 327.600 ;
        RECT 274.200 315.600 276.000 326.400 ;
        RECT 293.400 315.000 295.200 327.600 ;
        RECT 298.500 326.100 300.900 327.600 ;
        RECT 298.500 315.600 300.300 326.100 ;
        RECT 301.200 323.100 303.000 324.900 ;
        RECT 323.100 321.600 324.300 334.950 ;
        RECT 347.100 321.600 348.300 334.950 ;
        RECT 365.100 333.150 366.900 334.950 ;
        RECT 355.950 327.450 358.050 328.050 ;
        RECT 361.950 327.450 364.050 328.050 ;
        RECT 355.950 326.550 364.050 327.450 ;
        RECT 355.950 325.950 358.050 326.550 ;
        RECT 361.950 325.950 364.050 326.550 ;
        RECT 368.100 321.600 369.300 334.950 ;
        RECT 375.000 334.050 376.500 347.400 ;
        RECT 374.100 331.950 376.500 334.050 ;
        RECT 375.000 321.600 376.500 331.950 ;
        RECT 378.300 344.400 380.100 350.400 ;
        RECT 383.700 344.400 385.500 351.000 ;
        RECT 388.800 345.600 390.600 350.400 ;
        RECT 393.000 347.400 394.800 350.400 ;
        RECT 396.000 347.400 397.800 350.400 ;
        RECT 399.000 347.400 400.800 350.400 ;
        RECT 402.000 347.400 403.800 350.400 ;
        RECT 405.000 347.400 406.800 351.000 ;
        RECT 386.400 344.400 390.600 345.600 ;
        RECT 392.700 345.300 394.800 347.400 ;
        RECT 395.700 345.300 397.800 347.400 ;
        RECT 398.700 345.300 400.800 347.400 ;
        RECT 401.700 345.300 403.800 347.400 ;
        RECT 408.000 346.500 409.800 350.400 ;
        RECT 412.500 347.400 414.300 351.000 ;
        RECT 415.500 347.400 417.300 350.400 ;
        RECT 418.500 347.400 420.300 350.400 ;
        RECT 421.500 347.400 423.300 350.400 ;
        RECT 407.100 344.400 409.800 346.500 ;
        RECT 411.600 345.600 413.400 346.500 ;
        RECT 411.600 344.400 414.300 345.600 ;
        RECT 415.200 345.300 417.300 347.400 ;
        RECT 418.200 345.300 420.300 347.400 ;
        RECT 421.200 345.300 423.300 347.400 ;
        RECT 425.700 344.400 427.500 350.400 ;
        RECT 431.100 344.400 432.900 351.000 ;
        RECT 436.500 344.400 438.300 350.400 ;
        RECT 455.100 349.500 462.900 350.400 ;
        RECT 455.100 344.400 456.900 349.500 ;
        RECT 458.100 344.400 459.900 348.600 ;
        RECT 461.100 345.000 462.900 349.500 ;
        RECT 464.100 345.900 465.900 351.000 ;
        RECT 467.100 345.000 468.900 350.400 ;
        RECT 378.300 327.600 379.200 344.400 ;
        RECT 386.400 341.100 387.900 344.400 ;
        RECT 392.100 342.600 398.700 344.400 ;
        RECT 413.400 343.800 414.300 344.400 ;
        RECT 416.400 343.800 418.200 344.400 ;
        RECT 413.400 342.600 420.600 343.800 ;
        RECT 380.100 339.300 387.900 341.100 ;
        RECT 404.100 340.500 405.900 342.300 ;
        RECT 403.800 339.900 405.900 340.500 ;
        RECT 388.800 338.400 405.900 339.900 ;
        RECT 410.100 339.900 412.200 340.050 ;
        RECT 413.400 339.900 415.200 340.800 ;
        RECT 410.100 339.000 415.200 339.900 ;
        RECT 419.700 339.600 420.600 342.600 ;
        RECT 425.700 343.500 427.200 344.400 ;
        RECT 425.700 342.300 434.100 343.500 ;
        RECT 432.300 341.700 434.100 342.300 ;
        RECT 421.500 340.800 423.600 341.700 ;
        RECT 437.100 340.800 438.300 344.400 ;
        RECT 458.700 342.900 459.600 344.400 ;
        RECT 461.100 344.100 468.900 345.000 ;
        RECT 485.100 345.300 486.900 350.400 ;
        RECT 488.100 346.200 489.900 351.000 ;
        RECT 491.100 345.300 492.900 350.400 ;
        RECT 485.100 343.950 492.900 345.300 ;
        RECT 494.100 344.400 495.900 350.400 ;
        RECT 513.000 344.400 514.800 351.000 ;
        RECT 517.500 345.600 519.300 350.400 ;
        RECT 520.500 347.400 522.300 351.000 ;
        RECT 539.100 347.400 540.900 351.000 ;
        RECT 542.100 347.400 543.900 350.400 ;
        RECT 517.500 344.400 522.600 345.600 ;
        RECT 458.700 341.700 463.050 342.900 ;
        RECT 494.100 342.300 495.300 344.400 ;
        RECT 421.500 339.600 438.300 340.800 ;
        RECT 383.700 336.900 390.300 338.400 ;
        RECT 410.100 337.950 412.200 339.000 ;
        RECT 418.800 337.800 420.600 339.600 ;
        RECT 383.700 334.050 385.200 336.900 ;
        RECT 391.500 335.700 435.900 336.900 ;
        RECT 391.500 334.200 392.400 335.700 ;
        RECT 383.100 331.950 385.200 334.050 ;
        RECT 387.300 332.400 392.400 334.200 ;
        RECT 395.100 333.900 408.600 334.800 ;
        RECT 415.800 333.900 417.600 334.500 ;
        RECT 434.100 334.050 435.900 335.700 ;
        RECT 395.100 332.700 396.000 333.900 ;
        RECT 395.100 330.900 396.900 332.700 ;
        RECT 401.100 331.200 405.000 333.000 ;
        RECT 406.500 332.700 417.600 333.900 ;
        RECT 428.100 333.750 430.200 334.050 ;
        RECT 406.500 331.800 408.600 332.700 ;
        RECT 426.300 331.950 430.200 333.750 ;
        RECT 434.100 331.950 436.200 334.050 ;
        RECT 426.300 331.200 428.100 331.950 ;
        RECT 401.100 330.900 403.200 331.200 ;
        RECT 414.600 330.300 428.100 331.200 ;
        RECT 380.100 329.700 381.900 330.300 ;
        RECT 414.600 329.700 415.800 330.300 ;
        RECT 380.100 328.500 415.800 329.700 ;
        RECT 418.500 328.500 420.600 328.800 ;
        RECT 378.300 326.700 394.800 327.600 ;
        RECT 378.300 323.400 379.200 326.700 ;
        RECT 383.100 324.600 388.800 325.800 ;
        RECT 392.700 325.500 394.800 326.700 ;
        RECT 398.100 326.400 415.800 327.600 ;
        RECT 418.500 327.300 430.500 328.500 ;
        RECT 418.500 326.700 420.600 327.300 ;
        RECT 428.700 326.700 430.500 327.300 ;
        RECT 398.100 325.500 400.200 326.400 ;
        RECT 414.600 325.800 415.800 326.400 ;
        RECT 432.000 325.800 433.800 326.100 ;
        RECT 383.100 324.000 384.900 324.600 ;
        RECT 378.300 322.500 382.200 323.400 ;
        RECT 381.000 321.600 382.200 322.500 ;
        RECT 387.600 321.600 388.800 324.600 ;
        RECT 389.700 323.700 391.500 324.300 ;
        RECT 389.700 322.500 397.800 323.700 ;
        RECT 395.700 321.600 397.800 322.500 ;
        RECT 401.100 321.600 403.800 325.500 ;
        RECT 406.500 323.100 409.800 325.200 ;
        RECT 414.600 324.600 433.800 325.800 ;
        RECT 301.500 315.000 303.300 321.600 ;
        RECT 320.100 315.000 321.900 321.600 ;
        RECT 323.100 315.600 324.900 321.600 ;
        RECT 326.100 315.000 327.900 321.600 ;
        RECT 344.100 315.000 345.900 321.600 ;
        RECT 347.100 315.600 348.900 321.600 ;
        RECT 350.100 315.000 351.900 321.600 ;
        RECT 365.100 315.000 366.900 321.600 ;
        RECT 368.100 315.600 369.900 321.600 ;
        RECT 371.700 315.000 373.500 321.600 ;
        RECT 374.700 315.600 376.500 321.600 ;
        RECT 378.000 315.000 379.800 321.600 ;
        RECT 381.000 315.600 382.800 321.600 ;
        RECT 384.000 315.000 385.800 321.600 ;
        RECT 387.000 315.600 388.800 321.600 ;
        RECT 390.000 315.000 391.800 321.600 ;
        RECT 392.700 318.600 394.800 320.700 ;
        RECT 395.700 318.600 397.800 320.700 ;
        RECT 398.700 318.600 400.800 320.700 ;
        RECT 393.000 315.600 394.800 318.600 ;
        RECT 396.000 315.600 397.800 318.600 ;
        RECT 399.000 315.600 400.800 318.600 ;
        RECT 402.000 315.600 403.800 321.600 ;
        RECT 405.000 315.000 406.800 321.600 ;
        RECT 408.000 315.600 409.800 323.100 ;
        RECT 415.200 321.600 417.300 323.700 ;
        RECT 411.900 315.000 413.700 321.600 ;
        RECT 414.900 315.600 416.700 321.600 ;
        RECT 417.600 318.600 419.700 320.700 ;
        RECT 420.600 318.600 422.700 320.700 ;
        RECT 417.900 315.600 419.700 318.600 ;
        RECT 420.900 315.600 422.700 318.600 ;
        RECT 424.500 315.000 426.300 321.600 ;
        RECT 427.500 315.600 429.300 324.600 ;
        RECT 432.000 324.300 433.800 324.600 ;
        RECT 437.100 323.400 438.300 339.600 ;
        RECT 458.250 337.050 460.050 338.850 ;
        RECT 462.000 337.050 463.050 341.700 ;
        RECT 491.700 341.400 495.300 342.300 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 463.950 337.050 465.750 338.850 ;
        RECT 488.100 337.050 489.900 338.850 ;
        RECT 491.700 337.050 492.900 341.400 ;
        RECT 494.100 337.050 495.900 338.850 ;
        RECT 512.100 337.050 513.900 338.850 ;
        RECT 518.250 337.050 520.050 338.850 ;
        RECT 521.700 337.050 522.600 344.400 ;
        RECT 542.100 337.050 543.300 347.400 ;
        RECT 560.100 341.400 561.900 351.000 ;
        RECT 566.700 342.000 568.500 350.400 ;
        RECT 587.100 344.400 588.900 350.400 ;
        RECT 587.700 342.300 588.900 344.400 ;
        RECT 590.100 345.300 591.900 350.400 ;
        RECT 593.100 346.200 594.900 351.000 ;
        RECT 596.100 345.300 597.900 350.400 ;
        RECT 590.100 343.950 597.900 345.300 ;
        RECT 614.100 344.400 615.900 350.400 ;
        RECT 614.700 342.300 615.900 344.400 ;
        RECT 617.100 345.300 618.900 350.400 ;
        RECT 620.100 346.200 621.900 351.000 ;
        RECT 623.100 345.300 624.900 350.400 ;
        RECT 617.100 343.950 624.900 345.300 ;
        RECT 641.100 344.400 642.900 350.400 ;
        RECT 644.100 345.300 645.900 351.000 ;
        RECT 648.300 345.000 650.100 350.400 ;
        RECT 652.800 345.300 654.600 351.000 ;
        RECT 641.100 343.500 642.600 344.400 ;
        RECT 566.700 340.800 570.000 342.000 ;
        RECT 587.700 341.400 591.300 342.300 ;
        RECT 614.700 341.400 618.300 342.300 ;
        RECT 641.100 342.000 645.600 343.500 ;
        RECT 643.500 341.400 645.600 342.000 ;
        RECT 649.200 342.900 650.100 345.000 ;
        RECT 656.100 344.400 657.900 350.400 ;
        RECT 653.400 343.500 657.900 344.400 ;
        RECT 674.100 345.300 675.900 350.400 ;
        RECT 677.100 346.200 678.900 351.000 ;
        RECT 680.100 345.300 681.900 350.400 ;
        RECT 674.100 343.950 681.900 345.300 ;
        RECT 683.100 344.400 684.900 350.400 ;
        RECT 701.100 344.400 702.900 350.400 ;
        RECT 704.400 345.300 706.200 351.000 ;
        RECT 708.900 345.000 710.700 350.400 ;
        RECT 713.100 345.300 714.900 351.000 ;
        RECT 560.100 337.050 561.900 338.850 ;
        RECT 566.100 337.050 567.900 338.850 ;
        RECT 569.100 337.050 570.000 340.800 ;
        RECT 587.100 337.050 588.900 338.850 ;
        RECT 590.100 337.050 591.300 341.400 ;
        RECT 593.100 337.050 594.900 338.850 ;
        RECT 614.100 337.050 615.900 338.850 ;
        RECT 617.100 337.050 618.300 341.400 ;
        RECT 646.500 339.900 648.300 341.700 ;
        RECT 649.200 340.800 652.200 342.900 ;
        RECT 653.400 341.100 655.500 343.500 ;
        RECT 683.100 342.300 684.300 344.400 ;
        RECT 701.100 343.500 705.600 344.400 ;
        RECT 680.700 341.400 684.300 342.300 ;
        RECT 645.900 339.000 648.000 339.900 ;
        RECT 620.100 337.050 621.900 338.850 ;
        RECT 641.400 337.800 648.000 339.000 ;
        RECT 641.400 337.200 643.200 337.800 ;
        RECT 463.950 334.950 466.050 337.050 ;
        RECT 466.950 334.950 469.050 337.050 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 487.950 334.950 490.050 337.050 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 511.950 334.950 514.050 337.050 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 641.100 334.950 643.200 337.200 ;
        RECT 455.250 333.150 457.050 334.950 ;
        RECT 462.000 327.600 463.050 334.950 ;
        RECT 467.100 333.150 468.900 334.950 ;
        RECT 485.100 333.150 486.900 334.950 ;
        RECT 491.700 327.600 492.900 334.950 ;
        RECT 515.250 333.150 517.050 334.950 ;
        RECT 521.700 327.600 522.600 334.950 ;
        RECT 539.100 333.150 540.900 334.950 ;
        RECT 434.700 322.500 438.300 323.400 ;
        RECT 434.700 321.600 435.600 322.500 ;
        RECT 430.500 315.000 432.300 321.600 ;
        RECT 433.500 320.700 435.600 321.600 ;
        RECT 433.500 315.600 435.300 320.700 ;
        RECT 436.500 315.000 438.300 321.600 ;
        RECT 456.600 315.000 458.400 327.600 ;
        RECT 461.100 315.600 464.400 327.600 ;
        RECT 467.100 315.000 468.900 327.600 ;
        RECT 485.400 315.000 487.200 327.600 ;
        RECT 490.500 326.100 492.900 327.600 ;
        RECT 512.100 326.700 519.900 327.600 ;
        RECT 490.500 315.600 492.300 326.100 ;
        RECT 493.200 323.100 495.000 324.900 ;
        RECT 493.500 315.000 495.300 321.600 ;
        RECT 512.100 315.600 513.900 326.700 ;
        RECT 515.100 315.000 516.900 325.800 ;
        RECT 518.100 315.600 519.900 326.700 ;
        RECT 521.100 315.600 522.900 327.600 ;
        RECT 542.100 321.600 543.300 334.950 ;
        RECT 563.100 333.150 564.900 334.950 ;
        RECT 569.100 322.800 570.000 334.950 ;
        RECT 590.100 327.600 591.300 334.950 ;
        RECT 596.100 333.150 597.900 334.950 ;
        RECT 617.100 327.600 618.300 334.950 ;
        RECT 623.100 333.150 624.900 334.950 ;
        RECT 645.900 334.800 648.000 336.900 ;
        RECT 645.900 333.000 647.700 334.800 ;
        RECT 649.200 334.050 650.100 340.800 ;
        RECT 651.000 336.900 653.100 339.000 ;
        RECT 677.100 337.050 678.900 338.850 ;
        RECT 680.700 337.050 681.900 341.400 ;
        RECT 703.500 341.100 705.600 343.500 ;
        RECT 708.900 342.900 709.800 345.000 ;
        RECT 716.100 344.400 717.900 350.400 ;
        RECT 721.950 348.450 724.050 349.050 ;
        RECT 730.950 348.450 733.050 349.050 ;
        RECT 721.950 347.550 733.050 348.450 ;
        RECT 721.950 346.950 724.050 347.550 ;
        RECT 730.950 346.950 733.050 347.550 ;
        RECT 734.700 347.400 736.500 351.000 ;
        RECT 737.700 345.600 739.500 350.400 ;
        RECT 716.400 343.500 717.900 344.400 ;
        RECT 706.800 340.800 709.800 342.900 ;
        RECT 713.400 342.000 717.900 343.500 ;
        RECT 734.400 344.400 739.500 345.600 ;
        RECT 742.200 344.400 744.000 351.000 ;
        RECT 761.100 344.400 762.900 350.400 ;
        RECT 718.950 342.450 721.050 343.050 ;
        RECT 730.950 342.450 733.050 343.050 ;
        RECT 683.100 337.050 684.900 338.850 ;
        RECT 651.000 335.100 652.800 336.900 ;
        RECT 655.800 334.950 657.900 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 679.950 334.950 682.050 337.050 ;
        RECT 682.950 334.950 685.050 337.050 ;
        RECT 701.100 334.950 703.200 337.050 ;
        RECT 705.900 336.900 708.000 339.000 ;
        RECT 706.200 335.100 708.000 336.900 ;
        RECT 649.200 332.700 652.200 334.050 ;
        RECT 655.800 333.150 657.600 334.950 ;
        RECT 674.100 333.150 675.900 334.950 ;
        RECT 650.100 331.950 652.200 332.700 ;
        RECT 647.400 329.700 649.200 331.500 ;
        RECT 643.800 328.800 649.200 329.700 ;
        RECT 643.800 327.900 645.900 328.800 ;
        RECT 590.100 326.100 592.500 327.600 ;
        RECT 588.000 323.100 589.800 324.900 ;
        RECT 563.400 321.900 570.000 322.800 ;
        RECT 563.400 321.600 564.900 321.900 ;
        RECT 539.100 315.000 540.900 321.600 ;
        RECT 542.100 315.600 543.900 321.600 ;
        RECT 560.100 315.000 561.900 321.600 ;
        RECT 563.100 315.600 564.900 321.600 ;
        RECT 569.100 321.600 570.000 321.900 ;
        RECT 566.100 315.000 567.900 321.000 ;
        RECT 569.100 315.600 570.900 321.600 ;
        RECT 587.700 315.000 589.500 321.600 ;
        RECT 590.700 315.600 592.500 326.100 ;
        RECT 595.800 315.000 597.600 327.600 ;
        RECT 617.100 326.100 619.500 327.600 ;
        RECT 615.000 323.100 616.800 324.900 ;
        RECT 614.700 315.000 616.500 321.600 ;
        RECT 617.700 315.600 619.500 326.100 ;
        RECT 622.800 315.000 624.600 327.600 ;
        RECT 641.100 326.700 645.900 327.900 ;
        RECT 650.700 327.600 651.900 331.950 ;
        RECT 648.600 326.700 651.900 327.600 ;
        RECT 652.800 327.600 654.900 328.500 ;
        RECT 680.700 327.600 681.900 334.950 ;
        RECT 701.400 333.150 703.200 334.950 ;
        RECT 708.900 334.050 709.800 340.800 ;
        RECT 710.700 339.900 712.500 341.700 ;
        RECT 713.400 341.400 715.500 342.000 ;
        RECT 718.950 341.550 733.050 342.450 ;
        RECT 718.950 340.950 721.050 341.550 ;
        RECT 730.950 340.950 733.050 341.550 ;
        RECT 711.000 339.000 713.100 339.900 ;
        RECT 711.000 337.800 717.600 339.000 ;
        RECT 715.800 337.200 717.600 337.800 ;
        RECT 711.000 334.800 713.100 336.900 ;
        RECT 715.800 334.950 717.900 337.200 ;
        RECT 734.400 337.050 735.300 344.400 ;
        RECT 761.700 342.300 762.900 344.400 ;
        RECT 764.100 345.300 765.900 350.400 ;
        RECT 767.100 346.200 768.900 351.000 ;
        RECT 770.100 345.300 771.900 350.400 ;
        RECT 764.100 343.950 771.900 345.300 ;
        RECT 788.100 345.300 789.900 350.400 ;
        RECT 791.100 346.200 792.900 351.000 ;
        RECT 794.100 345.300 795.900 350.400 ;
        RECT 788.100 343.950 795.900 345.300 ;
        RECT 797.100 344.400 798.900 350.400 ;
        RECT 815.100 344.400 816.900 350.400 ;
        RECT 818.100 344.400 819.900 351.000 ;
        RECT 821.100 347.400 822.900 350.400 ;
        RECT 797.100 342.300 798.300 344.400 ;
        RECT 761.700 341.400 765.300 342.300 ;
        RECT 736.950 337.050 738.750 338.850 ;
        RECT 743.100 337.050 744.900 338.850 ;
        RECT 761.100 337.050 762.900 338.850 ;
        RECT 764.100 337.050 765.300 341.400 ;
        RECT 794.700 341.400 798.300 342.300 ;
        RECT 772.950 339.450 775.050 340.050 ;
        RECT 781.950 339.450 784.050 340.050 ;
        RECT 767.100 337.050 768.900 338.850 ;
        RECT 772.950 338.550 784.050 339.450 ;
        RECT 772.950 337.950 775.050 338.550 ;
        RECT 781.950 337.950 784.050 338.550 ;
        RECT 791.100 337.050 792.900 338.850 ;
        RECT 794.700 337.050 795.900 341.400 ;
        RECT 797.100 337.050 798.900 338.850 ;
        RECT 815.100 337.050 816.300 344.400 ;
        RECT 821.700 343.500 822.900 347.400 ;
        RECT 817.200 342.600 822.900 343.500 ;
        RECT 817.200 341.700 819.000 342.600 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 815.100 334.950 817.200 337.050 ;
        RECT 706.800 332.700 709.800 334.050 ;
        RECT 711.300 333.000 713.100 334.800 ;
        RECT 706.800 331.950 708.900 332.700 ;
        RECT 704.100 327.600 706.200 328.500 ;
        RECT 641.100 315.600 642.900 326.700 ;
        RECT 644.100 315.000 645.900 325.500 ;
        RECT 648.600 315.600 650.400 326.700 ;
        RECT 652.800 326.400 657.900 327.600 ;
        RECT 652.800 315.000 654.900 325.500 ;
        RECT 656.100 315.600 657.900 326.400 ;
        RECT 674.400 315.000 676.200 327.600 ;
        RECT 679.500 326.100 681.900 327.600 ;
        RECT 701.100 326.400 706.200 327.600 ;
        RECT 707.100 327.600 708.300 331.950 ;
        RECT 709.800 329.700 711.600 331.500 ;
        RECT 709.800 328.800 715.200 329.700 ;
        RECT 713.100 327.900 715.200 328.800 ;
        RECT 707.100 326.700 710.400 327.600 ;
        RECT 713.100 326.700 717.900 327.900 ;
        RECT 734.400 327.600 735.300 334.950 ;
        RECT 739.950 333.150 741.750 334.950 ;
        RECT 764.100 327.600 765.300 334.950 ;
        RECT 770.100 333.150 771.900 334.950 ;
        RECT 788.100 333.150 789.900 334.950 ;
        RECT 794.700 327.600 795.900 334.950 ;
        RECT 679.500 315.600 681.300 326.100 ;
        RECT 682.200 323.100 684.000 324.900 ;
        RECT 682.500 315.000 684.300 321.600 ;
        RECT 701.100 315.600 702.900 326.400 ;
        RECT 704.100 315.000 706.200 325.500 ;
        RECT 708.600 315.600 710.400 326.700 ;
        RECT 713.100 315.000 714.900 325.500 ;
        RECT 716.100 315.600 717.900 326.700 ;
        RECT 734.100 315.600 735.900 327.600 ;
        RECT 737.100 326.700 744.900 327.600 ;
        RECT 737.100 315.600 738.900 326.700 ;
        RECT 740.100 315.000 741.900 325.800 ;
        RECT 743.100 315.600 744.900 326.700 ;
        RECT 764.100 326.100 766.500 327.600 ;
        RECT 745.950 324.450 748.050 325.050 ;
        RECT 751.950 324.450 754.050 325.050 ;
        RECT 745.950 323.550 754.050 324.450 ;
        RECT 745.950 322.950 748.050 323.550 ;
        RECT 751.950 322.950 754.050 323.550 ;
        RECT 762.000 323.100 763.800 324.900 ;
        RECT 751.950 321.450 754.050 321.900 ;
        RECT 757.950 321.450 760.050 322.050 ;
        RECT 751.950 320.550 760.050 321.450 ;
        RECT 751.950 319.800 754.050 320.550 ;
        RECT 757.950 319.950 760.050 320.550 ;
        RECT 761.700 315.000 763.500 321.600 ;
        RECT 764.700 315.600 766.500 326.100 ;
        RECT 769.800 315.000 771.600 327.600 ;
        RECT 788.400 315.000 790.200 327.600 ;
        RECT 793.500 326.100 795.900 327.600 ;
        RECT 815.100 327.600 816.300 334.950 ;
        RECT 818.100 330.300 819.000 341.700 ;
        RECT 839.100 341.400 840.900 351.000 ;
        RECT 845.700 342.000 847.500 350.400 ;
        RECT 866.100 345.300 867.900 350.400 ;
        RECT 869.100 346.200 870.900 351.000 ;
        RECT 872.100 345.300 873.900 350.400 ;
        RECT 866.100 343.950 873.900 345.300 ;
        RECT 875.100 344.400 876.900 350.400 ;
        RECT 893.700 347.400 895.500 351.000 ;
        RECT 896.700 345.600 898.500 350.400 ;
        RECT 893.400 344.400 898.500 345.600 ;
        RECT 901.200 344.400 903.000 351.000 ;
        RECT 875.100 342.300 876.300 344.400 ;
        RECT 845.700 340.800 849.000 342.000 ;
        RECT 839.100 337.050 840.900 338.850 ;
        RECT 845.100 337.050 846.900 338.850 ;
        RECT 848.100 337.050 849.000 340.800 ;
        RECT 872.700 341.400 876.300 342.300 ;
        RECT 869.100 337.050 870.900 338.850 ;
        RECT 872.700 337.050 873.900 341.400 ;
        RECT 875.100 337.050 876.900 338.850 ;
        RECT 893.400 337.050 894.300 344.400 ;
        RECT 922.500 342.000 924.300 350.400 ;
        RECT 921.000 340.800 924.300 342.000 ;
        RECT 929.100 341.400 930.900 351.000 ;
        RECT 947.100 341.400 948.900 351.000 ;
        RECT 953.700 342.000 955.500 350.400 ;
        RECT 974.100 347.400 975.900 351.000 ;
        RECT 977.100 347.400 978.900 350.400 ;
        RECT 980.100 347.400 981.900 351.000 ;
        RECT 958.950 342.450 961.050 343.050 ;
        RECT 973.950 342.450 976.050 343.050 ;
        RECT 953.700 340.800 957.000 342.000 ;
        RECT 958.950 341.550 976.050 342.450 ;
        RECT 958.950 340.950 961.050 341.550 ;
        RECT 973.950 340.950 976.050 341.550 ;
        RECT 916.950 339.450 919.050 340.050 ;
        RECT 895.950 337.050 897.750 338.850 ;
        RECT 902.100 337.050 903.900 338.850 ;
        RECT 908.550 338.550 919.050 339.450 ;
        RECT 820.500 334.950 822.600 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 865.950 334.950 868.050 337.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 820.800 333.150 822.600 334.950 ;
        RECT 842.100 333.150 843.900 334.950 ;
        RECT 817.200 329.400 819.000 330.300 ;
        RECT 817.200 328.500 822.900 329.400 ;
        RECT 793.500 315.600 795.300 326.100 ;
        RECT 796.200 323.100 798.000 324.900 ;
        RECT 796.500 315.000 798.300 321.600 ;
        RECT 815.100 315.600 816.900 327.600 ;
        RECT 818.100 315.000 819.900 325.800 ;
        RECT 821.700 321.600 822.900 328.500 ;
        RECT 848.100 322.800 849.000 334.950 ;
        RECT 866.100 333.150 867.900 334.950 ;
        RECT 859.950 330.450 862.050 331.050 ;
        RECT 868.950 330.450 871.050 331.050 ;
        RECT 859.950 329.550 871.050 330.450 ;
        RECT 859.950 328.950 862.050 329.550 ;
        RECT 868.950 328.950 871.050 329.550 ;
        RECT 872.700 327.600 873.900 334.950 ;
        RECT 893.400 327.600 894.300 334.950 ;
        RECT 898.950 333.150 900.750 334.950 ;
        RECT 908.550 333.450 909.450 338.550 ;
        RECT 916.950 337.950 919.050 338.550 ;
        RECT 921.000 337.050 921.900 340.800 ;
        RECT 923.100 337.050 924.900 338.850 ;
        RECT 929.100 337.050 930.900 338.850 ;
        RECT 947.100 337.050 948.900 338.850 ;
        RECT 953.100 337.050 954.900 338.850 ;
        RECT 956.100 337.050 957.000 340.800 ;
        RECT 977.400 337.050 978.300 347.400 ;
        RECT 998.100 345.300 999.900 350.400 ;
        RECT 1001.100 346.200 1002.900 351.000 ;
        RECT 1004.100 345.300 1005.900 350.400 ;
        RECT 998.100 343.950 1005.900 345.300 ;
        RECT 1007.100 344.400 1008.900 350.400 ;
        RECT 1025.100 347.400 1026.900 351.000 ;
        RECT 1028.100 347.400 1029.900 350.400 ;
        RECT 1007.100 342.300 1008.300 344.400 ;
        RECT 1004.700 341.400 1008.300 342.300 ;
        RECT 1001.100 337.050 1002.900 338.850 ;
        RECT 1004.700 337.050 1005.900 341.400 ;
        RECT 1007.100 337.050 1008.900 338.850 ;
        RECT 1028.100 337.050 1029.300 347.400 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 928.950 334.950 931.050 337.050 ;
        RECT 946.950 334.950 949.050 337.050 ;
        RECT 949.950 334.950 952.050 337.050 ;
        RECT 952.950 334.950 955.050 337.050 ;
        RECT 955.950 334.950 958.050 337.050 ;
        RECT 973.950 334.950 976.050 337.050 ;
        RECT 976.950 334.950 979.050 337.050 ;
        RECT 979.950 334.950 982.050 337.050 ;
        RECT 997.950 334.950 1000.050 337.050 ;
        RECT 1000.950 334.950 1003.050 337.050 ;
        RECT 1003.950 334.950 1006.050 337.050 ;
        RECT 1006.950 334.950 1009.050 337.050 ;
        RECT 1024.950 334.950 1027.050 337.050 ;
        RECT 1027.950 334.950 1030.050 337.050 ;
        RECT 905.550 332.550 909.450 333.450 ;
        RECT 898.950 330.450 901.050 331.050 ;
        RECT 905.550 330.450 906.450 332.550 ;
        RECT 898.950 329.550 906.450 330.450 ;
        RECT 898.950 328.950 901.050 329.550 ;
        RECT 842.400 321.900 849.000 322.800 ;
        RECT 842.400 321.600 843.900 321.900 ;
        RECT 821.100 315.600 822.900 321.600 ;
        RECT 823.950 318.450 826.050 319.050 ;
        RECT 835.950 318.450 838.050 319.050 ;
        RECT 823.950 317.550 838.050 318.450 ;
        RECT 823.950 316.950 826.050 317.550 ;
        RECT 835.950 316.950 838.050 317.550 ;
        RECT 839.100 315.000 840.900 321.600 ;
        RECT 842.100 315.600 843.900 321.600 ;
        RECT 848.100 321.600 849.000 321.900 ;
        RECT 845.100 315.000 846.900 321.000 ;
        RECT 848.100 315.600 849.900 321.600 ;
        RECT 866.400 315.000 868.200 327.600 ;
        RECT 871.500 326.100 873.900 327.600 ;
        RECT 871.500 315.600 873.300 326.100 ;
        RECT 874.200 323.100 876.000 324.900 ;
        RECT 874.500 315.000 876.300 321.600 ;
        RECT 893.100 315.600 894.900 327.600 ;
        RECT 896.100 326.700 903.900 327.600 ;
        RECT 896.100 315.600 897.900 326.700 ;
        RECT 899.100 315.000 900.900 325.800 ;
        RECT 902.100 315.600 903.900 326.700 ;
        RECT 921.000 322.800 921.900 334.950 ;
        RECT 926.100 333.150 927.900 334.950 ;
        RECT 950.100 333.150 951.900 334.950 ;
        RECT 928.950 330.450 931.050 331.050 ;
        RECT 940.950 330.450 943.050 331.050 ;
        RECT 952.950 330.450 955.050 331.050 ;
        RECT 928.950 329.550 955.050 330.450 ;
        RECT 928.950 328.950 931.050 329.550 ;
        RECT 940.950 328.950 943.050 329.550 ;
        RECT 952.950 328.950 955.050 329.550 ;
        RECT 956.100 322.800 957.000 334.950 ;
        RECT 974.250 333.150 976.050 334.950 ;
        RECT 977.400 327.600 978.300 334.950 ;
        RECT 980.100 333.150 981.900 334.950 ;
        RECT 998.100 333.150 999.900 334.950 ;
        RECT 1004.700 327.600 1005.900 334.950 ;
        RECT 1025.100 333.150 1026.900 334.950 ;
        RECT 921.000 321.900 927.600 322.800 ;
        RECT 921.000 321.600 921.900 321.900 ;
        RECT 920.100 315.600 921.900 321.600 ;
        RECT 926.100 321.600 927.600 321.900 ;
        RECT 950.400 321.900 957.000 322.800 ;
        RECT 950.400 321.600 951.900 321.900 ;
        RECT 923.100 315.000 924.900 321.000 ;
        RECT 926.100 315.600 927.900 321.600 ;
        RECT 929.100 315.000 930.900 321.600 ;
        RECT 947.100 315.000 948.900 321.600 ;
        RECT 950.100 315.600 951.900 321.600 ;
        RECT 956.100 321.600 957.000 321.900 ;
        RECT 953.100 315.000 954.900 321.000 ;
        RECT 956.100 315.600 957.900 321.600 ;
        RECT 974.100 315.000 975.900 327.600 ;
        RECT 977.400 326.400 981.000 327.600 ;
        RECT 979.200 315.600 981.000 326.400 ;
        RECT 998.400 315.000 1000.200 327.600 ;
        RECT 1003.500 326.100 1005.900 327.600 ;
        RECT 1003.500 315.600 1005.300 326.100 ;
        RECT 1006.200 323.100 1008.000 324.900 ;
        RECT 1028.100 321.600 1029.300 334.950 ;
        RECT 1006.500 315.000 1008.300 321.600 ;
        RECT 1025.100 315.000 1026.900 321.600 ;
        RECT 1028.100 315.600 1029.900 321.600 ;
        RECT 17.100 300.300 18.900 311.400 ;
        RECT 20.100 301.200 21.900 312.000 ;
        RECT 23.100 300.300 24.900 311.400 ;
        RECT 17.100 299.400 24.900 300.300 ;
        RECT 26.100 299.400 27.900 311.400 ;
        RECT 44.100 300.300 45.900 311.400 ;
        RECT 47.100 301.200 48.900 312.000 ;
        RECT 50.100 300.300 51.900 311.400 ;
        RECT 44.100 299.400 51.900 300.300 ;
        RECT 53.100 299.400 54.900 311.400 ;
        RECT 71.100 305.400 72.900 312.000 ;
        RECT 74.100 305.400 75.900 311.400 ;
        RECT 77.100 305.400 78.900 312.000 ;
        RECT 95.100 310.500 102.900 311.400 ;
        RECT 20.250 292.050 22.050 293.850 ;
        RECT 26.700 292.050 27.600 299.400 ;
        RECT 47.250 292.050 49.050 293.850 ;
        RECT 53.700 292.050 54.600 299.400 ;
        RECT 74.700 292.050 75.900 305.400 ;
        RECT 95.100 299.400 96.900 310.500 ;
        RECT 98.100 298.500 99.900 309.600 ;
        RECT 101.100 300.600 102.900 310.500 ;
        RECT 104.100 301.500 105.900 312.000 ;
        RECT 107.100 300.600 108.900 311.400 ;
        RECT 125.700 305.400 127.500 312.000 ;
        RECT 126.000 302.100 127.800 303.900 ;
        RECT 128.700 300.900 130.500 311.400 ;
        RECT 101.100 299.700 108.900 300.600 ;
        RECT 128.100 299.400 130.500 300.900 ;
        RECT 133.800 299.400 135.600 312.000 ;
        RECT 153.000 300.600 154.800 311.400 ;
        RECT 153.000 299.400 156.600 300.600 ;
        RECT 158.100 299.400 159.900 312.000 ;
        RECT 176.100 299.400 177.900 311.400 ;
        RECT 179.100 300.300 180.900 311.400 ;
        RECT 182.100 301.200 183.900 312.000 ;
        RECT 185.100 300.300 186.900 311.400 ;
        RECT 179.100 299.400 186.900 300.300 ;
        RECT 204.000 300.600 205.800 311.400 ;
        RECT 204.000 299.400 207.600 300.600 ;
        RECT 209.100 299.400 210.900 312.000 ;
        RECT 227.700 305.400 229.500 312.000 ;
        RECT 228.000 302.100 229.800 303.900 ;
        RECT 230.700 300.900 232.500 311.400 ;
        RECT 230.100 299.400 232.500 300.900 ;
        RECT 235.800 299.400 237.600 312.000 ;
        RECT 254.100 305.400 255.900 312.000 ;
        RECT 257.100 305.400 258.900 311.400 ;
        RECT 260.100 305.400 261.900 312.000 ;
        RECT 98.100 297.600 102.900 298.500 ;
        RECT 98.100 292.050 99.900 293.850 ;
        RECT 102.000 292.050 102.900 297.600 ;
        RECT 103.950 292.050 105.750 293.850 ;
        RECT 128.100 292.050 129.300 299.400 ;
        RECT 134.100 292.050 135.900 293.850 ;
        RECT 152.100 292.050 153.900 293.850 ;
        RECT 155.700 292.050 156.600 299.400 ;
        RECT 157.950 292.050 159.750 293.850 ;
        RECT 176.400 292.050 177.300 299.400 ;
        RECT 181.950 292.050 183.750 293.850 ;
        RECT 203.100 292.050 204.900 293.850 ;
        RECT 206.700 292.050 207.600 299.400 ;
        RECT 211.950 297.450 214.050 298.050 ;
        RECT 226.950 297.450 229.050 298.050 ;
        RECT 211.950 296.550 229.050 297.450 ;
        RECT 211.950 295.950 214.050 296.550 ;
        RECT 226.950 295.950 229.050 296.550 ;
        RECT 208.950 292.050 210.750 293.850 ;
        RECT 230.100 292.050 231.300 299.400 ;
        RECT 236.100 292.050 237.900 293.850 ;
        RECT 257.700 292.050 258.900 305.400 ;
        RECT 259.950 300.450 262.050 301.050 ;
        RECT 271.950 300.450 274.050 301.050 ;
        RECT 259.950 299.550 274.050 300.450 ;
        RECT 259.950 298.950 262.050 299.550 ;
        RECT 271.950 298.950 274.050 299.550 ;
        RECT 279.000 300.600 280.800 311.400 ;
        RECT 279.000 299.400 282.600 300.600 ;
        RECT 284.100 299.400 285.900 312.000 ;
        RECT 302.100 305.400 303.900 312.000 ;
        RECT 305.100 305.400 306.900 311.400 ;
        RECT 308.100 306.000 309.900 312.000 ;
        RECT 305.400 305.100 306.900 305.400 ;
        RECT 311.100 305.400 312.900 311.400 ;
        RECT 329.100 305.400 330.900 312.000 ;
        RECT 332.100 305.400 333.900 311.400 ;
        RECT 335.100 305.400 336.900 312.000 ;
        RECT 353.100 305.400 354.900 311.400 ;
        RECT 356.100 305.400 357.900 312.000 ;
        RECT 311.100 305.100 312.000 305.400 ;
        RECT 305.400 304.200 312.000 305.100 ;
        RECT 278.100 292.050 279.900 293.850 ;
        RECT 281.700 292.050 282.600 299.400 ;
        RECT 283.950 292.050 285.750 293.850 ;
        RECT 305.100 292.050 306.900 293.850 ;
        RECT 311.100 292.050 312.000 304.200 ;
        RECT 332.100 292.050 333.300 305.400 ;
        RECT 353.700 292.050 354.900 305.400 ;
        RECT 374.100 299.400 375.900 312.000 ;
        RECT 379.200 300.600 381.000 311.400 ;
        RECT 377.400 299.400 381.000 300.600 ;
        RECT 398.100 299.400 399.900 312.000 ;
        RECT 356.100 292.050 357.900 293.850 ;
        RECT 374.250 292.050 376.050 293.850 ;
        RECT 377.400 292.050 378.300 299.400 ;
        RECT 401.100 298.500 402.900 311.400 ;
        RECT 404.100 299.400 405.900 312.000 ;
        RECT 407.100 298.500 408.900 311.400 ;
        RECT 410.100 299.400 411.900 312.000 ;
        RECT 413.100 298.500 414.900 311.400 ;
        RECT 416.100 299.400 417.900 312.000 ;
        RECT 419.100 298.500 420.900 311.400 ;
        RECT 422.100 299.400 423.900 312.000 ;
        RECT 440.100 299.400 441.900 312.000 ;
        RECT 445.200 300.600 447.000 311.400 ;
        RECT 449.700 305.400 451.500 312.000 ;
        RECT 452.700 306.300 454.500 311.400 ;
        RECT 452.400 305.400 454.500 306.300 ;
        RECT 455.700 305.400 457.500 312.000 ;
        RECT 452.400 304.500 453.300 305.400 ;
        RECT 443.400 299.400 447.000 300.600 ;
        RECT 449.700 303.600 453.300 304.500 ;
        RECT 401.100 297.300 405.000 298.500 ;
        RECT 407.100 297.300 411.000 298.500 ;
        RECT 413.100 297.300 417.000 298.500 ;
        RECT 419.100 297.300 421.950 298.500 ;
        RECT 380.100 292.050 381.900 293.850 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 22.950 289.950 25.050 292.050 ;
        RECT 25.950 289.950 28.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 49.950 289.950 52.050 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 70.950 289.950 73.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 157.950 289.950 160.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 277.950 289.950 280.050 292.050 ;
        RECT 280.950 289.950 283.050 292.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 301.950 289.950 304.050 292.050 ;
        RECT 304.950 289.950 307.050 292.050 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 400.800 289.950 402.900 292.050 ;
        RECT 17.100 288.150 18.900 289.950 ;
        RECT 23.250 288.150 25.050 289.950 ;
        RECT 10.950 285.450 13.050 286.050 ;
        RECT 19.950 285.450 22.050 286.050 ;
        RECT 10.950 284.550 22.050 285.450 ;
        RECT 10.950 283.950 13.050 284.550 ;
        RECT 19.950 283.950 22.050 284.550 ;
        RECT 26.700 282.600 27.600 289.950 ;
        RECT 44.100 288.150 45.900 289.950 ;
        RECT 50.250 288.150 52.050 289.950 ;
        RECT 53.700 282.600 54.600 289.950 ;
        RECT 71.100 288.150 72.900 289.950 ;
        RECT 74.700 284.700 75.900 289.950 ;
        RECT 76.950 288.150 78.750 289.950 ;
        RECT 95.100 288.150 96.900 289.950 ;
        RECT 18.000 276.000 19.800 282.600 ;
        RECT 22.500 281.400 27.600 282.600 ;
        RECT 22.500 276.600 24.300 281.400 ;
        RECT 25.500 276.000 27.300 279.600 ;
        RECT 45.000 276.000 46.800 282.600 ;
        RECT 49.500 281.400 54.600 282.600 ;
        RECT 71.700 283.800 75.900 284.700 ;
        RECT 49.500 276.600 51.300 281.400 ;
        RECT 52.500 276.000 54.300 279.600 ;
        RECT 71.700 276.600 73.500 283.800 ;
        RECT 101.700 282.600 102.900 289.950 ;
        RECT 106.950 288.150 108.750 289.950 ;
        RECT 125.100 288.150 126.900 289.950 ;
        RECT 128.100 285.600 129.300 289.950 ;
        RECT 131.100 288.150 132.900 289.950 ;
        RECT 125.700 284.700 129.300 285.600 ;
        RECT 125.700 282.600 126.900 284.700 ;
        RECT 76.800 276.000 78.600 282.600 ;
        RECT 97.500 276.000 99.300 282.600 ;
        RECT 102.000 276.600 103.800 282.600 ;
        RECT 106.500 276.000 108.300 282.600 ;
        RECT 125.100 276.600 126.900 282.600 ;
        RECT 128.100 281.700 135.900 283.050 ;
        RECT 128.100 276.600 129.900 281.700 ;
        RECT 131.100 276.000 132.900 280.800 ;
        RECT 134.100 276.600 135.900 281.700 ;
        RECT 155.700 279.600 156.600 289.950 ;
        RECT 176.400 282.600 177.300 289.950 ;
        RECT 178.950 288.150 180.750 289.950 ;
        RECT 185.100 288.150 186.900 289.950 ;
        RECT 193.950 285.450 196.050 286.050 ;
        RECT 202.950 285.450 205.050 286.050 ;
        RECT 193.950 284.550 205.050 285.450 ;
        RECT 193.950 283.950 196.050 284.550 ;
        RECT 202.950 283.950 205.050 284.550 ;
        RECT 176.400 281.400 181.500 282.600 ;
        RECT 152.100 276.000 153.900 279.600 ;
        RECT 155.100 276.600 156.900 279.600 ;
        RECT 158.100 276.000 159.900 279.600 ;
        RECT 176.700 276.000 178.500 279.600 ;
        RECT 179.700 276.600 181.500 281.400 ;
        RECT 184.200 276.000 186.000 282.600 ;
        RECT 206.700 279.600 207.600 289.950 ;
        RECT 227.100 288.150 228.900 289.950 ;
        RECT 230.100 285.600 231.300 289.950 ;
        RECT 233.100 288.150 234.900 289.950 ;
        RECT 254.100 288.150 255.900 289.950 ;
        RECT 227.700 284.700 231.300 285.600 ;
        RECT 257.700 284.700 258.900 289.950 ;
        RECT 259.950 288.150 261.750 289.950 ;
        RECT 227.700 282.600 228.900 284.700 ;
        RECT 254.700 283.800 258.900 284.700 ;
        RECT 203.100 276.000 204.900 279.600 ;
        RECT 206.100 276.600 207.900 279.600 ;
        RECT 209.100 276.000 210.900 279.600 ;
        RECT 227.100 276.600 228.900 282.600 ;
        RECT 230.100 281.700 237.900 283.050 ;
        RECT 230.100 276.600 231.900 281.700 ;
        RECT 233.100 276.000 234.900 280.800 ;
        RECT 236.100 276.600 237.900 281.700 ;
        RECT 254.700 276.600 256.500 283.800 ;
        RECT 259.800 276.000 261.600 282.600 ;
        RECT 262.950 282.450 265.050 283.050 ;
        RECT 277.950 282.450 280.050 283.050 ;
        RECT 262.950 281.550 280.050 282.450 ;
        RECT 262.950 280.950 265.050 281.550 ;
        RECT 277.950 280.950 280.050 281.550 ;
        RECT 281.700 279.600 282.600 289.950 ;
        RECT 302.100 288.150 303.900 289.950 ;
        RECT 308.100 288.150 309.900 289.950 ;
        RECT 311.100 286.200 312.000 289.950 ;
        RECT 329.250 288.150 331.050 289.950 ;
        RECT 278.100 276.000 279.900 279.600 ;
        RECT 281.100 276.600 282.900 279.600 ;
        RECT 284.100 276.000 285.900 279.600 ;
        RECT 286.950 279.450 289.050 280.050 ;
        RECT 295.950 279.450 298.050 280.050 ;
        RECT 286.950 278.550 298.050 279.450 ;
        RECT 286.950 277.950 289.050 278.550 ;
        RECT 295.950 277.950 298.050 278.550 ;
        RECT 302.100 276.000 303.900 285.600 ;
        RECT 308.700 285.000 312.000 286.200 ;
        RECT 308.700 276.600 310.500 285.000 ;
        RECT 332.100 284.700 333.300 289.950 ;
        RECT 335.100 288.150 336.900 289.950 ;
        RECT 332.100 283.800 336.300 284.700 ;
        RECT 329.400 276.000 331.200 282.600 ;
        RECT 334.500 276.600 336.300 283.800 ;
        RECT 353.700 279.600 354.900 289.950 ;
        RECT 377.400 279.600 378.300 289.950 ;
        RECT 382.950 288.450 385.050 289.050 ;
        RECT 394.950 288.450 397.050 289.050 ;
        RECT 382.950 287.550 397.050 288.450 ;
        RECT 400.800 288.150 402.600 289.950 ;
        RECT 382.950 286.950 385.050 287.550 ;
        RECT 394.950 286.950 397.050 287.550 ;
        RECT 403.800 286.800 405.000 297.300 ;
        RECT 406.200 286.800 408.000 287.400 ;
        RECT 403.800 285.600 408.000 286.800 ;
        RECT 409.800 286.800 411.000 297.300 ;
        RECT 412.200 286.800 414.000 287.400 ;
        RECT 409.800 285.600 414.000 286.800 ;
        RECT 415.800 286.800 417.000 297.300 ;
        RECT 420.900 292.050 421.950 297.300 ;
        RECT 440.250 292.050 442.050 293.850 ;
        RECT 443.400 292.050 444.300 299.400 ;
        RECT 446.100 292.050 447.900 293.850 ;
        RECT 418.800 289.950 421.950 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 418.200 286.800 420.000 287.400 ;
        RECT 415.800 285.600 420.000 286.800 ;
        RECT 403.800 284.700 405.000 285.600 ;
        RECT 409.800 284.700 411.000 285.600 ;
        RECT 415.800 284.700 417.000 285.600 ;
        RECT 420.900 284.700 421.950 289.950 ;
        RECT 401.100 283.500 405.000 284.700 ;
        RECT 407.100 283.500 411.000 284.700 ;
        RECT 413.100 283.500 417.000 284.700 ;
        RECT 419.100 283.500 421.950 284.700 ;
        RECT 427.950 285.450 430.050 286.050 ;
        RECT 439.950 285.450 442.050 286.050 ;
        RECT 427.950 284.550 442.050 285.450 ;
        RECT 427.950 283.950 430.050 284.550 ;
        RECT 439.950 283.950 442.050 284.550 ;
        RECT 353.100 276.600 354.900 279.600 ;
        RECT 356.100 276.000 357.900 279.600 ;
        RECT 374.100 276.000 375.900 279.600 ;
        RECT 377.100 276.600 378.900 279.600 ;
        RECT 380.100 276.000 381.900 279.600 ;
        RECT 398.100 276.000 399.900 282.600 ;
        RECT 401.100 276.600 402.900 283.500 ;
        RECT 404.100 276.000 405.900 282.600 ;
        RECT 407.100 276.600 408.900 283.500 ;
        RECT 410.100 276.000 411.900 282.600 ;
        RECT 413.100 276.600 414.900 283.500 ;
        RECT 416.100 276.000 417.900 282.600 ;
        RECT 419.100 276.600 420.900 283.500 ;
        RECT 422.100 276.000 423.900 282.600 ;
        RECT 443.400 279.600 444.300 289.950 ;
        RECT 449.700 287.400 450.900 303.600 ;
        RECT 454.200 302.400 456.000 302.700 ;
        RECT 458.700 302.400 460.500 311.400 ;
        RECT 461.700 305.400 463.500 312.000 ;
        RECT 465.300 308.400 467.100 311.400 ;
        RECT 468.300 308.400 470.100 311.400 ;
        RECT 465.300 306.300 467.400 308.400 ;
        RECT 468.300 306.300 470.400 308.400 ;
        RECT 471.300 305.400 473.100 311.400 ;
        RECT 474.300 305.400 476.100 312.000 ;
        RECT 470.700 303.300 472.800 305.400 ;
        RECT 478.200 303.900 480.000 311.400 ;
        RECT 481.200 305.400 483.000 312.000 ;
        RECT 484.200 305.400 486.000 311.400 ;
        RECT 487.200 308.400 489.000 311.400 ;
        RECT 490.200 308.400 492.000 311.400 ;
        RECT 493.200 308.400 495.000 311.400 ;
        RECT 487.200 306.300 489.300 308.400 ;
        RECT 490.200 306.300 492.300 308.400 ;
        RECT 493.200 306.300 495.300 308.400 ;
        RECT 496.200 305.400 498.000 312.000 ;
        RECT 499.200 305.400 501.000 311.400 ;
        RECT 502.200 305.400 504.000 312.000 ;
        RECT 505.200 305.400 507.000 311.400 ;
        RECT 508.200 305.400 510.000 312.000 ;
        RECT 511.500 305.400 513.300 311.400 ;
        RECT 514.500 305.400 516.300 312.000 ;
        RECT 518.700 305.400 520.500 312.000 ;
        RECT 521.700 306.300 523.500 311.400 ;
        RECT 521.400 305.400 523.500 306.300 ;
        RECT 524.700 305.400 526.500 312.000 ;
        RECT 454.200 301.200 473.400 302.400 ;
        RECT 478.200 301.800 481.500 303.900 ;
        RECT 484.200 301.500 486.900 305.400 ;
        RECT 490.200 304.500 492.300 305.400 ;
        RECT 490.200 303.300 498.300 304.500 ;
        RECT 496.500 302.700 498.300 303.300 ;
        RECT 499.200 302.400 500.400 305.400 ;
        RECT 505.800 304.500 507.000 305.400 ;
        RECT 505.800 303.600 509.700 304.500 ;
        RECT 503.100 302.400 504.900 303.000 ;
        RECT 454.200 300.900 456.000 301.200 ;
        RECT 472.200 300.600 473.400 301.200 ;
        RECT 487.800 300.600 489.900 301.500 ;
        RECT 457.500 299.700 459.300 300.300 ;
        RECT 467.400 299.700 469.500 300.300 ;
        RECT 457.500 298.500 469.500 299.700 ;
        RECT 472.200 299.400 489.900 300.600 ;
        RECT 493.200 300.300 495.300 301.500 ;
        RECT 499.200 301.200 504.900 302.400 ;
        RECT 508.800 300.300 509.700 303.600 ;
        RECT 493.200 299.400 509.700 300.300 ;
        RECT 467.400 298.200 469.500 298.500 ;
        RECT 472.200 297.300 507.900 298.500 ;
        RECT 472.200 296.700 473.400 297.300 ;
        RECT 506.100 296.700 507.900 297.300 ;
        RECT 459.900 295.800 473.400 296.700 ;
        RECT 484.800 295.800 486.900 296.100 ;
        RECT 459.900 295.050 461.700 295.800 ;
        RECT 451.800 292.950 453.900 295.050 ;
        RECT 457.800 293.250 461.700 295.050 ;
        RECT 479.400 294.300 481.500 295.200 ;
        RECT 457.800 292.950 459.900 293.250 ;
        RECT 470.400 293.100 481.500 294.300 ;
        RECT 483.000 294.000 486.900 295.800 ;
        RECT 491.100 294.300 492.900 296.100 ;
        RECT 492.000 293.100 492.900 294.300 ;
        RECT 452.100 291.300 453.900 292.950 ;
        RECT 470.400 292.500 472.200 293.100 ;
        RECT 479.400 292.200 492.900 293.100 ;
        RECT 495.600 292.800 500.700 294.600 ;
        RECT 502.800 292.950 504.900 295.050 ;
        RECT 495.600 291.300 496.500 292.800 ;
        RECT 452.100 290.100 496.500 291.300 ;
        RECT 502.800 290.100 504.300 292.950 ;
        RECT 467.400 287.400 469.200 289.200 ;
        RECT 475.800 288.000 477.900 289.050 ;
        RECT 497.700 288.600 504.300 290.100 ;
        RECT 449.700 286.200 466.500 287.400 ;
        RECT 449.700 282.600 450.900 286.200 ;
        RECT 464.400 285.300 466.500 286.200 ;
        RECT 453.900 284.700 455.700 285.300 ;
        RECT 453.900 283.500 462.300 284.700 ;
        RECT 460.800 282.600 462.300 283.500 ;
        RECT 467.400 284.400 468.300 287.400 ;
        RECT 472.800 287.100 477.900 288.000 ;
        RECT 472.800 286.200 474.600 287.100 ;
        RECT 475.800 286.950 477.900 287.100 ;
        RECT 482.100 287.100 499.200 288.600 ;
        RECT 482.100 286.500 484.200 287.100 ;
        RECT 482.100 284.700 483.900 286.500 ;
        RECT 500.100 285.900 507.900 287.700 ;
        RECT 467.400 283.200 474.600 284.400 ;
        RECT 469.800 282.600 471.600 283.200 ;
        RECT 473.700 282.600 474.600 283.200 ;
        RECT 489.300 282.600 495.900 284.400 ;
        RECT 500.100 282.600 501.600 285.900 ;
        RECT 508.800 282.600 509.700 299.400 ;
        RECT 440.100 276.000 441.900 279.600 ;
        RECT 443.100 276.600 444.900 279.600 ;
        RECT 446.100 276.000 447.900 279.600 ;
        RECT 449.700 276.600 451.500 282.600 ;
        RECT 455.100 276.000 456.900 282.600 ;
        RECT 460.500 276.600 462.300 282.600 ;
        RECT 464.700 279.600 466.800 281.700 ;
        RECT 467.700 279.600 469.800 281.700 ;
        RECT 470.700 279.600 472.800 281.700 ;
        RECT 473.700 281.400 476.400 282.600 ;
        RECT 474.600 280.500 476.400 281.400 ;
        RECT 478.200 280.500 480.900 282.600 ;
        RECT 464.700 276.600 466.500 279.600 ;
        RECT 467.700 276.600 469.500 279.600 ;
        RECT 470.700 276.600 472.500 279.600 ;
        RECT 473.700 276.000 475.500 279.600 ;
        RECT 478.200 276.600 480.000 280.500 ;
        RECT 484.200 279.600 486.300 281.700 ;
        RECT 487.200 279.600 489.300 281.700 ;
        RECT 490.200 279.600 492.300 281.700 ;
        RECT 493.200 279.600 495.300 281.700 ;
        RECT 497.400 281.400 501.600 282.600 ;
        RECT 481.200 276.000 483.000 279.600 ;
        RECT 484.200 276.600 486.000 279.600 ;
        RECT 487.200 276.600 489.000 279.600 ;
        RECT 490.200 276.600 492.000 279.600 ;
        RECT 493.200 276.600 495.000 279.600 ;
        RECT 497.400 276.600 499.200 281.400 ;
        RECT 502.500 276.000 504.300 282.600 ;
        RECT 507.900 276.600 509.700 282.600 ;
        RECT 511.500 295.050 513.000 305.400 ;
        RECT 521.400 304.500 522.300 305.400 ;
        RECT 518.700 303.600 522.300 304.500 ;
        RECT 511.500 292.950 513.900 295.050 ;
        RECT 511.500 279.600 513.000 292.950 ;
        RECT 518.700 287.400 519.900 303.600 ;
        RECT 523.200 302.400 525.000 302.700 ;
        RECT 527.700 302.400 529.500 311.400 ;
        RECT 530.700 305.400 532.500 312.000 ;
        RECT 534.300 308.400 536.100 311.400 ;
        RECT 537.300 308.400 539.100 311.400 ;
        RECT 534.300 306.300 536.400 308.400 ;
        RECT 537.300 306.300 539.400 308.400 ;
        RECT 540.300 305.400 542.100 311.400 ;
        RECT 543.300 305.400 545.100 312.000 ;
        RECT 539.700 303.300 541.800 305.400 ;
        RECT 547.200 303.900 549.000 311.400 ;
        RECT 550.200 305.400 552.000 312.000 ;
        RECT 553.200 305.400 555.000 311.400 ;
        RECT 556.200 308.400 558.000 311.400 ;
        RECT 559.200 308.400 561.000 311.400 ;
        RECT 562.200 308.400 564.000 311.400 ;
        RECT 556.200 306.300 558.300 308.400 ;
        RECT 559.200 306.300 561.300 308.400 ;
        RECT 562.200 306.300 564.300 308.400 ;
        RECT 565.200 305.400 567.000 312.000 ;
        RECT 568.200 305.400 570.000 311.400 ;
        RECT 571.200 305.400 573.000 312.000 ;
        RECT 574.200 305.400 576.000 311.400 ;
        RECT 577.200 305.400 579.000 312.000 ;
        RECT 580.500 305.400 582.300 311.400 ;
        RECT 583.500 305.400 585.300 312.000 ;
        RECT 523.200 301.200 542.400 302.400 ;
        RECT 547.200 301.800 550.500 303.900 ;
        RECT 553.200 301.500 555.900 305.400 ;
        RECT 559.200 304.500 561.300 305.400 ;
        RECT 559.200 303.300 567.300 304.500 ;
        RECT 565.500 302.700 567.300 303.300 ;
        RECT 568.200 302.400 569.400 305.400 ;
        RECT 574.800 304.500 576.000 305.400 ;
        RECT 574.800 303.600 578.700 304.500 ;
        RECT 572.100 302.400 573.900 303.000 ;
        RECT 523.200 300.900 525.000 301.200 ;
        RECT 541.200 300.600 542.400 301.200 ;
        RECT 556.800 300.600 558.900 301.500 ;
        RECT 526.500 299.700 528.300 300.300 ;
        RECT 536.400 299.700 538.500 300.300 ;
        RECT 526.500 298.500 538.500 299.700 ;
        RECT 541.200 299.400 558.900 300.600 ;
        RECT 562.200 300.300 564.300 301.500 ;
        RECT 568.200 301.200 573.900 302.400 ;
        RECT 577.800 300.300 578.700 303.600 ;
        RECT 562.200 299.400 578.700 300.300 ;
        RECT 536.400 298.200 538.500 298.500 ;
        RECT 541.200 297.300 576.900 298.500 ;
        RECT 541.200 296.700 542.400 297.300 ;
        RECT 575.100 296.700 576.900 297.300 ;
        RECT 528.900 295.800 542.400 296.700 ;
        RECT 553.800 295.800 555.900 296.100 ;
        RECT 528.900 295.050 530.700 295.800 ;
        RECT 520.800 292.950 522.900 295.050 ;
        RECT 526.800 293.250 530.700 295.050 ;
        RECT 548.400 294.300 550.500 295.200 ;
        RECT 526.800 292.950 528.900 293.250 ;
        RECT 539.400 293.100 550.500 294.300 ;
        RECT 552.000 294.000 555.900 295.800 ;
        RECT 560.100 294.300 561.900 296.100 ;
        RECT 561.000 293.100 561.900 294.300 ;
        RECT 521.100 291.300 522.900 292.950 ;
        RECT 539.400 292.500 541.200 293.100 ;
        RECT 548.400 292.200 561.900 293.100 ;
        RECT 564.600 292.800 569.700 294.600 ;
        RECT 571.800 292.950 573.900 295.050 ;
        RECT 564.600 291.300 565.500 292.800 ;
        RECT 521.100 290.100 565.500 291.300 ;
        RECT 571.800 290.100 573.300 292.950 ;
        RECT 536.400 287.400 538.200 289.200 ;
        RECT 544.800 288.000 546.900 289.050 ;
        RECT 566.700 288.600 573.300 290.100 ;
        RECT 518.700 286.200 535.500 287.400 ;
        RECT 518.700 282.600 519.900 286.200 ;
        RECT 533.400 285.300 535.500 286.200 ;
        RECT 522.900 284.700 524.700 285.300 ;
        RECT 522.900 283.500 531.300 284.700 ;
        RECT 529.800 282.600 531.300 283.500 ;
        RECT 536.400 284.400 537.300 287.400 ;
        RECT 541.800 287.100 546.900 288.000 ;
        RECT 541.800 286.200 543.600 287.100 ;
        RECT 544.800 286.950 546.900 287.100 ;
        RECT 551.100 287.100 568.200 288.600 ;
        RECT 551.100 286.500 553.200 287.100 ;
        RECT 551.100 284.700 552.900 286.500 ;
        RECT 569.100 285.900 576.900 287.700 ;
        RECT 536.400 283.200 543.600 284.400 ;
        RECT 538.800 282.600 540.600 283.200 ;
        RECT 542.700 282.600 543.600 283.200 ;
        RECT 558.300 282.600 564.900 284.400 ;
        RECT 569.100 282.600 570.600 285.900 ;
        RECT 577.800 282.600 578.700 299.400 ;
        RECT 511.500 276.600 513.300 279.600 ;
        RECT 514.500 276.000 516.300 279.600 ;
        RECT 518.700 276.600 520.500 282.600 ;
        RECT 524.100 276.000 525.900 282.600 ;
        RECT 529.500 276.600 531.300 282.600 ;
        RECT 533.700 279.600 535.800 281.700 ;
        RECT 536.700 279.600 538.800 281.700 ;
        RECT 539.700 279.600 541.800 281.700 ;
        RECT 542.700 281.400 545.400 282.600 ;
        RECT 543.600 280.500 545.400 281.400 ;
        RECT 547.200 280.500 549.900 282.600 ;
        RECT 533.700 276.600 535.500 279.600 ;
        RECT 536.700 276.600 538.500 279.600 ;
        RECT 539.700 276.600 541.500 279.600 ;
        RECT 542.700 276.000 544.500 279.600 ;
        RECT 547.200 276.600 549.000 280.500 ;
        RECT 553.200 279.600 555.300 281.700 ;
        RECT 556.200 279.600 558.300 281.700 ;
        RECT 559.200 279.600 561.300 281.700 ;
        RECT 562.200 279.600 564.300 281.700 ;
        RECT 566.400 281.400 570.600 282.600 ;
        RECT 550.200 276.000 552.000 279.600 ;
        RECT 553.200 276.600 555.000 279.600 ;
        RECT 556.200 276.600 558.000 279.600 ;
        RECT 559.200 276.600 561.000 279.600 ;
        RECT 562.200 276.600 564.000 279.600 ;
        RECT 566.400 276.600 568.200 281.400 ;
        RECT 571.500 276.000 573.300 282.600 ;
        RECT 576.900 276.600 578.700 282.600 ;
        RECT 580.500 295.050 582.000 305.400 ;
        RECT 602.400 299.400 604.200 312.000 ;
        RECT 607.500 300.900 609.300 311.400 ;
        RECT 610.500 305.400 612.300 312.000 ;
        RECT 629.700 305.400 631.500 312.000 ;
        RECT 610.200 302.100 612.000 303.900 ;
        RECT 630.000 302.100 631.800 303.900 ;
        RECT 632.700 300.900 634.500 311.400 ;
        RECT 607.500 299.400 609.900 300.900 ;
        RECT 580.500 292.950 582.900 295.050 ;
        RECT 580.500 279.600 582.000 292.950 ;
        RECT 602.100 292.050 603.900 293.850 ;
        RECT 608.700 292.050 609.900 299.400 ;
        RECT 632.100 299.400 634.500 300.900 ;
        RECT 637.800 299.400 639.600 312.000 ;
        RECT 656.400 299.400 658.200 312.000 ;
        RECT 661.500 300.900 663.300 311.400 ;
        RECT 664.500 305.400 666.300 312.000 ;
        RECT 683.700 305.400 685.500 312.000 ;
        RECT 664.200 302.100 666.000 303.900 ;
        RECT 684.000 302.100 685.800 303.900 ;
        RECT 686.700 300.900 688.500 311.400 ;
        RECT 661.500 299.400 663.900 300.900 ;
        RECT 632.100 292.050 633.300 299.400 ;
        RECT 638.100 292.050 639.900 293.850 ;
        RECT 656.100 292.050 657.900 293.850 ;
        RECT 662.700 292.050 663.900 299.400 ;
        RECT 686.100 299.400 688.500 300.900 ;
        RECT 691.800 299.400 693.600 312.000 ;
        RECT 710.700 305.400 712.500 312.000 ;
        RECT 711.000 302.100 712.800 303.900 ;
        RECT 713.700 300.900 715.500 311.400 ;
        RECT 713.100 299.400 715.500 300.900 ;
        RECT 718.800 299.400 720.600 312.000 ;
        RECT 738.000 300.600 739.800 311.400 ;
        RECT 738.000 299.400 741.600 300.600 ;
        RECT 743.100 299.400 744.900 312.000 ;
        RECT 761.100 305.400 762.900 312.000 ;
        RECT 764.100 305.400 765.900 311.400 ;
        RECT 767.100 305.400 768.900 312.000 ;
        RECT 686.100 292.050 687.300 299.400 ;
        RECT 688.950 297.450 691.050 298.200 ;
        RECT 697.950 297.450 700.050 298.050 ;
        RECT 688.950 296.550 700.050 297.450 ;
        RECT 688.950 296.100 691.050 296.550 ;
        RECT 697.950 295.950 700.050 296.550 ;
        RECT 700.950 294.450 703.050 295.050 ;
        RECT 706.950 294.450 709.050 295.050 ;
        RECT 692.100 292.050 693.900 293.850 ;
        RECT 700.950 293.550 709.050 294.450 ;
        RECT 700.950 292.950 703.050 293.550 ;
        RECT 706.950 292.950 709.050 293.550 ;
        RECT 713.100 292.050 714.300 299.400 ;
        RECT 719.100 292.050 720.900 293.850 ;
        RECT 737.100 292.050 738.900 293.850 ;
        RECT 740.700 292.050 741.600 299.400 ;
        RECT 742.950 297.450 745.050 298.050 ;
        RECT 760.950 297.450 763.050 298.050 ;
        RECT 742.950 296.550 763.050 297.450 ;
        RECT 742.950 295.950 745.050 296.550 ;
        RECT 760.950 295.950 763.050 296.550 ;
        RECT 745.950 294.450 748.050 295.050 ;
        RECT 742.950 292.050 744.750 293.850 ;
        RECT 745.950 293.550 756.450 294.450 ;
        RECT 745.950 292.950 748.050 293.550 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 610.950 289.950 613.050 292.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 605.100 288.150 606.900 289.950 ;
        RECT 608.700 285.600 609.900 289.950 ;
        RECT 611.100 288.150 612.900 289.950 ;
        RECT 629.100 288.150 630.900 289.950 ;
        RECT 632.100 285.600 633.300 289.950 ;
        RECT 635.100 288.150 636.900 289.950 ;
        RECT 659.100 288.150 660.900 289.950 ;
        RECT 608.700 284.700 612.300 285.600 ;
        RECT 602.100 281.700 609.900 283.050 ;
        RECT 580.500 276.600 582.300 279.600 ;
        RECT 583.500 276.000 585.300 279.600 ;
        RECT 602.100 276.600 603.900 281.700 ;
        RECT 605.100 276.000 606.900 280.800 ;
        RECT 608.100 276.600 609.900 281.700 ;
        RECT 611.100 282.600 612.300 284.700 ;
        RECT 629.700 284.700 633.300 285.600 ;
        RECT 662.700 285.600 663.900 289.950 ;
        RECT 665.100 288.150 666.900 289.950 ;
        RECT 683.100 288.150 684.900 289.950 ;
        RECT 686.100 285.600 687.300 289.950 ;
        RECT 689.100 288.150 690.900 289.950 ;
        RECT 710.100 288.150 711.900 289.950 ;
        RECT 713.100 285.600 714.300 289.950 ;
        RECT 716.100 288.150 717.900 289.950 ;
        RECT 662.700 284.700 666.300 285.600 ;
        RECT 629.700 282.600 630.900 284.700 ;
        RECT 611.100 276.600 612.900 282.600 ;
        RECT 629.100 276.600 630.900 282.600 ;
        RECT 632.100 281.700 639.900 283.050 ;
        RECT 632.100 276.600 633.900 281.700 ;
        RECT 635.100 276.000 636.900 280.800 ;
        RECT 638.100 276.600 639.900 281.700 ;
        RECT 656.100 281.700 663.900 283.050 ;
        RECT 656.100 276.600 657.900 281.700 ;
        RECT 659.100 276.000 660.900 280.800 ;
        RECT 662.100 276.600 663.900 281.700 ;
        RECT 665.100 282.600 666.300 284.700 ;
        RECT 683.700 284.700 687.300 285.600 ;
        RECT 710.700 284.700 714.300 285.600 ;
        RECT 683.700 282.600 684.900 284.700 ;
        RECT 665.100 276.600 666.900 282.600 ;
        RECT 683.100 276.600 684.900 282.600 ;
        RECT 686.100 281.700 693.900 283.050 ;
        RECT 710.700 282.600 711.900 284.700 ;
        RECT 686.100 276.600 687.900 281.700 ;
        RECT 689.100 276.000 690.900 280.800 ;
        RECT 692.100 276.600 693.900 281.700 ;
        RECT 710.100 276.600 711.900 282.600 ;
        RECT 713.100 281.700 720.900 283.050 ;
        RECT 713.100 276.600 714.900 281.700 ;
        RECT 716.100 276.000 717.900 280.800 ;
        RECT 719.100 276.600 720.900 281.700 ;
        RECT 740.700 279.600 741.600 289.950 ;
        RECT 755.550 289.050 756.450 293.550 ;
        RECT 764.100 292.050 765.300 305.400 ;
        RECT 766.950 303.450 769.050 304.050 ;
        RECT 778.950 303.450 781.050 304.050 ;
        RECT 766.950 302.550 781.050 303.450 ;
        RECT 766.950 301.950 769.050 302.550 ;
        RECT 778.950 301.950 781.050 302.550 ;
        RECT 785.100 300.600 786.900 311.400 ;
        RECT 788.100 301.500 790.200 312.000 ;
        RECT 785.100 299.400 790.200 300.600 ;
        RECT 792.600 300.300 794.400 311.400 ;
        RECT 797.100 301.500 798.900 312.000 ;
        RECT 800.100 300.300 801.900 311.400 ;
        RECT 803.700 305.400 805.500 312.000 ;
        RECT 806.700 305.400 808.500 311.400 ;
        RECT 810.000 305.400 811.800 312.000 ;
        RECT 813.000 305.400 814.800 311.400 ;
        RECT 816.000 305.400 817.800 312.000 ;
        RECT 819.000 305.400 820.800 311.400 ;
        RECT 822.000 305.400 823.800 312.000 ;
        RECT 825.000 308.400 826.800 311.400 ;
        RECT 828.000 308.400 829.800 311.400 ;
        RECT 831.000 308.400 832.800 311.400 ;
        RECT 824.700 306.300 826.800 308.400 ;
        RECT 827.700 306.300 829.800 308.400 ;
        RECT 830.700 306.300 832.800 308.400 ;
        RECT 834.000 305.400 835.800 311.400 ;
        RECT 837.000 305.400 838.800 312.000 ;
        RECT 788.100 298.500 790.200 299.400 ;
        RECT 791.100 299.400 794.400 300.300 ;
        RECT 791.100 295.050 792.300 299.400 ;
        RECT 797.100 299.100 801.900 300.300 ;
        RECT 797.100 298.200 799.200 299.100 ;
        RECT 793.800 297.300 799.200 298.200 ;
        RECT 793.800 295.500 795.600 297.300 ;
        RECT 807.000 295.050 808.500 305.400 ;
        RECT 813.000 304.500 814.200 305.400 ;
        RECT 790.800 294.300 792.900 295.050 ;
        RECT 785.400 292.050 787.200 293.850 ;
        RECT 790.800 292.950 793.800 294.300 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 785.100 289.950 787.200 292.050 ;
        RECT 790.200 290.100 792.000 291.900 ;
        RECT 755.550 287.550 760.050 289.050 ;
        RECT 761.250 288.150 763.050 289.950 ;
        RECT 756.000 286.950 760.050 287.550 ;
        RECT 764.100 284.700 765.300 289.950 ;
        RECT 767.100 288.150 768.900 289.950 ;
        RECT 789.900 288.000 792.000 290.100 ;
        RECT 792.900 286.200 793.800 292.950 ;
        RECT 795.300 292.200 797.100 294.000 ;
        RECT 806.100 292.950 808.500 295.050 ;
        RECT 795.000 290.100 797.100 292.200 ;
        RECT 799.800 289.800 801.900 292.050 ;
        RECT 799.800 289.200 801.600 289.800 ;
        RECT 795.000 288.000 801.600 289.200 ;
        RECT 795.000 287.100 797.100 288.000 ;
        RECT 764.100 283.800 768.300 284.700 ;
        RECT 737.100 276.000 738.900 279.600 ;
        RECT 740.100 276.600 741.900 279.600 ;
        RECT 743.100 276.000 744.900 279.600 ;
        RECT 761.400 276.000 763.200 282.600 ;
        RECT 766.500 276.600 768.300 283.800 ;
        RECT 787.500 283.500 789.600 285.900 ;
        RECT 790.800 284.100 793.800 286.200 ;
        RECT 794.700 285.300 796.500 287.100 ;
        RECT 785.100 282.600 789.600 283.500 ;
        RECT 785.100 276.600 786.900 282.600 ;
        RECT 792.900 282.000 793.800 284.100 ;
        RECT 797.400 285.000 799.500 285.600 ;
        RECT 797.400 283.500 801.900 285.000 ;
        RECT 800.400 282.600 801.900 283.500 ;
        RECT 788.400 276.000 790.200 281.700 ;
        RECT 792.900 276.600 794.700 282.000 ;
        RECT 797.100 276.000 798.900 281.700 ;
        RECT 800.100 276.600 801.900 282.600 ;
        RECT 807.000 279.600 808.500 292.950 ;
        RECT 803.700 276.000 805.500 279.600 ;
        RECT 806.700 276.600 808.500 279.600 ;
        RECT 810.300 303.600 814.200 304.500 ;
        RECT 810.300 300.300 811.200 303.600 ;
        RECT 815.100 302.400 816.900 303.000 ;
        RECT 819.600 302.400 820.800 305.400 ;
        RECT 827.700 304.500 829.800 305.400 ;
        RECT 821.700 303.300 829.800 304.500 ;
        RECT 821.700 302.700 823.500 303.300 ;
        RECT 815.100 301.200 820.800 302.400 ;
        RECT 833.100 301.500 835.800 305.400 ;
        RECT 840.000 303.900 841.800 311.400 ;
        RECT 843.900 305.400 845.700 312.000 ;
        RECT 846.900 305.400 848.700 311.400 ;
        RECT 849.900 308.400 851.700 311.400 ;
        RECT 852.900 308.400 854.700 311.400 ;
        RECT 849.600 306.300 851.700 308.400 ;
        RECT 852.600 306.300 854.700 308.400 ;
        RECT 856.500 305.400 858.300 312.000 ;
        RECT 838.500 301.800 841.800 303.900 ;
        RECT 847.200 303.300 849.300 305.400 ;
        RECT 859.500 302.400 861.300 311.400 ;
        RECT 862.500 305.400 864.300 312.000 ;
        RECT 865.500 306.300 867.300 311.400 ;
        RECT 865.500 305.400 867.600 306.300 ;
        RECT 868.500 305.400 870.300 312.000 ;
        RECT 874.950 309.450 877.050 310.050 ;
        RECT 883.950 309.450 886.050 310.050 ;
        RECT 874.950 308.550 886.050 309.450 ;
        RECT 874.950 307.950 877.050 308.550 ;
        RECT 883.950 307.950 886.050 308.550 ;
        RECT 866.700 304.500 867.600 305.400 ;
        RECT 866.700 303.600 870.300 304.500 ;
        RECT 864.000 302.400 865.800 302.700 ;
        RECT 824.700 300.300 826.800 301.500 ;
        RECT 810.300 299.400 826.800 300.300 ;
        RECT 830.100 300.600 832.200 301.500 ;
        RECT 846.600 301.200 865.800 302.400 ;
        RECT 846.600 300.600 847.800 301.200 ;
        RECT 864.000 300.900 865.800 301.200 ;
        RECT 830.100 299.400 847.800 300.600 ;
        RECT 850.500 299.700 852.600 300.300 ;
        RECT 860.700 299.700 862.500 300.300 ;
        RECT 810.300 282.600 811.200 299.400 ;
        RECT 850.500 298.500 862.500 299.700 ;
        RECT 812.100 297.300 847.800 298.500 ;
        RECT 850.500 298.200 852.600 298.500 ;
        RECT 812.100 296.700 813.900 297.300 ;
        RECT 846.600 296.700 847.800 297.300 ;
        RECT 815.100 292.950 817.200 295.050 ;
        RECT 815.700 290.100 817.200 292.950 ;
        RECT 819.300 292.800 824.400 294.600 ;
        RECT 823.500 291.300 824.400 292.800 ;
        RECT 827.100 294.300 828.900 296.100 ;
        RECT 833.100 295.800 835.200 296.100 ;
        RECT 846.600 295.800 860.100 296.700 ;
        RECT 827.100 293.100 828.000 294.300 ;
        RECT 833.100 294.000 837.000 295.800 ;
        RECT 838.500 294.300 840.600 295.200 ;
        RECT 858.300 295.050 860.100 295.800 ;
        RECT 838.500 293.100 849.600 294.300 ;
        RECT 858.300 293.250 862.200 295.050 ;
        RECT 827.100 292.200 840.600 293.100 ;
        RECT 847.800 292.500 849.600 293.100 ;
        RECT 860.100 292.950 862.200 293.250 ;
        RECT 866.100 292.950 868.200 295.050 ;
        RECT 866.100 291.300 867.900 292.950 ;
        RECT 823.500 290.100 867.900 291.300 ;
        RECT 815.700 288.600 822.300 290.100 ;
        RECT 812.100 285.900 819.900 287.700 ;
        RECT 820.800 287.100 837.900 288.600 ;
        RECT 835.800 286.500 837.900 287.100 ;
        RECT 842.100 288.000 844.200 289.050 ;
        RECT 842.100 287.100 847.200 288.000 ;
        RECT 850.800 287.400 852.600 289.200 ;
        RECT 869.100 287.400 870.300 303.600 ;
        RECT 887.400 299.400 889.200 312.000 ;
        RECT 892.500 300.900 894.300 311.400 ;
        RECT 895.500 305.400 897.300 312.000 ;
        RECT 895.200 302.100 897.000 303.900 ;
        RECT 892.500 299.400 894.900 300.900 ;
        RECT 880.950 297.450 883.050 298.050 ;
        RECT 889.950 297.450 892.050 298.050 ;
        RECT 880.950 296.550 892.050 297.450 ;
        RECT 880.950 295.950 883.050 296.550 ;
        RECT 889.950 295.950 892.050 296.550 ;
        RECT 887.100 292.050 888.900 293.850 ;
        RECT 893.700 292.050 894.900 299.400 ;
        RECT 901.950 300.450 904.050 301.050 ;
        RECT 907.950 300.450 910.050 301.050 ;
        RECT 901.950 299.550 910.050 300.450 ;
        RECT 901.950 298.950 904.050 299.550 ;
        RECT 907.950 298.950 910.050 299.550 ;
        RECT 914.400 299.400 916.200 312.000 ;
        RECT 919.500 300.900 921.300 311.400 ;
        RECT 922.500 305.400 924.300 312.000 ;
        RECT 922.200 302.100 924.000 303.900 ;
        RECT 919.500 299.400 921.900 300.900 ;
        RECT 941.100 300.300 942.900 311.400 ;
        RECT 944.100 301.500 945.900 312.000 ;
        RECT 941.100 299.400 945.600 300.300 ;
        RECT 948.600 299.400 950.400 311.400 ;
        RECT 953.100 301.500 954.900 312.000 ;
        RECT 956.100 300.600 957.900 311.400 ;
        RECT 974.100 305.400 975.900 311.400 ;
        RECT 977.100 306.000 978.900 312.000 ;
        RECT 975.000 305.100 975.900 305.400 ;
        RECT 980.100 305.400 981.900 311.400 ;
        RECT 983.100 305.400 984.900 312.000 ;
        RECT 980.100 305.100 981.600 305.400 ;
        RECT 975.000 304.200 981.600 305.100 ;
        RECT 958.950 303.450 961.050 304.050 ;
        RECT 967.950 303.450 970.050 304.050 ;
        RECT 958.950 302.550 970.050 303.450 ;
        RECT 958.950 301.950 961.050 302.550 ;
        RECT 967.950 301.950 970.050 302.550 ;
        RECT 895.950 297.450 898.050 298.050 ;
        RECT 904.950 297.450 907.050 298.050 ;
        RECT 895.950 296.550 907.050 297.450 ;
        RECT 895.950 295.950 898.050 296.550 ;
        RECT 904.950 295.950 907.050 296.550 ;
        RECT 914.100 292.050 915.900 293.850 ;
        RECT 920.700 292.050 921.900 299.400 ;
        RECT 943.500 297.300 945.600 299.400 ;
        RECT 949.200 298.050 950.400 299.400 ;
        RECT 953.100 299.400 957.900 300.600 ;
        RECT 953.100 298.500 955.200 299.400 ;
        RECT 949.200 297.000 950.700 298.050 ;
        RECT 946.800 295.500 948.900 295.800 ;
        RECT 945.000 293.700 948.900 295.500 ;
        RECT 949.800 295.050 950.700 297.000 ;
        RECT 949.800 292.950 951.900 295.050 ;
        RECT 949.800 292.800 951.300 292.950 ;
        RECT 946.200 292.050 948.000 292.500 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 892.950 289.950 895.050 292.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 913.950 289.950 916.050 292.050 ;
        RECT 916.950 289.950 919.050 292.050 ;
        RECT 919.950 289.950 922.050 292.050 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 941.100 290.700 948.000 292.050 ;
        RECT 948.900 291.900 951.300 292.800 ;
        RECT 955.800 292.050 957.600 293.850 ;
        RECT 975.000 292.050 975.900 304.200 ;
        RECT 985.950 303.450 988.050 304.050 ;
        RECT 991.950 303.450 994.050 303.900 ;
        RECT 985.950 302.550 994.050 303.450 ;
        RECT 985.950 301.950 988.050 302.550 ;
        RECT 991.950 301.800 994.050 302.550 ;
        RECT 1002.600 300.900 1004.400 311.400 ;
        RECT 1002.000 299.400 1004.400 300.900 ;
        RECT 1005.600 299.400 1007.400 312.000 ;
        RECT 1010.100 299.400 1011.900 311.400 ;
        RECT 1028.100 305.400 1029.900 312.000 ;
        RECT 1031.100 305.400 1032.900 311.400 ;
        RECT 1034.100 305.400 1035.900 312.000 ;
        RECT 985.950 294.450 988.050 295.050 ;
        RECT 997.950 294.450 1000.050 295.050 ;
        RECT 980.100 292.050 981.900 293.850 ;
        RECT 985.950 293.550 1000.050 294.450 ;
        RECT 985.950 292.950 988.050 293.550 ;
        RECT 997.950 292.950 1000.050 293.550 ;
        RECT 1002.000 292.050 1003.200 299.400 ;
        RECT 1010.700 297.900 1011.900 299.400 ;
        RECT 1004.100 296.700 1011.900 297.900 ;
        RECT 1004.100 296.100 1005.900 296.700 ;
        RECT 941.100 289.950 943.200 290.700 ;
        RECT 890.100 288.150 891.900 289.950 ;
        RECT 842.100 286.950 844.200 287.100 ;
        RECT 818.400 282.600 819.900 285.900 ;
        RECT 836.100 284.700 837.900 286.500 ;
        RECT 845.400 286.200 847.200 287.100 ;
        RECT 851.700 284.400 852.600 287.400 ;
        RECT 853.500 286.200 870.300 287.400 ;
        RECT 853.500 285.300 855.600 286.200 ;
        RECT 864.300 284.700 866.100 285.300 ;
        RECT 824.100 282.600 830.700 284.400 ;
        RECT 845.400 283.200 852.600 284.400 ;
        RECT 857.700 283.500 866.100 284.700 ;
        RECT 845.400 282.600 846.300 283.200 ;
        RECT 848.400 282.600 850.200 283.200 ;
        RECT 857.700 282.600 859.200 283.500 ;
        RECT 869.100 282.600 870.300 286.200 ;
        RECT 893.700 285.600 894.900 289.950 ;
        RECT 896.100 288.150 897.900 289.950 ;
        RECT 917.100 288.150 918.900 289.950 ;
        RECT 920.700 285.600 921.900 289.950 ;
        RECT 923.100 288.150 924.900 289.950 ;
        RECT 941.400 288.150 943.200 289.950 ;
        RECT 946.200 287.400 948.000 289.200 ;
        RECT 893.700 284.700 897.300 285.600 ;
        RECT 920.700 284.700 924.300 285.600 ;
        RECT 945.900 285.300 948.000 287.400 ;
        RECT 810.300 276.600 812.100 282.600 ;
        RECT 815.700 276.000 817.500 282.600 ;
        RECT 818.400 281.400 822.600 282.600 ;
        RECT 820.800 276.600 822.600 281.400 ;
        RECT 824.700 279.600 826.800 281.700 ;
        RECT 827.700 279.600 829.800 281.700 ;
        RECT 830.700 279.600 832.800 281.700 ;
        RECT 833.700 279.600 835.800 281.700 ;
        RECT 839.100 280.500 841.800 282.600 ;
        RECT 843.600 281.400 846.300 282.600 ;
        RECT 843.600 280.500 845.400 281.400 ;
        RECT 825.000 276.600 826.800 279.600 ;
        RECT 828.000 276.600 829.800 279.600 ;
        RECT 831.000 276.600 832.800 279.600 ;
        RECT 834.000 276.600 835.800 279.600 ;
        RECT 837.000 276.000 838.800 279.600 ;
        RECT 840.000 276.600 841.800 280.500 ;
        RECT 847.200 279.600 849.300 281.700 ;
        RECT 850.200 279.600 852.300 281.700 ;
        RECT 853.200 279.600 855.300 281.700 ;
        RECT 844.500 276.000 846.300 279.600 ;
        RECT 847.500 276.600 849.300 279.600 ;
        RECT 850.500 276.600 852.300 279.600 ;
        RECT 853.500 276.600 855.300 279.600 ;
        RECT 857.700 276.600 859.500 282.600 ;
        RECT 863.100 276.000 864.900 282.600 ;
        RECT 868.500 276.600 870.300 282.600 ;
        RECT 887.100 281.700 894.900 283.050 ;
        RECT 887.100 276.600 888.900 281.700 ;
        RECT 890.100 276.000 891.900 280.800 ;
        RECT 893.100 276.600 894.900 281.700 ;
        RECT 896.100 282.600 897.300 284.700 ;
        RECT 896.100 276.600 897.900 282.600 ;
        RECT 914.100 281.700 921.900 283.050 ;
        RECT 914.100 276.600 915.900 281.700 ;
        RECT 917.100 276.000 918.900 280.800 ;
        RECT 920.100 276.600 921.900 281.700 ;
        RECT 923.100 282.600 924.300 284.700 ;
        RECT 941.700 284.400 948.000 285.300 ;
        RECT 948.900 286.200 950.100 291.900 ;
        RECT 951.300 289.200 953.100 291.000 ;
        RECT 955.800 289.950 957.900 292.050 ;
        RECT 973.950 289.950 976.050 292.050 ;
        RECT 976.950 289.950 979.050 292.050 ;
        RECT 979.950 289.950 982.050 292.050 ;
        RECT 982.950 289.950 985.050 292.050 ;
        RECT 1001.100 289.950 1003.200 292.050 ;
        RECT 951.000 287.100 953.100 289.200 ;
        RECT 975.000 286.200 975.900 289.950 ;
        RECT 977.100 288.150 978.900 289.950 ;
        RECT 983.100 288.150 984.900 289.950 ;
        RECT 941.700 282.600 942.900 284.400 ;
        RECT 948.900 284.100 951.900 286.200 ;
        RECT 975.000 285.000 978.300 286.200 ;
        RECT 948.900 282.600 950.100 284.100 ;
        RECT 953.100 283.500 955.200 284.700 ;
        RECT 953.100 282.600 957.900 283.500 ;
        RECT 923.100 276.600 924.900 282.600 ;
        RECT 941.100 276.600 942.900 282.600 ;
        RECT 944.100 276.000 945.900 281.700 ;
        RECT 948.600 276.600 950.400 282.600 ;
        RECT 953.100 276.000 954.900 281.700 ;
        RECT 956.100 276.600 957.900 282.600 ;
        RECT 961.950 282.450 964.050 283.050 ;
        RECT 970.950 282.450 973.050 283.050 ;
        RECT 961.950 281.550 973.050 282.450 ;
        RECT 961.950 280.950 964.050 281.550 ;
        RECT 970.950 280.950 973.050 281.550 ;
        RECT 976.500 276.600 978.300 285.000 ;
        RECT 983.100 276.000 984.900 285.600 ;
        RECT 1001.100 282.600 1002.000 289.950 ;
        RECT 1004.400 285.600 1005.300 296.100 ;
        RECT 1006.200 292.050 1008.000 293.850 ;
        RECT 1031.700 292.050 1032.900 305.400 ;
        RECT 1006.500 289.950 1008.600 292.050 ;
        RECT 1009.800 289.950 1011.900 292.050 ;
        RECT 1027.950 289.950 1030.050 292.050 ;
        RECT 1030.950 289.950 1033.050 292.050 ;
        RECT 1033.950 289.950 1036.050 292.050 ;
        RECT 1009.800 288.150 1011.600 289.950 ;
        RECT 1028.100 288.150 1029.900 289.950 ;
        RECT 1003.200 284.700 1005.300 285.600 ;
        RECT 1031.700 284.700 1032.900 289.950 ;
        RECT 1033.950 288.150 1035.750 289.950 ;
        RECT 1003.200 283.800 1008.600 284.700 ;
        RECT 1001.100 276.600 1002.900 282.600 ;
        RECT 1004.100 276.000 1005.900 282.000 ;
        RECT 1007.700 279.600 1008.600 283.800 ;
        RECT 1028.700 283.800 1032.900 284.700 ;
        RECT 1007.100 276.600 1008.900 279.600 ;
        RECT 1010.100 276.600 1011.900 279.600 ;
        RECT 1028.700 276.600 1030.500 283.800 ;
        RECT 1010.700 276.000 1011.900 276.600 ;
        RECT 1033.800 276.000 1035.600 282.600 ;
        RECT 17.100 266.400 18.900 272.400 ;
        RECT 20.100 267.300 21.900 273.000 ;
        RECT 24.600 266.400 26.400 272.400 ;
        RECT 29.100 267.300 30.900 273.000 ;
        RECT 32.100 266.400 33.900 272.400 ;
        RECT 50.100 269.400 51.900 272.400 ;
        RECT 53.100 269.400 54.900 273.000 ;
        RECT 17.100 265.500 21.900 266.400 ;
        RECT 19.800 264.300 21.900 265.500 ;
        RECT 24.900 264.900 26.100 266.400 ;
        RECT 23.100 262.800 26.100 264.900 ;
        RECT 32.100 264.600 33.300 266.400 ;
        RECT 21.900 259.800 24.000 261.900 ;
        RECT 17.100 256.950 19.200 259.050 ;
        RECT 21.900 258.000 23.700 259.800 ;
        RECT 24.900 257.100 26.100 262.800 ;
        RECT 27.000 263.700 33.300 264.600 ;
        RECT 27.000 261.600 29.100 263.700 ;
        RECT 27.000 259.800 28.800 261.600 ;
        RECT 31.800 259.050 33.600 260.850 ;
        RECT 50.700 259.050 51.900 269.400 ;
        RECT 71.400 266.400 73.200 273.000 ;
        RECT 76.500 265.200 78.300 272.400 ;
        RECT 74.100 264.300 78.300 265.200 ;
        RECT 71.250 259.050 73.050 260.850 ;
        RECT 74.100 259.050 75.300 264.300 ;
        RECT 95.100 263.400 96.900 273.000 ;
        RECT 101.700 264.000 103.500 272.400 ;
        RECT 122.100 264.600 123.900 272.400 ;
        RECT 126.600 266.400 128.400 273.000 ;
        RECT 129.600 268.200 131.400 272.400 ;
        RECT 149.100 269.400 150.900 273.000 ;
        RECT 152.100 269.400 153.900 272.400 ;
        RECT 155.100 269.400 156.900 273.000 ;
        RECT 129.600 266.400 132.300 268.200 ;
        RECT 128.700 264.600 130.500 265.500 ;
        RECT 101.700 262.800 105.000 264.000 ;
        RECT 122.100 263.700 130.500 264.600 ;
        RECT 77.100 259.050 78.900 260.850 ;
        RECT 95.100 259.050 96.900 260.850 ;
        RECT 101.100 259.050 102.900 260.850 ;
        RECT 104.100 259.050 105.000 262.800 ;
        RECT 122.250 259.050 124.050 260.850 ;
        RECT 31.800 258.300 33.900 259.050 ;
        RECT 17.400 255.150 19.200 256.950 ;
        RECT 23.700 256.200 26.100 257.100 ;
        RECT 27.000 256.950 33.900 258.300 ;
        RECT 49.950 256.950 52.050 259.050 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 70.950 256.950 73.050 259.050 ;
        RECT 73.950 256.950 76.050 259.050 ;
        RECT 76.950 256.950 79.050 259.050 ;
        RECT 94.950 256.950 97.050 259.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 122.100 256.950 124.200 259.050 ;
        RECT 27.000 256.500 28.800 256.950 ;
        RECT 23.700 256.050 25.200 256.200 ;
        RECT 23.100 253.950 25.200 256.050 ;
        RECT 24.300 252.000 25.200 253.950 ;
        RECT 26.100 253.500 30.000 255.300 ;
        RECT 26.100 253.200 28.200 253.500 ;
        RECT 24.300 250.950 25.800 252.000 ;
        RECT 19.800 249.600 21.900 250.500 ;
        RECT 17.100 248.400 21.900 249.600 ;
        RECT 24.600 249.600 25.800 250.950 ;
        RECT 29.400 249.600 31.500 251.700 ;
        RECT 17.100 237.600 18.900 248.400 ;
        RECT 20.100 237.000 21.900 247.500 ;
        RECT 24.600 237.600 26.400 249.600 ;
        RECT 29.400 248.700 33.900 249.600 ;
        RECT 29.100 237.000 30.900 247.500 ;
        RECT 32.100 237.600 33.900 248.700 ;
        RECT 50.700 243.600 51.900 256.950 ;
        RECT 53.100 255.150 54.900 256.950 ;
        RECT 74.100 243.600 75.300 256.950 ;
        RECT 98.100 255.150 99.900 256.950 ;
        RECT 104.100 244.800 105.000 256.950 ;
        RECT 98.400 243.900 105.000 244.800 ;
        RECT 98.400 243.600 99.900 243.900 ;
        RECT 50.100 237.600 51.900 243.600 ;
        RECT 53.100 237.000 54.900 243.600 ;
        RECT 71.100 237.000 72.900 243.600 ;
        RECT 74.100 237.600 75.900 243.600 ;
        RECT 77.100 237.000 78.900 243.600 ;
        RECT 95.100 237.000 96.900 243.600 ;
        RECT 98.100 237.600 99.900 243.600 ;
        RECT 104.100 243.600 105.000 243.900 ;
        RECT 125.100 243.600 126.000 263.700 ;
        RECT 131.400 259.050 132.300 266.400 ;
        RECT 152.400 259.050 153.300 269.400 ;
        RECT 173.100 266.400 174.900 272.400 ;
        RECT 173.700 264.300 174.900 266.400 ;
        RECT 176.100 267.300 177.900 272.400 ;
        RECT 179.100 268.200 180.900 273.000 ;
        RECT 182.100 267.300 183.900 272.400 ;
        RECT 176.100 265.950 183.900 267.300 ;
        RECT 200.700 265.200 202.500 272.400 ;
        RECT 205.800 266.400 207.600 273.000 ;
        RECT 224.700 265.200 226.500 272.400 ;
        RECT 229.800 266.400 231.600 273.000 ;
        RECT 248.100 269.400 249.900 272.400 ;
        RECT 251.100 269.400 252.900 273.000 ;
        RECT 269.100 269.400 270.900 273.000 ;
        RECT 272.100 269.400 273.900 272.400 ;
        RECT 275.100 269.400 276.900 273.000 ;
        RECT 293.100 269.400 294.900 272.400 ;
        RECT 296.100 269.400 297.900 273.000 ;
        RECT 200.700 264.300 204.900 265.200 ;
        RECT 224.700 264.300 228.900 265.200 ;
        RECT 173.700 263.400 177.300 264.300 ;
        RECT 160.950 261.450 163.050 262.050 ;
        RECT 169.950 261.450 172.050 262.050 ;
        RECT 160.950 260.550 172.050 261.450 ;
        RECT 160.950 259.950 163.050 260.550 ;
        RECT 169.950 259.950 172.050 260.550 ;
        RECT 173.100 259.050 174.900 260.850 ;
        RECT 176.100 259.050 177.300 263.400 ;
        RECT 179.100 259.050 180.900 260.850 ;
        RECT 200.100 259.050 201.900 260.850 ;
        RECT 203.700 259.050 204.900 264.300 ;
        RECT 205.950 259.050 207.750 260.850 ;
        RECT 224.100 259.050 225.900 260.850 ;
        RECT 227.700 259.050 228.900 264.300 ;
        RECT 232.950 261.450 235.050 262.050 ;
        RECT 244.950 261.450 247.050 262.050 ;
        RECT 229.950 259.050 231.750 260.850 ;
        RECT 232.950 260.550 247.050 261.450 ;
        RECT 232.950 259.950 235.050 260.550 ;
        RECT 244.950 259.950 247.050 260.550 ;
        RECT 248.700 259.050 249.900 269.400 ;
        RECT 272.400 259.050 273.300 269.400 ;
        RECT 293.700 259.050 294.900 269.400 ;
        RECT 314.700 265.200 316.500 272.400 ;
        RECT 319.800 266.400 321.600 273.000 ;
        RECT 323.700 269.400 325.500 273.000 ;
        RECT 326.700 269.400 328.500 272.400 ;
        RECT 314.700 264.300 318.900 265.200 ;
        RECT 314.100 259.050 315.900 260.850 ;
        RECT 317.700 259.050 318.900 264.300 ;
        RECT 319.950 259.050 321.750 260.850 ;
        RECT 127.500 256.950 129.600 259.050 ;
        RECT 130.800 256.950 132.900 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 199.950 256.950 202.050 259.050 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 127.200 255.150 129.000 256.950 ;
        RECT 131.400 249.600 132.300 256.950 ;
        RECT 136.950 255.450 139.050 256.050 ;
        RECT 145.950 255.450 148.050 256.050 ;
        RECT 136.950 254.550 148.050 255.450 ;
        RECT 149.250 255.150 151.050 256.950 ;
        RECT 136.950 253.950 139.050 254.550 ;
        RECT 145.950 253.950 148.050 254.550 ;
        RECT 152.400 249.600 153.300 256.950 ;
        RECT 155.100 255.150 156.900 256.950 ;
        RECT 176.100 249.600 177.300 256.950 ;
        RECT 182.100 255.150 183.900 256.950 ;
        RECT 101.100 237.000 102.900 243.000 ;
        RECT 104.100 237.600 105.900 243.600 ;
        RECT 122.100 237.000 123.900 243.600 ;
        RECT 125.100 237.600 126.900 243.600 ;
        RECT 128.100 237.000 129.900 249.000 ;
        RECT 131.100 237.600 132.900 249.600 ;
        RECT 149.100 237.000 150.900 249.600 ;
        RECT 152.400 248.400 156.000 249.600 ;
        RECT 154.200 237.600 156.000 248.400 ;
        RECT 176.100 248.100 178.500 249.600 ;
        RECT 174.000 245.100 175.800 246.900 ;
        RECT 173.700 237.000 175.500 243.600 ;
        RECT 176.700 237.600 178.500 248.100 ;
        RECT 181.800 237.000 183.600 249.600 ;
        RECT 203.700 243.600 204.900 256.950 ;
        RECT 227.700 243.600 228.900 256.950 ;
        RECT 229.950 252.450 232.050 252.750 ;
        RECT 235.950 252.450 238.050 253.050 ;
        RECT 229.950 251.550 238.050 252.450 ;
        RECT 229.950 250.650 232.050 251.550 ;
        RECT 235.950 250.950 238.050 251.550 ;
        RECT 248.700 243.600 249.900 256.950 ;
        RECT 251.100 255.150 252.900 256.950 ;
        RECT 269.250 255.150 271.050 256.950 ;
        RECT 272.400 249.600 273.300 256.950 ;
        RECT 275.100 255.150 276.900 256.950 ;
        RECT 200.100 237.000 201.900 243.600 ;
        RECT 203.100 237.600 204.900 243.600 ;
        RECT 206.100 237.000 207.900 243.600 ;
        RECT 224.100 237.000 225.900 243.600 ;
        RECT 227.100 237.600 228.900 243.600 ;
        RECT 230.100 237.000 231.900 243.600 ;
        RECT 248.100 237.600 249.900 243.600 ;
        RECT 251.100 237.000 252.900 243.600 ;
        RECT 269.100 237.000 270.900 249.600 ;
        RECT 272.400 248.400 276.000 249.600 ;
        RECT 274.200 237.600 276.000 248.400 ;
        RECT 293.700 243.600 294.900 256.950 ;
        RECT 296.100 255.150 297.900 256.950 ;
        RECT 317.700 243.600 318.900 256.950 ;
        RECT 327.000 256.050 328.500 269.400 ;
        RECT 326.100 253.950 328.500 256.050 ;
        RECT 327.000 243.600 328.500 253.950 ;
        RECT 330.300 266.400 332.100 272.400 ;
        RECT 335.700 266.400 337.500 273.000 ;
        RECT 340.800 267.600 342.600 272.400 ;
        RECT 345.000 269.400 346.800 272.400 ;
        RECT 348.000 269.400 349.800 272.400 ;
        RECT 351.000 269.400 352.800 272.400 ;
        RECT 354.000 269.400 355.800 272.400 ;
        RECT 357.000 269.400 358.800 273.000 ;
        RECT 338.400 266.400 342.600 267.600 ;
        RECT 344.700 267.300 346.800 269.400 ;
        RECT 347.700 267.300 349.800 269.400 ;
        RECT 350.700 267.300 352.800 269.400 ;
        RECT 353.700 267.300 355.800 269.400 ;
        RECT 360.000 268.500 361.800 272.400 ;
        RECT 364.500 269.400 366.300 273.000 ;
        RECT 367.500 269.400 369.300 272.400 ;
        RECT 370.500 269.400 372.300 272.400 ;
        RECT 373.500 269.400 375.300 272.400 ;
        RECT 359.100 266.400 361.800 268.500 ;
        RECT 363.600 267.600 365.400 268.500 ;
        RECT 363.600 266.400 366.300 267.600 ;
        RECT 367.200 267.300 369.300 269.400 ;
        RECT 370.200 267.300 372.300 269.400 ;
        RECT 373.200 267.300 375.300 269.400 ;
        RECT 377.700 266.400 379.500 272.400 ;
        RECT 383.100 266.400 384.900 273.000 ;
        RECT 388.500 266.400 390.300 272.400 ;
        RECT 392.700 269.400 394.500 273.000 ;
        RECT 395.700 269.400 397.500 272.400 ;
        RECT 330.300 249.600 331.200 266.400 ;
        RECT 338.400 263.100 339.900 266.400 ;
        RECT 344.100 264.600 350.700 266.400 ;
        RECT 365.400 265.800 366.300 266.400 ;
        RECT 368.400 265.800 370.200 266.400 ;
        RECT 365.400 264.600 372.600 265.800 ;
        RECT 332.100 261.300 339.900 263.100 ;
        RECT 356.100 262.500 357.900 264.300 ;
        RECT 355.800 261.900 357.900 262.500 ;
        RECT 340.800 260.400 357.900 261.900 ;
        RECT 362.100 261.900 364.200 262.050 ;
        RECT 365.400 261.900 367.200 262.800 ;
        RECT 362.100 261.000 367.200 261.900 ;
        RECT 371.700 261.600 372.600 264.600 ;
        RECT 377.700 265.500 379.200 266.400 ;
        RECT 377.700 264.300 386.100 265.500 ;
        RECT 384.300 263.700 386.100 264.300 ;
        RECT 373.500 262.800 375.600 263.700 ;
        RECT 389.100 262.800 390.300 266.400 ;
        RECT 373.500 261.600 390.300 262.800 ;
        RECT 335.700 258.900 342.300 260.400 ;
        RECT 362.100 259.950 364.200 261.000 ;
        RECT 370.800 259.800 372.600 261.600 ;
        RECT 335.700 256.050 337.200 258.900 ;
        RECT 343.500 257.700 387.900 258.900 ;
        RECT 343.500 256.200 344.400 257.700 ;
        RECT 335.100 253.950 337.200 256.050 ;
        RECT 339.300 254.400 344.400 256.200 ;
        RECT 347.100 255.900 360.600 256.800 ;
        RECT 367.800 255.900 369.600 256.500 ;
        RECT 386.100 256.050 387.900 257.700 ;
        RECT 347.100 254.700 348.000 255.900 ;
        RECT 347.100 252.900 348.900 254.700 ;
        RECT 353.100 253.200 357.000 255.000 ;
        RECT 358.500 254.700 369.600 255.900 ;
        RECT 380.100 255.750 382.200 256.050 ;
        RECT 358.500 253.800 360.600 254.700 ;
        RECT 378.300 253.950 382.200 255.750 ;
        RECT 386.100 253.950 388.200 256.050 ;
        RECT 378.300 253.200 380.100 253.950 ;
        RECT 353.100 252.900 355.200 253.200 ;
        RECT 366.600 252.300 380.100 253.200 ;
        RECT 332.100 251.700 333.900 252.300 ;
        RECT 366.600 251.700 367.800 252.300 ;
        RECT 332.100 250.500 367.800 251.700 ;
        RECT 370.500 250.500 372.600 250.800 ;
        RECT 330.300 248.700 346.800 249.600 ;
        RECT 330.300 245.400 331.200 248.700 ;
        RECT 335.100 246.600 340.800 247.800 ;
        RECT 344.700 247.500 346.800 248.700 ;
        RECT 350.100 248.400 367.800 249.600 ;
        RECT 370.500 249.300 382.500 250.500 ;
        RECT 370.500 248.700 372.600 249.300 ;
        RECT 380.700 248.700 382.500 249.300 ;
        RECT 350.100 247.500 352.200 248.400 ;
        RECT 366.600 247.800 367.800 248.400 ;
        RECT 384.000 247.800 385.800 248.100 ;
        RECT 335.100 246.000 336.900 246.600 ;
        RECT 330.300 244.500 334.200 245.400 ;
        RECT 333.000 243.600 334.200 244.500 ;
        RECT 339.600 243.600 340.800 246.600 ;
        RECT 341.700 245.700 343.500 246.300 ;
        RECT 341.700 244.500 349.800 245.700 ;
        RECT 347.700 243.600 349.800 244.500 ;
        RECT 353.100 243.600 355.800 247.500 ;
        RECT 358.500 245.100 361.800 247.200 ;
        RECT 366.600 246.600 385.800 247.800 ;
        RECT 293.100 237.600 294.900 243.600 ;
        RECT 296.100 237.000 297.900 243.600 ;
        RECT 314.100 237.000 315.900 243.600 ;
        RECT 317.100 237.600 318.900 243.600 ;
        RECT 320.100 237.000 321.900 243.600 ;
        RECT 323.700 237.000 325.500 243.600 ;
        RECT 326.700 237.600 328.500 243.600 ;
        RECT 330.000 237.000 331.800 243.600 ;
        RECT 333.000 237.600 334.800 243.600 ;
        RECT 336.000 237.000 337.800 243.600 ;
        RECT 339.000 237.600 340.800 243.600 ;
        RECT 342.000 237.000 343.800 243.600 ;
        RECT 344.700 240.600 346.800 242.700 ;
        RECT 347.700 240.600 349.800 242.700 ;
        RECT 350.700 240.600 352.800 242.700 ;
        RECT 345.000 237.600 346.800 240.600 ;
        RECT 348.000 237.600 349.800 240.600 ;
        RECT 351.000 237.600 352.800 240.600 ;
        RECT 354.000 237.600 355.800 243.600 ;
        RECT 357.000 237.000 358.800 243.600 ;
        RECT 360.000 237.600 361.800 245.100 ;
        RECT 367.200 243.600 369.300 245.700 ;
        RECT 363.900 237.000 365.700 243.600 ;
        RECT 366.900 237.600 368.700 243.600 ;
        RECT 369.600 240.600 371.700 242.700 ;
        RECT 372.600 240.600 374.700 242.700 ;
        RECT 369.900 237.600 371.700 240.600 ;
        RECT 372.900 237.600 374.700 240.600 ;
        RECT 376.500 237.000 378.300 243.600 ;
        RECT 379.500 237.600 381.300 246.600 ;
        RECT 384.000 246.300 385.800 246.600 ;
        RECT 389.100 245.400 390.300 261.600 ;
        RECT 396.000 256.050 397.500 269.400 ;
        RECT 395.100 253.950 397.500 256.050 ;
        RECT 386.700 244.500 390.300 245.400 ;
        RECT 386.700 243.600 387.600 244.500 ;
        RECT 396.000 243.600 397.500 253.950 ;
        RECT 399.300 266.400 401.100 272.400 ;
        RECT 404.700 266.400 406.500 273.000 ;
        RECT 409.800 267.600 411.600 272.400 ;
        RECT 414.000 269.400 415.800 272.400 ;
        RECT 417.000 269.400 418.800 272.400 ;
        RECT 420.000 269.400 421.800 272.400 ;
        RECT 423.000 269.400 424.800 272.400 ;
        RECT 426.000 269.400 427.800 273.000 ;
        RECT 407.400 266.400 411.600 267.600 ;
        RECT 413.700 267.300 415.800 269.400 ;
        RECT 416.700 267.300 418.800 269.400 ;
        RECT 419.700 267.300 421.800 269.400 ;
        RECT 422.700 267.300 424.800 269.400 ;
        RECT 429.000 268.500 430.800 272.400 ;
        RECT 433.500 269.400 435.300 273.000 ;
        RECT 436.500 269.400 438.300 272.400 ;
        RECT 439.500 269.400 441.300 272.400 ;
        RECT 442.500 269.400 444.300 272.400 ;
        RECT 428.100 266.400 430.800 268.500 ;
        RECT 432.600 267.600 434.400 268.500 ;
        RECT 432.600 266.400 435.300 267.600 ;
        RECT 436.200 267.300 438.300 269.400 ;
        RECT 439.200 267.300 441.300 269.400 ;
        RECT 442.200 267.300 444.300 269.400 ;
        RECT 446.700 266.400 448.500 272.400 ;
        RECT 452.100 266.400 453.900 273.000 ;
        RECT 457.500 266.400 459.300 272.400 ;
        RECT 399.300 249.600 400.200 266.400 ;
        RECT 407.400 263.100 408.900 266.400 ;
        RECT 413.100 264.600 419.700 266.400 ;
        RECT 434.400 265.800 435.300 266.400 ;
        RECT 437.400 265.800 439.200 266.400 ;
        RECT 434.400 264.600 441.600 265.800 ;
        RECT 401.100 261.300 408.900 263.100 ;
        RECT 425.100 262.500 426.900 264.300 ;
        RECT 424.800 261.900 426.900 262.500 ;
        RECT 409.800 260.400 426.900 261.900 ;
        RECT 431.100 261.900 433.200 262.050 ;
        RECT 434.400 261.900 436.200 262.800 ;
        RECT 431.100 261.000 436.200 261.900 ;
        RECT 440.700 261.600 441.600 264.600 ;
        RECT 446.700 265.500 448.200 266.400 ;
        RECT 446.700 264.300 455.100 265.500 ;
        RECT 453.300 263.700 455.100 264.300 ;
        RECT 442.500 262.800 444.600 263.700 ;
        RECT 458.100 262.800 459.300 266.400 ;
        RECT 442.500 261.600 459.300 262.800 ;
        RECT 404.700 258.900 411.300 260.400 ;
        RECT 431.100 259.950 433.200 261.000 ;
        RECT 439.800 259.800 441.600 261.600 ;
        RECT 404.700 256.050 406.200 258.900 ;
        RECT 412.500 257.700 456.900 258.900 ;
        RECT 412.500 256.200 413.400 257.700 ;
        RECT 404.100 253.950 406.200 256.050 ;
        RECT 408.300 254.400 413.400 256.200 ;
        RECT 416.100 255.900 429.600 256.800 ;
        RECT 436.800 255.900 438.600 256.500 ;
        RECT 455.100 256.050 456.900 257.700 ;
        RECT 416.100 254.700 417.000 255.900 ;
        RECT 416.100 252.900 417.900 254.700 ;
        RECT 422.100 253.200 426.000 255.000 ;
        RECT 427.500 254.700 438.600 255.900 ;
        RECT 449.100 255.750 451.200 256.050 ;
        RECT 427.500 253.800 429.600 254.700 ;
        RECT 447.300 253.950 451.200 255.750 ;
        RECT 455.100 253.950 457.200 256.050 ;
        RECT 447.300 253.200 449.100 253.950 ;
        RECT 422.100 252.900 424.200 253.200 ;
        RECT 435.600 252.300 449.100 253.200 ;
        RECT 401.100 251.700 402.900 252.300 ;
        RECT 435.600 251.700 436.800 252.300 ;
        RECT 401.100 250.500 436.800 251.700 ;
        RECT 439.500 250.500 441.600 250.800 ;
        RECT 399.300 248.700 415.800 249.600 ;
        RECT 399.300 245.400 400.200 248.700 ;
        RECT 404.100 246.600 409.800 247.800 ;
        RECT 413.700 247.500 415.800 248.700 ;
        RECT 419.100 248.400 436.800 249.600 ;
        RECT 439.500 249.300 451.500 250.500 ;
        RECT 439.500 248.700 441.600 249.300 ;
        RECT 449.700 248.700 451.500 249.300 ;
        RECT 419.100 247.500 421.200 248.400 ;
        RECT 435.600 247.800 436.800 248.400 ;
        RECT 453.000 247.800 454.800 248.100 ;
        RECT 404.100 246.000 405.900 246.600 ;
        RECT 399.300 244.500 403.200 245.400 ;
        RECT 402.000 243.600 403.200 244.500 ;
        RECT 408.600 243.600 409.800 246.600 ;
        RECT 410.700 245.700 412.500 246.300 ;
        RECT 410.700 244.500 418.800 245.700 ;
        RECT 416.700 243.600 418.800 244.500 ;
        RECT 422.100 243.600 424.800 247.500 ;
        RECT 427.500 245.100 430.800 247.200 ;
        RECT 435.600 246.600 454.800 247.800 ;
        RECT 382.500 237.000 384.300 243.600 ;
        RECT 385.500 242.700 387.600 243.600 ;
        RECT 385.500 237.600 387.300 242.700 ;
        RECT 388.500 237.000 390.300 243.600 ;
        RECT 392.700 237.000 394.500 243.600 ;
        RECT 395.700 237.600 397.500 243.600 ;
        RECT 399.000 237.000 400.800 243.600 ;
        RECT 402.000 237.600 403.800 243.600 ;
        RECT 405.000 237.000 406.800 243.600 ;
        RECT 408.000 237.600 409.800 243.600 ;
        RECT 411.000 237.000 412.800 243.600 ;
        RECT 413.700 240.600 415.800 242.700 ;
        RECT 416.700 240.600 418.800 242.700 ;
        RECT 419.700 240.600 421.800 242.700 ;
        RECT 414.000 237.600 415.800 240.600 ;
        RECT 417.000 237.600 418.800 240.600 ;
        RECT 420.000 237.600 421.800 240.600 ;
        RECT 423.000 237.600 424.800 243.600 ;
        RECT 426.000 237.000 427.800 243.600 ;
        RECT 429.000 237.600 430.800 245.100 ;
        RECT 436.200 243.600 438.300 245.700 ;
        RECT 432.900 237.000 434.700 243.600 ;
        RECT 435.900 237.600 437.700 243.600 ;
        RECT 438.600 240.600 440.700 242.700 ;
        RECT 441.600 240.600 443.700 242.700 ;
        RECT 438.900 237.600 440.700 240.600 ;
        RECT 441.900 237.600 443.700 240.600 ;
        RECT 445.500 237.000 447.300 243.600 ;
        RECT 448.500 237.600 450.300 246.600 ;
        RECT 453.000 246.300 454.800 246.600 ;
        RECT 458.100 245.400 459.300 261.600 ;
        RECT 455.700 244.500 459.300 245.400 ;
        RECT 461.700 266.400 463.500 272.400 ;
        RECT 467.100 266.400 468.900 273.000 ;
        RECT 472.500 266.400 474.300 272.400 ;
        RECT 476.700 269.400 478.500 272.400 ;
        RECT 479.700 269.400 481.500 272.400 ;
        RECT 482.700 269.400 484.500 272.400 ;
        RECT 485.700 269.400 487.500 273.000 ;
        RECT 476.700 267.300 478.800 269.400 ;
        RECT 479.700 267.300 481.800 269.400 ;
        RECT 482.700 267.300 484.800 269.400 ;
        RECT 490.200 268.500 492.000 272.400 ;
        RECT 493.200 269.400 495.000 273.000 ;
        RECT 496.200 269.400 498.000 272.400 ;
        RECT 499.200 269.400 501.000 272.400 ;
        RECT 502.200 269.400 504.000 272.400 ;
        RECT 505.200 269.400 507.000 272.400 ;
        RECT 486.600 267.600 488.400 268.500 ;
        RECT 485.700 266.400 488.400 267.600 ;
        RECT 490.200 266.400 492.900 268.500 ;
        RECT 496.200 267.300 498.300 269.400 ;
        RECT 499.200 267.300 501.300 269.400 ;
        RECT 502.200 267.300 504.300 269.400 ;
        RECT 505.200 267.300 507.300 269.400 ;
        RECT 509.400 267.600 511.200 272.400 ;
        RECT 509.400 266.400 513.600 267.600 ;
        RECT 514.500 266.400 516.300 273.000 ;
        RECT 519.900 266.400 521.700 272.400 ;
        RECT 461.700 262.800 462.900 266.400 ;
        RECT 472.800 265.500 474.300 266.400 ;
        RECT 481.800 265.800 483.600 266.400 ;
        RECT 485.700 265.800 486.600 266.400 ;
        RECT 465.900 264.300 474.300 265.500 ;
        RECT 479.400 264.600 486.600 265.800 ;
        RECT 501.300 264.600 507.900 266.400 ;
        RECT 465.900 263.700 467.700 264.300 ;
        RECT 476.400 262.800 478.500 263.700 ;
        RECT 461.700 261.600 478.500 262.800 ;
        RECT 479.400 261.600 480.300 264.600 ;
        RECT 484.800 261.900 486.600 262.800 ;
        RECT 494.100 262.500 495.900 264.300 ;
        RECT 512.100 263.100 513.600 266.400 ;
        RECT 487.800 261.900 489.900 262.050 ;
        RECT 461.700 245.400 462.900 261.600 ;
        RECT 479.400 259.800 481.200 261.600 ;
        RECT 484.800 261.000 489.900 261.900 ;
        RECT 487.800 259.950 489.900 261.000 ;
        RECT 494.100 261.900 496.200 262.500 ;
        RECT 494.100 260.400 511.200 261.900 ;
        RECT 512.100 261.300 519.900 263.100 ;
        RECT 509.700 258.900 516.300 260.400 ;
        RECT 464.100 257.700 508.500 258.900 ;
        RECT 464.100 256.050 465.900 257.700 ;
        RECT 463.800 253.950 465.900 256.050 ;
        RECT 469.800 255.750 471.900 256.050 ;
        RECT 482.400 255.900 484.200 256.500 ;
        RECT 491.400 255.900 504.900 256.800 ;
        RECT 469.800 253.950 473.700 255.750 ;
        RECT 482.400 254.700 493.500 255.900 ;
        RECT 471.900 253.200 473.700 253.950 ;
        RECT 491.400 253.800 493.500 254.700 ;
        RECT 495.000 253.200 498.900 255.000 ;
        RECT 504.000 254.700 504.900 255.900 ;
        RECT 471.900 252.300 485.400 253.200 ;
        RECT 496.800 252.900 498.900 253.200 ;
        RECT 503.100 252.900 504.900 254.700 ;
        RECT 507.600 256.200 508.500 257.700 ;
        RECT 507.600 254.400 512.700 256.200 ;
        RECT 514.800 256.050 516.300 258.900 ;
        RECT 514.800 253.950 516.900 256.050 ;
        RECT 484.200 251.700 485.400 252.300 ;
        RECT 518.100 251.700 519.900 252.300 ;
        RECT 479.400 250.500 481.500 250.800 ;
        RECT 484.200 250.500 519.900 251.700 ;
        RECT 469.500 249.300 481.500 250.500 ;
        RECT 520.800 249.600 521.700 266.400 ;
        RECT 469.500 248.700 471.300 249.300 ;
        RECT 479.400 248.700 481.500 249.300 ;
        RECT 484.200 248.400 501.900 249.600 ;
        RECT 466.200 247.800 468.000 248.100 ;
        RECT 484.200 247.800 485.400 248.400 ;
        RECT 466.200 246.600 485.400 247.800 ;
        RECT 499.800 247.500 501.900 248.400 ;
        RECT 505.200 248.700 521.700 249.600 ;
        RECT 505.200 247.500 507.300 248.700 ;
        RECT 466.200 246.300 468.000 246.600 ;
        RECT 461.700 244.500 465.300 245.400 ;
        RECT 455.700 243.600 456.600 244.500 ;
        RECT 464.400 243.600 465.300 244.500 ;
        RECT 451.500 237.000 453.300 243.600 ;
        RECT 454.500 242.700 456.600 243.600 ;
        RECT 454.500 237.600 456.300 242.700 ;
        RECT 457.500 237.000 459.300 243.600 ;
        RECT 461.700 237.000 463.500 243.600 ;
        RECT 464.400 242.700 466.500 243.600 ;
        RECT 464.700 237.600 466.500 242.700 ;
        RECT 467.700 237.000 469.500 243.600 ;
        RECT 470.700 237.600 472.500 246.600 ;
        RECT 482.700 243.600 484.800 245.700 ;
        RECT 490.200 245.100 493.500 247.200 ;
        RECT 473.700 237.000 475.500 243.600 ;
        RECT 477.300 240.600 479.400 242.700 ;
        RECT 480.300 240.600 482.400 242.700 ;
        RECT 477.300 237.600 479.100 240.600 ;
        RECT 480.300 237.600 482.100 240.600 ;
        RECT 483.300 237.600 485.100 243.600 ;
        RECT 486.300 237.000 488.100 243.600 ;
        RECT 490.200 237.600 492.000 245.100 ;
        RECT 496.200 243.600 498.900 247.500 ;
        RECT 511.200 246.600 516.900 247.800 ;
        RECT 508.500 245.700 510.300 246.300 ;
        RECT 502.200 244.500 510.300 245.700 ;
        RECT 502.200 243.600 504.300 244.500 ;
        RECT 511.200 243.600 512.400 246.600 ;
        RECT 515.100 246.000 516.900 246.600 ;
        RECT 520.800 245.400 521.700 248.700 ;
        RECT 517.800 244.500 521.700 245.400 ;
        RECT 523.500 269.400 525.300 272.400 ;
        RECT 526.500 269.400 528.300 273.000 ;
        RECT 523.500 256.050 525.000 269.400 ;
        RECT 545.400 266.400 547.200 273.000 ;
        RECT 550.500 265.200 552.300 272.400 ;
        RECT 569.100 269.400 570.900 273.000 ;
        RECT 572.100 269.400 573.900 272.400 ;
        RECT 590.100 269.400 591.900 273.000 ;
        RECT 593.100 269.400 594.900 272.400 ;
        RECT 548.100 264.300 552.300 265.200 ;
        RECT 556.950 264.450 559.050 265.050 ;
        RECT 568.950 264.450 571.050 265.050 ;
        RECT 545.250 259.050 547.050 260.850 ;
        RECT 548.100 259.050 549.300 264.300 ;
        RECT 556.950 263.550 571.050 264.450 ;
        RECT 556.950 262.950 559.050 263.550 ;
        RECT 568.950 262.950 571.050 263.550 ;
        RECT 551.100 259.050 552.900 260.850 ;
        RECT 572.100 259.050 573.300 269.400 ;
        RECT 574.950 267.450 577.050 268.050 ;
        RECT 580.950 267.450 583.050 268.050 ;
        RECT 574.950 266.550 583.050 267.450 ;
        RECT 574.950 265.950 577.050 266.550 ;
        RECT 580.950 265.950 583.050 266.550 ;
        RECT 593.100 259.050 594.300 269.400 ;
        RECT 611.400 266.400 613.200 273.000 ;
        RECT 616.500 265.200 618.300 272.400 ;
        RECT 635.100 266.400 636.900 272.400 ;
        RECT 614.100 264.300 618.300 265.200 ;
        RECT 635.700 264.300 636.900 266.400 ;
        RECT 638.100 267.300 639.900 272.400 ;
        RECT 641.100 268.200 642.900 273.000 ;
        RECT 644.100 267.300 645.900 272.400 ;
        RECT 638.100 265.950 645.900 267.300 ;
        RECT 662.100 267.300 663.900 272.400 ;
        RECT 665.100 268.200 666.900 273.000 ;
        RECT 668.100 267.300 669.900 272.400 ;
        RECT 662.100 265.950 669.900 267.300 ;
        RECT 671.100 266.400 672.900 272.400 ;
        RECT 674.700 269.400 676.500 273.000 ;
        RECT 677.700 269.400 679.500 272.400 ;
        RECT 671.100 264.300 672.300 266.400 ;
        RECT 611.250 259.050 613.050 260.850 ;
        RECT 614.100 259.050 615.300 264.300 ;
        RECT 635.700 263.400 639.300 264.300 ;
        RECT 617.100 259.050 618.900 260.850 ;
        RECT 635.100 259.050 636.900 260.850 ;
        RECT 638.100 259.050 639.300 263.400 ;
        RECT 668.700 263.400 672.300 264.300 ;
        RECT 641.100 259.050 642.900 260.850 ;
        RECT 665.100 259.050 666.900 260.850 ;
        RECT 668.700 259.050 669.900 263.400 ;
        RECT 671.100 259.050 672.900 260.850 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 640.950 256.950 643.050 259.050 ;
        RECT 643.950 256.950 646.050 259.050 ;
        RECT 661.950 256.950 664.050 259.050 ;
        RECT 664.950 256.950 667.050 259.050 ;
        RECT 667.950 256.950 670.050 259.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 523.500 253.950 525.900 256.050 ;
        RECT 517.800 243.600 519.000 244.500 ;
        RECT 523.500 243.600 525.000 253.950 ;
        RECT 548.100 243.600 549.300 256.950 ;
        RECT 569.100 255.150 570.900 256.950 ;
        RECT 572.100 243.600 573.300 256.950 ;
        RECT 590.100 255.150 591.900 256.950 ;
        RECT 593.100 243.600 594.300 256.950 ;
        RECT 614.100 243.600 615.300 256.950 ;
        RECT 638.100 249.600 639.300 256.950 ;
        RECT 644.100 255.150 645.900 256.950 ;
        RECT 662.100 255.150 663.900 256.950 ;
        RECT 668.700 249.600 669.900 256.950 ;
        RECT 678.000 256.050 679.500 269.400 ;
        RECT 677.100 253.950 679.500 256.050 ;
        RECT 638.100 248.100 640.500 249.600 ;
        RECT 636.000 245.100 637.800 246.900 ;
        RECT 493.200 237.000 495.000 243.600 ;
        RECT 496.200 237.600 498.000 243.600 ;
        RECT 499.200 240.600 501.300 242.700 ;
        RECT 502.200 240.600 504.300 242.700 ;
        RECT 505.200 240.600 507.300 242.700 ;
        RECT 499.200 237.600 501.000 240.600 ;
        RECT 502.200 237.600 504.000 240.600 ;
        RECT 505.200 237.600 507.000 240.600 ;
        RECT 508.200 237.000 510.000 243.600 ;
        RECT 511.200 237.600 513.000 243.600 ;
        RECT 514.200 237.000 516.000 243.600 ;
        RECT 517.200 237.600 519.000 243.600 ;
        RECT 520.200 237.000 522.000 243.600 ;
        RECT 523.500 237.600 525.300 243.600 ;
        RECT 526.500 237.000 528.300 243.600 ;
        RECT 545.100 237.000 546.900 243.600 ;
        RECT 548.100 237.600 549.900 243.600 ;
        RECT 551.100 237.000 552.900 243.600 ;
        RECT 569.100 237.000 570.900 243.600 ;
        RECT 572.100 237.600 573.900 243.600 ;
        RECT 590.100 237.000 591.900 243.600 ;
        RECT 593.100 237.600 594.900 243.600 ;
        RECT 611.100 237.000 612.900 243.600 ;
        RECT 614.100 237.600 615.900 243.600 ;
        RECT 617.100 237.000 618.900 243.600 ;
        RECT 635.700 237.000 637.500 243.600 ;
        RECT 638.700 237.600 640.500 248.100 ;
        RECT 643.800 237.000 645.600 249.600 ;
        RECT 662.400 237.000 664.200 249.600 ;
        RECT 667.500 248.100 669.900 249.600 ;
        RECT 667.500 237.600 669.300 248.100 ;
        RECT 670.200 245.100 672.000 246.900 ;
        RECT 678.000 243.600 679.500 253.950 ;
        RECT 681.300 266.400 683.100 272.400 ;
        RECT 686.700 266.400 688.500 273.000 ;
        RECT 691.800 267.600 693.600 272.400 ;
        RECT 696.000 269.400 697.800 272.400 ;
        RECT 699.000 269.400 700.800 272.400 ;
        RECT 702.000 269.400 703.800 272.400 ;
        RECT 705.000 269.400 706.800 272.400 ;
        RECT 708.000 269.400 709.800 273.000 ;
        RECT 689.400 266.400 693.600 267.600 ;
        RECT 695.700 267.300 697.800 269.400 ;
        RECT 698.700 267.300 700.800 269.400 ;
        RECT 701.700 267.300 703.800 269.400 ;
        RECT 704.700 267.300 706.800 269.400 ;
        RECT 711.000 268.500 712.800 272.400 ;
        RECT 715.500 269.400 717.300 273.000 ;
        RECT 718.500 269.400 720.300 272.400 ;
        RECT 721.500 269.400 723.300 272.400 ;
        RECT 724.500 269.400 726.300 272.400 ;
        RECT 710.100 266.400 712.800 268.500 ;
        RECT 714.600 267.600 716.400 268.500 ;
        RECT 714.600 266.400 717.300 267.600 ;
        RECT 718.200 267.300 720.300 269.400 ;
        RECT 721.200 267.300 723.300 269.400 ;
        RECT 724.200 267.300 726.300 269.400 ;
        RECT 728.700 266.400 730.500 272.400 ;
        RECT 734.100 266.400 735.900 273.000 ;
        RECT 739.500 266.400 741.300 272.400 ;
        RECT 758.100 266.400 759.900 272.400 ;
        RECT 761.100 267.300 762.900 273.000 ;
        RECT 765.600 266.400 767.400 272.400 ;
        RECT 770.100 267.300 771.900 273.000 ;
        RECT 773.100 266.400 774.900 272.400 ;
        RECT 791.100 269.400 792.900 273.000 ;
        RECT 794.100 269.400 795.900 272.400 ;
        RECT 812.100 269.400 813.900 273.000 ;
        RECT 815.100 269.400 816.900 272.400 ;
        RECT 818.100 269.400 819.900 273.000 ;
        RECT 681.300 249.600 682.200 266.400 ;
        RECT 689.400 263.100 690.900 266.400 ;
        RECT 695.100 264.600 701.700 266.400 ;
        RECT 716.400 265.800 717.300 266.400 ;
        RECT 719.400 265.800 721.200 266.400 ;
        RECT 716.400 264.600 723.600 265.800 ;
        RECT 683.100 261.300 690.900 263.100 ;
        RECT 707.100 262.500 708.900 264.300 ;
        RECT 706.800 261.900 708.900 262.500 ;
        RECT 691.800 260.400 708.900 261.900 ;
        RECT 713.100 261.900 715.200 262.050 ;
        RECT 716.400 261.900 718.200 262.800 ;
        RECT 713.100 261.000 718.200 261.900 ;
        RECT 722.700 261.600 723.600 264.600 ;
        RECT 728.700 265.500 730.200 266.400 ;
        RECT 728.700 264.300 737.100 265.500 ;
        RECT 735.300 263.700 737.100 264.300 ;
        RECT 724.500 262.800 726.600 263.700 ;
        RECT 740.100 262.800 741.300 266.400 ;
        RECT 758.700 264.600 759.900 266.400 ;
        RECT 765.900 264.900 767.100 266.400 ;
        RECT 770.100 265.500 774.900 266.400 ;
        RECT 758.700 263.700 765.000 264.600 ;
        RECT 724.500 261.600 741.300 262.800 ;
        RECT 762.900 261.600 765.000 263.700 ;
        RECT 686.700 258.900 693.300 260.400 ;
        RECT 713.100 259.950 715.200 261.000 ;
        RECT 721.800 259.800 723.600 261.600 ;
        RECT 686.700 256.050 688.200 258.900 ;
        RECT 694.500 257.700 738.900 258.900 ;
        RECT 694.500 256.200 695.400 257.700 ;
        RECT 686.100 253.950 688.200 256.050 ;
        RECT 690.300 254.400 695.400 256.200 ;
        RECT 698.100 255.900 711.600 256.800 ;
        RECT 718.800 255.900 720.600 256.500 ;
        RECT 737.100 256.050 738.900 257.700 ;
        RECT 698.100 254.700 699.000 255.900 ;
        RECT 698.100 252.900 699.900 254.700 ;
        RECT 704.100 253.200 708.000 255.000 ;
        RECT 709.500 254.700 720.600 255.900 ;
        RECT 731.100 255.750 733.200 256.050 ;
        RECT 709.500 253.800 711.600 254.700 ;
        RECT 729.300 253.950 733.200 255.750 ;
        RECT 737.100 253.950 739.200 256.050 ;
        RECT 729.300 253.200 731.100 253.950 ;
        RECT 704.100 252.900 706.200 253.200 ;
        RECT 717.600 252.300 731.100 253.200 ;
        RECT 683.100 251.700 684.900 252.300 ;
        RECT 717.600 251.700 718.800 252.300 ;
        RECT 683.100 250.500 718.800 251.700 ;
        RECT 721.500 250.500 723.600 250.800 ;
        RECT 681.300 248.700 697.800 249.600 ;
        RECT 681.300 245.400 682.200 248.700 ;
        RECT 686.100 246.600 691.800 247.800 ;
        RECT 695.700 247.500 697.800 248.700 ;
        RECT 701.100 248.400 718.800 249.600 ;
        RECT 721.500 249.300 733.500 250.500 ;
        RECT 721.500 248.700 723.600 249.300 ;
        RECT 731.700 248.700 733.500 249.300 ;
        RECT 701.100 247.500 703.200 248.400 ;
        RECT 717.600 247.800 718.800 248.400 ;
        RECT 735.000 247.800 736.800 248.100 ;
        RECT 686.100 246.000 687.900 246.600 ;
        RECT 681.300 244.500 685.200 245.400 ;
        RECT 684.000 243.600 685.200 244.500 ;
        RECT 690.600 243.600 691.800 246.600 ;
        RECT 692.700 245.700 694.500 246.300 ;
        RECT 692.700 244.500 700.800 245.700 ;
        RECT 698.700 243.600 700.800 244.500 ;
        RECT 704.100 243.600 706.800 247.500 ;
        RECT 709.500 245.100 712.800 247.200 ;
        RECT 717.600 246.600 736.800 247.800 ;
        RECT 670.500 237.000 672.300 243.600 ;
        RECT 674.700 237.000 676.500 243.600 ;
        RECT 677.700 237.600 679.500 243.600 ;
        RECT 681.000 237.000 682.800 243.600 ;
        RECT 684.000 237.600 685.800 243.600 ;
        RECT 687.000 237.000 688.800 243.600 ;
        RECT 690.000 237.600 691.800 243.600 ;
        RECT 693.000 237.000 694.800 243.600 ;
        RECT 695.700 240.600 697.800 242.700 ;
        RECT 698.700 240.600 700.800 242.700 ;
        RECT 701.700 240.600 703.800 242.700 ;
        RECT 696.000 237.600 697.800 240.600 ;
        RECT 699.000 237.600 700.800 240.600 ;
        RECT 702.000 237.600 703.800 240.600 ;
        RECT 705.000 237.600 706.800 243.600 ;
        RECT 708.000 237.000 709.800 243.600 ;
        RECT 711.000 237.600 712.800 245.100 ;
        RECT 718.200 243.600 720.300 245.700 ;
        RECT 714.900 237.000 716.700 243.600 ;
        RECT 717.900 237.600 719.700 243.600 ;
        RECT 720.600 240.600 722.700 242.700 ;
        RECT 723.600 240.600 725.700 242.700 ;
        RECT 720.900 237.600 722.700 240.600 ;
        RECT 723.900 237.600 725.700 240.600 ;
        RECT 727.500 237.000 729.300 243.600 ;
        RECT 730.500 237.600 732.300 246.600 ;
        RECT 735.000 246.300 736.800 246.600 ;
        RECT 740.100 245.400 741.300 261.600 ;
        RECT 758.400 259.050 760.200 260.850 ;
        RECT 763.200 259.800 765.000 261.600 ;
        RECT 765.900 262.800 768.900 264.900 ;
        RECT 770.100 264.300 772.200 265.500 ;
        RECT 758.100 258.300 760.200 259.050 ;
        RECT 758.100 256.950 765.000 258.300 ;
        RECT 763.200 256.500 765.000 256.950 ;
        RECT 765.900 257.100 767.100 262.800 ;
        RECT 768.000 259.800 770.100 261.900 ;
        RECT 768.300 258.000 770.100 259.800 ;
        RECT 794.100 259.050 795.300 269.400 ;
        RECT 815.400 259.050 816.300 269.400 ;
        RECT 821.700 266.400 823.500 272.400 ;
        RECT 827.100 266.400 828.900 273.000 ;
        RECT 832.500 266.400 834.300 272.400 ;
        RECT 836.700 269.400 838.500 272.400 ;
        RECT 839.700 269.400 841.500 272.400 ;
        RECT 842.700 269.400 844.500 272.400 ;
        RECT 845.700 269.400 847.500 273.000 ;
        RECT 836.700 267.300 838.800 269.400 ;
        RECT 839.700 267.300 841.800 269.400 ;
        RECT 842.700 267.300 844.800 269.400 ;
        RECT 850.200 268.500 852.000 272.400 ;
        RECT 853.200 269.400 855.000 273.000 ;
        RECT 856.200 269.400 858.000 272.400 ;
        RECT 859.200 269.400 861.000 272.400 ;
        RECT 862.200 269.400 864.000 272.400 ;
        RECT 865.200 269.400 867.000 272.400 ;
        RECT 846.600 267.600 848.400 268.500 ;
        RECT 845.700 266.400 848.400 267.600 ;
        RECT 850.200 266.400 852.900 268.500 ;
        RECT 856.200 267.300 858.300 269.400 ;
        RECT 859.200 267.300 861.300 269.400 ;
        RECT 862.200 267.300 864.300 269.400 ;
        RECT 865.200 267.300 867.300 269.400 ;
        RECT 869.400 267.600 871.200 272.400 ;
        RECT 869.400 266.400 873.600 267.600 ;
        RECT 874.500 266.400 876.300 273.000 ;
        RECT 879.900 266.400 881.700 272.400 ;
        RECT 821.700 262.800 822.900 266.400 ;
        RECT 832.800 265.500 834.300 266.400 ;
        RECT 841.800 265.800 843.600 266.400 ;
        RECT 845.700 265.800 846.600 266.400 ;
        RECT 825.900 264.300 834.300 265.500 ;
        RECT 839.400 264.600 846.600 265.800 ;
        RECT 861.300 264.600 867.900 266.400 ;
        RECT 825.900 263.700 827.700 264.300 ;
        RECT 836.400 262.800 838.500 263.700 ;
        RECT 821.700 261.600 838.500 262.800 ;
        RECT 839.400 261.600 840.300 264.600 ;
        RECT 844.800 261.900 846.600 262.800 ;
        RECT 854.100 262.500 855.900 264.300 ;
        RECT 872.100 263.100 873.600 266.400 ;
        RECT 847.800 261.900 849.900 262.050 ;
        RECT 765.900 256.200 768.300 257.100 ;
        RECT 766.800 256.050 768.300 256.200 ;
        RECT 772.800 256.950 774.900 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 762.000 253.500 765.900 255.300 ;
        RECT 763.800 253.200 765.900 253.500 ;
        RECT 766.800 253.950 768.900 256.050 ;
        RECT 772.800 255.150 774.600 256.950 ;
        RECT 791.100 255.150 792.900 256.950 ;
        RECT 766.800 252.000 767.700 253.950 ;
        RECT 760.500 249.600 762.600 251.700 ;
        RECT 766.200 250.950 767.700 252.000 ;
        RECT 766.200 249.600 767.400 250.950 ;
        RECT 737.700 244.500 741.300 245.400 ;
        RECT 758.100 248.700 762.600 249.600 ;
        RECT 737.700 243.600 738.600 244.500 ;
        RECT 733.500 237.000 735.300 243.600 ;
        RECT 736.500 242.700 738.600 243.600 ;
        RECT 736.500 237.600 738.300 242.700 ;
        RECT 739.500 237.000 741.300 243.600 ;
        RECT 758.100 237.600 759.900 248.700 ;
        RECT 761.100 237.000 762.900 247.500 ;
        RECT 765.600 237.600 767.400 249.600 ;
        RECT 770.100 249.600 772.200 250.500 ;
        RECT 770.100 248.400 774.900 249.600 ;
        RECT 770.100 237.000 771.900 247.500 ;
        RECT 773.100 237.600 774.900 248.400 ;
        RECT 794.100 243.600 795.300 256.950 ;
        RECT 812.250 255.150 814.050 256.950 ;
        RECT 815.400 249.600 816.300 256.950 ;
        RECT 818.100 255.150 819.900 256.950 ;
        RECT 791.100 237.000 792.900 243.600 ;
        RECT 794.100 237.600 795.900 243.600 ;
        RECT 812.100 237.000 813.900 249.600 ;
        RECT 815.400 248.400 819.000 249.600 ;
        RECT 817.200 237.600 819.000 248.400 ;
        RECT 821.700 245.400 822.900 261.600 ;
        RECT 839.400 259.800 841.200 261.600 ;
        RECT 844.800 261.000 849.900 261.900 ;
        RECT 847.800 259.950 849.900 261.000 ;
        RECT 854.100 261.900 856.200 262.500 ;
        RECT 854.100 260.400 871.200 261.900 ;
        RECT 872.100 261.300 879.900 263.100 ;
        RECT 869.700 258.900 876.300 260.400 ;
        RECT 824.100 257.700 868.500 258.900 ;
        RECT 824.100 256.050 825.900 257.700 ;
        RECT 823.800 253.950 825.900 256.050 ;
        RECT 829.800 255.750 831.900 256.050 ;
        RECT 842.400 255.900 844.200 256.500 ;
        RECT 851.400 255.900 864.900 256.800 ;
        RECT 829.800 253.950 833.700 255.750 ;
        RECT 842.400 254.700 853.500 255.900 ;
        RECT 831.900 253.200 833.700 253.950 ;
        RECT 851.400 253.800 853.500 254.700 ;
        RECT 855.000 253.200 858.900 255.000 ;
        RECT 864.000 254.700 864.900 255.900 ;
        RECT 831.900 252.300 845.400 253.200 ;
        RECT 856.800 252.900 858.900 253.200 ;
        RECT 863.100 252.900 864.900 254.700 ;
        RECT 867.600 256.200 868.500 257.700 ;
        RECT 867.600 254.400 872.700 256.200 ;
        RECT 874.800 256.050 876.300 258.900 ;
        RECT 874.800 253.950 876.900 256.050 ;
        RECT 844.200 251.700 845.400 252.300 ;
        RECT 878.100 251.700 879.900 252.300 ;
        RECT 839.400 250.500 841.500 250.800 ;
        RECT 844.200 250.500 879.900 251.700 ;
        RECT 829.500 249.300 841.500 250.500 ;
        RECT 880.800 249.600 881.700 266.400 ;
        RECT 829.500 248.700 831.300 249.300 ;
        RECT 839.400 248.700 841.500 249.300 ;
        RECT 844.200 248.400 861.900 249.600 ;
        RECT 826.200 247.800 828.000 248.100 ;
        RECT 844.200 247.800 845.400 248.400 ;
        RECT 826.200 246.600 845.400 247.800 ;
        RECT 859.800 247.500 861.900 248.400 ;
        RECT 865.200 248.700 881.700 249.600 ;
        RECT 865.200 247.500 867.300 248.700 ;
        RECT 826.200 246.300 828.000 246.600 ;
        RECT 821.700 244.500 825.300 245.400 ;
        RECT 824.400 243.600 825.300 244.500 ;
        RECT 821.700 237.000 823.500 243.600 ;
        RECT 824.400 242.700 826.500 243.600 ;
        RECT 824.700 237.600 826.500 242.700 ;
        RECT 827.700 237.000 829.500 243.600 ;
        RECT 830.700 237.600 832.500 246.600 ;
        RECT 842.700 243.600 844.800 245.700 ;
        RECT 850.200 245.100 853.500 247.200 ;
        RECT 833.700 237.000 835.500 243.600 ;
        RECT 837.300 240.600 839.400 242.700 ;
        RECT 840.300 240.600 842.400 242.700 ;
        RECT 837.300 237.600 839.100 240.600 ;
        RECT 840.300 237.600 842.100 240.600 ;
        RECT 843.300 237.600 845.100 243.600 ;
        RECT 846.300 237.000 848.100 243.600 ;
        RECT 850.200 237.600 852.000 245.100 ;
        RECT 856.200 243.600 858.900 247.500 ;
        RECT 871.200 246.600 876.900 247.800 ;
        RECT 868.500 245.700 870.300 246.300 ;
        RECT 862.200 244.500 870.300 245.700 ;
        RECT 862.200 243.600 864.300 244.500 ;
        RECT 871.200 243.600 872.400 246.600 ;
        RECT 875.100 246.000 876.900 246.600 ;
        RECT 880.800 245.400 881.700 248.700 ;
        RECT 877.800 244.500 881.700 245.400 ;
        RECT 883.500 269.400 885.300 272.400 ;
        RECT 886.500 269.400 888.300 273.000 ;
        RECT 883.500 256.050 885.000 269.400 ;
        RECT 907.500 264.000 909.300 272.400 ;
        RECT 906.000 262.800 909.300 264.000 ;
        RECT 914.100 263.400 915.900 273.000 ;
        RECT 932.400 266.400 934.200 273.000 ;
        RECT 937.500 265.200 939.300 272.400 ;
        RECT 931.950 264.450 934.050 265.050 ;
        RECT 926.550 263.550 934.050 264.450 ;
        RECT 886.950 261.450 889.050 262.050 ;
        RECT 901.950 261.450 904.050 262.050 ;
        RECT 886.950 260.550 904.050 261.450 ;
        RECT 886.950 259.950 889.050 260.550 ;
        RECT 901.950 259.950 904.050 260.550 ;
        RECT 906.000 259.050 906.900 262.800 ;
        RECT 908.100 259.050 909.900 260.850 ;
        RECT 914.100 259.050 915.900 260.850 ;
        RECT 904.950 256.950 907.050 259.050 ;
        RECT 907.950 256.950 910.050 259.050 ;
        RECT 910.950 256.950 913.050 259.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 883.500 253.950 885.900 256.050 ;
        RECT 877.800 243.600 879.000 244.500 ;
        RECT 883.500 243.600 885.000 253.950 ;
        RECT 906.000 244.800 906.900 256.950 ;
        RECT 911.100 255.150 912.900 256.950 ;
        RECT 926.550 256.050 927.450 263.550 ;
        RECT 931.950 262.950 934.050 263.550 ;
        RECT 935.100 264.300 939.300 265.200 ;
        RECT 932.250 259.050 934.050 260.850 ;
        RECT 935.100 259.050 936.300 264.300 ;
        RECT 958.500 264.000 960.300 272.400 ;
        RECT 957.000 262.800 960.300 264.000 ;
        RECT 965.100 263.400 966.900 273.000 ;
        RECT 983.100 266.400 984.900 272.400 ;
        RECT 986.100 266.400 987.900 273.000 ;
        RECT 1004.100 266.400 1005.900 272.400 ;
        RECT 938.100 259.050 939.900 260.850 ;
        RECT 957.000 259.050 957.900 262.800 ;
        RECT 959.100 259.050 960.900 260.850 ;
        RECT 965.100 259.050 966.900 260.850 ;
        RECT 983.700 259.050 984.900 266.400 ;
        RECT 1004.700 264.300 1005.900 266.400 ;
        RECT 1007.100 267.300 1008.900 272.400 ;
        RECT 1010.100 268.200 1011.900 273.000 ;
        RECT 1013.100 267.300 1014.900 272.400 ;
        RECT 1007.100 265.950 1014.900 267.300 ;
        RECT 1031.100 266.400 1032.900 272.400 ;
        RECT 1015.950 264.450 1018.050 265.050 ;
        RECT 1004.700 263.400 1008.300 264.300 ;
        RECT 999.000 261.450 1003.050 262.050 ;
        RECT 986.100 259.050 987.900 260.850 ;
        RECT 998.550 259.950 1003.050 261.450 ;
        RECT 931.950 256.950 934.050 259.050 ;
        RECT 934.950 256.950 937.050 259.050 ;
        RECT 937.950 256.950 940.050 259.050 ;
        RECT 955.950 256.950 958.050 259.050 ;
        RECT 958.950 256.950 961.050 259.050 ;
        RECT 961.950 256.950 964.050 259.050 ;
        RECT 964.950 256.950 967.050 259.050 ;
        RECT 982.950 256.950 985.050 259.050 ;
        RECT 985.950 256.950 988.050 259.050 ;
        RECT 926.550 254.550 931.050 256.050 ;
        RECT 927.000 253.950 931.050 254.550 ;
        RECT 906.000 243.900 912.600 244.800 ;
        RECT 906.000 243.600 906.900 243.900 ;
        RECT 853.200 237.000 855.000 243.600 ;
        RECT 856.200 237.600 858.000 243.600 ;
        RECT 859.200 240.600 861.300 242.700 ;
        RECT 862.200 240.600 864.300 242.700 ;
        RECT 865.200 240.600 867.300 242.700 ;
        RECT 859.200 237.600 861.000 240.600 ;
        RECT 862.200 237.600 864.000 240.600 ;
        RECT 865.200 237.600 867.000 240.600 ;
        RECT 868.200 237.000 870.000 243.600 ;
        RECT 871.200 237.600 873.000 243.600 ;
        RECT 874.200 237.000 876.000 243.600 ;
        RECT 877.200 237.600 879.000 243.600 ;
        RECT 880.200 237.000 882.000 243.600 ;
        RECT 883.500 237.600 885.300 243.600 ;
        RECT 886.500 237.000 888.300 243.600 ;
        RECT 905.100 237.600 906.900 243.600 ;
        RECT 911.100 243.600 912.600 243.900 ;
        RECT 935.100 243.600 936.300 256.950 ;
        RECT 957.000 244.800 957.900 256.950 ;
        RECT 962.100 255.150 963.900 256.950 ;
        RECT 958.950 252.450 961.050 253.050 ;
        RECT 973.950 252.450 976.050 253.050 ;
        RECT 958.950 251.550 976.050 252.450 ;
        RECT 958.950 250.950 961.050 251.550 ;
        RECT 973.950 250.950 976.050 251.550 ;
        RECT 983.700 249.600 984.900 256.950 ;
        RECT 998.550 256.050 999.450 259.950 ;
        RECT 1004.100 259.050 1005.900 260.850 ;
        RECT 1007.100 259.050 1008.300 263.400 ;
        RECT 1015.950 263.550 1026.450 264.450 ;
        RECT 1015.950 262.950 1018.050 263.550 ;
        RECT 1010.100 259.050 1011.900 260.850 ;
        RECT 1003.950 256.950 1006.050 259.050 ;
        RECT 1006.950 256.950 1009.050 259.050 ;
        RECT 1009.950 256.950 1012.050 259.050 ;
        RECT 1012.950 256.950 1015.050 259.050 ;
        RECT 998.550 254.550 1003.050 256.050 ;
        RECT 999.000 253.950 1003.050 254.550 ;
        RECT 985.950 252.450 988.050 253.050 ;
        RECT 994.950 252.450 997.050 253.050 ;
        RECT 985.950 251.550 997.050 252.450 ;
        RECT 985.950 250.950 988.050 251.550 ;
        RECT 994.950 250.950 997.050 251.550 ;
        RECT 1007.100 249.600 1008.300 256.950 ;
        RECT 1013.100 255.150 1014.900 256.950 ;
        RECT 1025.550 256.050 1026.450 263.550 ;
        RECT 1031.700 264.300 1032.900 266.400 ;
        RECT 1034.100 267.300 1035.900 272.400 ;
        RECT 1037.100 268.200 1038.900 273.000 ;
        RECT 1040.100 267.300 1041.900 272.400 ;
        RECT 1034.100 265.950 1041.900 267.300 ;
        RECT 1031.700 263.400 1035.300 264.300 ;
        RECT 1031.100 259.050 1032.900 260.850 ;
        RECT 1034.100 259.050 1035.300 263.400 ;
        RECT 1037.100 259.050 1038.900 260.850 ;
        RECT 1030.950 256.950 1033.050 259.050 ;
        RECT 1033.950 256.950 1036.050 259.050 ;
        RECT 1036.950 256.950 1039.050 259.050 ;
        RECT 1039.950 256.950 1042.050 259.050 ;
        RECT 1025.550 254.550 1030.050 256.050 ;
        RECT 1026.000 253.950 1030.050 254.550 ;
        RECT 1034.100 249.600 1035.300 256.950 ;
        RECT 1040.100 255.150 1041.900 256.950 ;
        RECT 957.000 243.900 963.600 244.800 ;
        RECT 957.000 243.600 957.900 243.900 ;
        RECT 908.100 237.000 909.900 243.000 ;
        RECT 911.100 237.600 912.900 243.600 ;
        RECT 914.100 237.000 915.900 243.600 ;
        RECT 932.100 237.000 933.900 243.600 ;
        RECT 935.100 237.600 936.900 243.600 ;
        RECT 938.100 237.000 939.900 243.600 ;
        RECT 956.100 237.600 957.900 243.600 ;
        RECT 962.100 243.600 963.600 243.900 ;
        RECT 959.100 237.000 960.900 243.000 ;
        RECT 962.100 237.600 963.900 243.600 ;
        RECT 965.100 237.000 966.900 243.600 ;
        RECT 983.100 237.600 984.900 249.600 ;
        RECT 986.100 237.000 987.900 249.600 ;
        RECT 1007.100 248.100 1009.500 249.600 ;
        RECT 1005.000 245.100 1006.800 246.900 ;
        RECT 1004.700 237.000 1006.500 243.600 ;
        RECT 1007.700 237.600 1009.500 248.100 ;
        RECT 1012.800 237.000 1014.600 249.600 ;
        RECT 1034.100 248.100 1036.500 249.600 ;
        RECT 1032.000 245.100 1033.800 246.900 ;
        RECT 1031.700 237.000 1033.500 243.600 ;
        RECT 1034.700 237.600 1036.500 248.100 ;
        RECT 1039.800 237.000 1041.600 249.600 ;
        RECT 17.100 227.400 18.900 234.000 ;
        RECT 20.100 227.400 21.900 233.400 ;
        RECT 23.100 227.400 24.900 234.000 ;
        RECT 41.100 227.400 42.900 234.000 ;
        RECT 44.100 227.400 45.900 233.400 ;
        RECT 47.100 227.400 48.900 234.000 ;
        RECT 65.100 227.400 66.900 233.400 ;
        RECT 68.100 227.400 69.900 234.000 ;
        RECT 86.700 227.400 88.500 234.000 ;
        RECT 20.100 214.050 21.300 227.400 ;
        RECT 44.700 214.050 45.900 227.400 ;
        RECT 65.700 214.050 66.900 227.400 ;
        RECT 87.000 224.100 88.800 225.900 ;
        RECT 89.700 222.900 91.500 233.400 ;
        RECT 89.100 221.400 91.500 222.900 ;
        RECT 94.800 221.400 96.600 234.000 ;
        RECT 113.100 227.400 114.900 234.000 ;
        RECT 116.100 227.400 117.900 233.400 ;
        RECT 119.100 227.400 120.900 234.000 ;
        RECT 137.100 227.400 138.900 233.400 ;
        RECT 140.100 228.000 141.900 234.000 ;
        RECT 76.950 219.450 79.050 220.050 ;
        RECT 85.950 219.450 88.050 220.200 ;
        RECT 76.950 218.550 88.050 219.450 ;
        RECT 76.950 217.950 79.050 218.550 ;
        RECT 85.950 218.100 88.050 218.550 ;
        RECT 68.100 214.050 69.900 215.850 ;
        RECT 89.100 214.050 90.300 221.400 ;
        RECT 95.100 214.050 96.900 215.850 ;
        RECT 116.700 214.050 117.900 227.400 ;
        RECT 138.000 227.100 138.900 227.400 ;
        RECT 143.100 227.400 144.900 233.400 ;
        RECT 146.100 227.400 147.900 234.000 ;
        RECT 143.100 227.100 144.600 227.400 ;
        RECT 138.000 226.200 144.600 227.100 ;
        RECT 121.950 216.450 126.000 217.050 ;
        RECT 121.950 214.950 126.450 216.450 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 19.950 211.950 22.050 214.050 ;
        RECT 22.950 211.950 25.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 46.950 211.950 49.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 17.250 210.150 19.050 211.950 ;
        RECT 20.100 206.700 21.300 211.950 ;
        RECT 23.100 210.150 24.900 211.950 ;
        RECT 41.100 210.150 42.900 211.950 ;
        RECT 44.700 206.700 45.900 211.950 ;
        RECT 46.950 210.150 48.750 211.950 ;
        RECT 20.100 205.800 24.300 206.700 ;
        RECT 17.400 198.000 19.200 204.600 ;
        RECT 22.500 198.600 24.300 205.800 ;
        RECT 41.700 205.800 45.900 206.700 ;
        RECT 46.950 207.450 49.050 208.050 ;
        RECT 52.950 207.450 55.050 208.050 ;
        RECT 46.950 206.550 55.050 207.450 ;
        RECT 46.950 205.950 49.050 206.550 ;
        RECT 52.950 205.950 55.050 206.550 ;
        RECT 41.700 198.600 43.500 205.800 ;
        RECT 46.800 198.000 48.600 204.600 ;
        RECT 65.700 201.600 66.900 211.950 ;
        RECT 86.100 210.150 87.900 211.950 ;
        RECT 89.100 207.600 90.300 211.950 ;
        RECT 92.100 210.150 93.900 211.950 ;
        RECT 113.100 210.150 114.900 211.950 ;
        RECT 86.700 206.700 90.300 207.600 ;
        RECT 116.700 206.700 117.900 211.950 ;
        RECT 118.950 210.150 120.750 211.950 ;
        RECT 125.550 211.050 126.450 214.950 ;
        RECT 138.000 214.050 138.900 226.200 ;
        RECT 139.950 222.450 142.050 223.050 ;
        RECT 154.950 222.450 157.050 223.050 ;
        RECT 139.950 221.550 157.050 222.450 ;
        RECT 139.950 220.950 142.050 221.550 ;
        RECT 154.950 220.950 157.050 221.550 ;
        RECT 165.000 222.600 166.800 233.400 ;
        RECT 165.000 221.400 168.600 222.600 ;
        RECT 170.100 221.400 171.900 234.000 ;
        RECT 188.100 227.400 189.900 234.000 ;
        RECT 191.100 227.400 192.900 233.400 ;
        RECT 194.100 227.400 195.900 234.000 ;
        RECT 143.100 214.050 144.900 215.850 ;
        RECT 164.100 214.050 165.900 215.850 ;
        RECT 167.700 214.050 168.600 221.400 ;
        RECT 169.950 214.050 171.750 215.850 ;
        RECT 191.700 214.050 192.900 227.400 ;
        RECT 212.100 221.400 213.900 233.400 ;
        RECT 215.100 222.000 216.900 234.000 ;
        RECT 218.100 227.400 219.900 233.400 ;
        RECT 221.100 227.400 222.900 234.000 ;
        RECT 239.100 227.400 240.900 234.000 ;
        RECT 242.100 227.400 243.900 233.400 ;
        RECT 245.100 227.400 246.900 234.000 ;
        RECT 263.100 227.400 264.900 233.400 ;
        RECT 266.100 228.000 267.900 234.000 ;
        RECT 212.700 214.050 213.600 221.400 ;
        RECT 216.000 214.050 217.800 215.850 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 145.950 211.950 148.050 214.050 ;
        RECT 163.950 211.950 166.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 212.100 211.950 214.200 214.050 ;
        RECT 215.400 211.950 217.500 214.050 ;
        RECT 121.950 209.550 126.450 211.050 ;
        RECT 121.950 208.950 126.000 209.550 ;
        RECT 138.000 208.200 138.900 211.950 ;
        RECT 140.100 210.150 141.900 211.950 ;
        RECT 146.100 210.150 147.900 211.950 ;
        RECT 138.000 207.000 141.300 208.200 ;
        RECT 86.700 204.600 87.900 206.700 ;
        RECT 113.700 205.800 117.900 206.700 ;
        RECT 65.100 198.600 66.900 201.600 ;
        RECT 68.100 198.000 69.900 201.600 ;
        RECT 86.100 198.600 87.900 204.600 ;
        RECT 89.100 203.700 96.900 205.050 ;
        RECT 89.100 198.600 90.900 203.700 ;
        RECT 92.100 198.000 93.900 202.800 ;
        RECT 95.100 198.600 96.900 203.700 ;
        RECT 113.700 198.600 115.500 205.800 ;
        RECT 118.800 198.000 120.600 204.600 ;
        RECT 139.500 198.600 141.300 207.000 ;
        RECT 146.100 198.000 147.900 207.600 ;
        RECT 167.700 201.600 168.600 211.950 ;
        RECT 188.100 210.150 189.900 211.950 ;
        RECT 191.700 206.700 192.900 211.950 ;
        RECT 193.950 210.150 195.750 211.950 ;
        RECT 188.700 205.800 192.900 206.700 ;
        RECT 164.100 198.000 165.900 201.600 ;
        RECT 167.100 198.600 168.900 201.600 ;
        RECT 170.100 198.000 171.900 201.600 ;
        RECT 188.700 198.600 190.500 205.800 ;
        RECT 212.700 204.600 213.600 211.950 ;
        RECT 219.000 207.300 219.900 227.400 ;
        RECT 242.100 214.050 243.300 227.400 ;
        RECT 264.000 227.100 264.900 227.400 ;
        RECT 269.100 227.400 270.900 233.400 ;
        RECT 272.100 227.400 273.900 234.000 ;
        RECT 290.700 227.400 292.500 234.000 ;
        RECT 269.100 227.100 270.600 227.400 ;
        RECT 264.000 226.200 270.600 227.100 ;
        RECT 264.000 214.050 264.900 226.200 ;
        RECT 291.000 224.100 292.800 225.900 ;
        RECT 293.700 222.900 295.500 233.400 ;
        RECT 293.100 221.400 295.500 222.900 ;
        RECT 298.800 221.400 300.600 234.000 ;
        RECT 317.100 227.400 318.900 234.000 ;
        RECT 320.100 227.400 321.900 233.400 ;
        RECT 323.100 227.400 324.900 234.000 ;
        RECT 341.100 227.400 342.900 234.000 ;
        RECT 344.100 227.400 345.900 233.400 ;
        RECT 347.100 227.400 348.900 234.000 ;
        RECT 365.100 227.400 366.900 234.000 ;
        RECT 368.100 227.400 369.900 233.400 ;
        RECT 371.100 227.400 372.900 234.000 ;
        RECT 374.700 227.400 376.500 234.000 ;
        RECT 377.700 227.400 379.500 233.400 ;
        RECT 381.000 227.400 382.800 234.000 ;
        RECT 384.000 227.400 385.800 233.400 ;
        RECT 387.000 227.400 388.800 234.000 ;
        RECT 390.000 227.400 391.800 233.400 ;
        RECT 393.000 227.400 394.800 234.000 ;
        RECT 396.000 230.400 397.800 233.400 ;
        RECT 399.000 230.400 400.800 233.400 ;
        RECT 402.000 230.400 403.800 233.400 ;
        RECT 395.700 228.300 397.800 230.400 ;
        RECT 398.700 228.300 400.800 230.400 ;
        RECT 401.700 228.300 403.800 230.400 ;
        RECT 405.000 227.400 406.800 233.400 ;
        RECT 408.000 227.400 409.800 234.000 ;
        RECT 269.100 214.050 270.900 215.850 ;
        RECT 293.100 214.050 294.300 221.400 ;
        RECT 299.100 214.050 300.900 215.850 ;
        RECT 320.100 214.050 321.300 227.400 ;
        RECT 344.100 214.050 345.300 227.400 ;
        RECT 349.950 216.450 354.000 217.050 ;
        RECT 349.950 214.950 354.450 216.450 ;
        RECT 220.800 211.950 222.900 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 346.950 211.950 349.050 214.050 ;
        RECT 220.950 210.150 222.750 211.950 ;
        RECT 239.250 210.150 241.050 211.950 ;
        RECT 214.500 206.400 222.900 207.300 ;
        RECT 214.500 205.500 216.300 206.400 ;
        RECT 193.800 198.000 195.600 204.600 ;
        RECT 212.700 202.800 215.400 204.600 ;
        RECT 213.600 198.600 215.400 202.800 ;
        RECT 216.600 198.000 218.400 204.600 ;
        RECT 221.100 198.600 222.900 206.400 ;
        RECT 242.100 206.700 243.300 211.950 ;
        RECT 245.100 210.150 246.900 211.950 ;
        RECT 264.000 208.200 264.900 211.950 ;
        RECT 266.100 210.150 267.900 211.950 ;
        RECT 272.100 210.150 273.900 211.950 ;
        RECT 290.100 210.150 291.900 211.950 ;
        RECT 264.000 207.000 267.300 208.200 ;
        RECT 293.100 207.600 294.300 211.950 ;
        RECT 296.100 210.150 297.900 211.950 ;
        RECT 317.250 210.150 319.050 211.950 ;
        RECT 242.100 205.800 246.300 206.700 ;
        RECT 239.400 198.000 241.200 204.600 ;
        RECT 244.500 198.600 246.300 205.800 ;
        RECT 265.500 198.600 267.300 207.000 ;
        RECT 272.100 198.000 273.900 207.600 ;
        RECT 290.700 206.700 294.300 207.600 ;
        RECT 320.100 206.700 321.300 211.950 ;
        RECT 323.100 210.150 324.900 211.950 ;
        RECT 341.250 210.150 343.050 211.950 ;
        RECT 344.100 206.700 345.300 211.950 ;
        RECT 347.100 210.150 348.900 211.950 ;
        RECT 353.550 210.450 354.450 214.950 ;
        RECT 368.700 214.050 369.900 227.400 ;
        RECT 378.000 217.050 379.500 227.400 ;
        RECT 384.000 226.500 385.200 227.400 ;
        RECT 377.100 214.950 379.500 217.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 361.950 210.450 364.050 211.050 ;
        RECT 353.550 209.550 364.050 210.450 ;
        RECT 365.100 210.150 366.900 211.950 ;
        RECT 361.950 208.950 364.050 209.550 ;
        RECT 368.700 206.700 369.900 211.950 ;
        RECT 370.950 210.150 372.750 211.950 ;
        RECT 290.700 204.600 291.900 206.700 ;
        RECT 320.100 205.800 324.300 206.700 ;
        RECT 344.100 205.800 348.300 206.700 ;
        RECT 290.100 198.600 291.900 204.600 ;
        RECT 293.100 203.700 300.900 205.050 ;
        RECT 293.100 198.600 294.900 203.700 ;
        RECT 296.100 198.000 297.900 202.800 ;
        RECT 299.100 198.600 300.900 203.700 ;
        RECT 317.400 198.000 319.200 204.600 ;
        RECT 322.500 198.600 324.300 205.800 ;
        RECT 341.400 198.000 343.200 204.600 ;
        RECT 346.500 198.600 348.300 205.800 ;
        RECT 365.700 205.800 369.900 206.700 ;
        RECT 365.700 198.600 367.500 205.800 ;
        RECT 370.800 198.000 372.600 204.600 ;
        RECT 378.000 201.600 379.500 214.950 ;
        RECT 374.700 198.000 376.500 201.600 ;
        RECT 377.700 198.600 379.500 201.600 ;
        RECT 381.300 225.600 385.200 226.500 ;
        RECT 381.300 222.300 382.200 225.600 ;
        RECT 386.100 224.400 387.900 225.000 ;
        RECT 390.600 224.400 391.800 227.400 ;
        RECT 398.700 226.500 400.800 227.400 ;
        RECT 392.700 225.300 400.800 226.500 ;
        RECT 392.700 224.700 394.500 225.300 ;
        RECT 386.100 223.200 391.800 224.400 ;
        RECT 404.100 223.500 406.800 227.400 ;
        RECT 411.000 225.900 412.800 233.400 ;
        RECT 414.900 227.400 416.700 234.000 ;
        RECT 417.900 227.400 419.700 233.400 ;
        RECT 420.900 230.400 422.700 233.400 ;
        RECT 423.900 230.400 425.700 233.400 ;
        RECT 420.600 228.300 422.700 230.400 ;
        RECT 423.600 228.300 425.700 230.400 ;
        RECT 427.500 227.400 429.300 234.000 ;
        RECT 409.500 223.800 412.800 225.900 ;
        RECT 418.200 225.300 420.300 227.400 ;
        RECT 430.500 224.400 432.300 233.400 ;
        RECT 433.500 227.400 435.300 234.000 ;
        RECT 436.500 228.300 438.300 233.400 ;
        RECT 436.500 227.400 438.600 228.300 ;
        RECT 439.500 227.400 441.300 234.000 ;
        RECT 437.700 226.500 438.600 227.400 ;
        RECT 437.700 225.600 441.300 226.500 ;
        RECT 435.000 224.400 436.800 224.700 ;
        RECT 395.700 222.300 397.800 223.500 ;
        RECT 381.300 221.400 397.800 222.300 ;
        RECT 401.100 222.600 403.200 223.500 ;
        RECT 417.600 223.200 436.800 224.400 ;
        RECT 417.600 222.600 418.800 223.200 ;
        RECT 435.000 222.900 436.800 223.200 ;
        RECT 401.100 221.400 418.800 222.600 ;
        RECT 421.500 221.700 423.600 222.300 ;
        RECT 431.700 221.700 433.500 222.300 ;
        RECT 381.300 204.600 382.200 221.400 ;
        RECT 421.500 220.500 433.500 221.700 ;
        RECT 383.100 219.300 418.800 220.500 ;
        RECT 421.500 220.200 423.600 220.500 ;
        RECT 383.100 218.700 384.900 219.300 ;
        RECT 417.600 218.700 418.800 219.300 ;
        RECT 386.100 214.950 388.200 217.050 ;
        RECT 386.700 212.100 388.200 214.950 ;
        RECT 390.300 214.800 395.400 216.600 ;
        RECT 394.500 213.300 395.400 214.800 ;
        RECT 398.100 216.300 399.900 218.100 ;
        RECT 404.100 217.800 406.200 218.100 ;
        RECT 417.600 217.800 431.100 218.700 ;
        RECT 398.100 215.100 399.000 216.300 ;
        RECT 404.100 216.000 408.000 217.800 ;
        RECT 409.500 216.300 411.600 217.200 ;
        RECT 429.300 217.050 431.100 217.800 ;
        RECT 409.500 215.100 420.600 216.300 ;
        RECT 429.300 215.250 433.200 217.050 ;
        RECT 398.100 214.200 411.600 215.100 ;
        RECT 418.800 214.500 420.600 215.100 ;
        RECT 431.100 214.950 433.200 215.250 ;
        RECT 437.100 214.950 439.200 217.050 ;
        RECT 437.100 213.300 438.900 214.950 ;
        RECT 394.500 212.100 438.900 213.300 ;
        RECT 386.700 210.600 393.300 212.100 ;
        RECT 383.100 207.900 390.900 209.700 ;
        RECT 391.800 209.100 408.900 210.600 ;
        RECT 406.800 208.500 408.900 209.100 ;
        RECT 413.100 210.000 415.200 211.050 ;
        RECT 413.100 209.100 418.200 210.000 ;
        RECT 421.800 209.400 423.600 211.200 ;
        RECT 440.100 209.400 441.300 225.600 ;
        RECT 458.400 221.400 460.200 234.000 ;
        RECT 463.500 222.900 465.300 233.400 ;
        RECT 466.500 227.400 468.300 234.000 ;
        RECT 466.200 224.100 468.000 225.900 ;
        RECT 463.500 221.400 465.900 222.900 ;
        RECT 485.400 221.400 487.200 234.000 ;
        RECT 490.500 222.900 492.300 233.400 ;
        RECT 493.500 227.400 495.300 234.000 ;
        RECT 512.100 227.400 513.900 233.400 ;
        RECT 493.200 224.100 495.000 225.900 ;
        RECT 490.500 221.400 492.900 222.900 ;
        RECT 458.100 214.050 459.900 215.850 ;
        RECT 464.700 214.050 465.900 221.400 ;
        RECT 485.100 214.050 486.900 215.850 ;
        RECT 491.700 214.050 492.900 221.400 ;
        RECT 512.100 220.500 513.300 227.400 ;
        RECT 515.100 223.200 516.900 234.000 ;
        RECT 518.100 221.400 519.900 233.400 ;
        RECT 521.700 227.400 523.500 234.000 ;
        RECT 524.700 228.300 526.500 233.400 ;
        RECT 524.400 227.400 526.500 228.300 ;
        RECT 527.700 227.400 529.500 234.000 ;
        RECT 524.400 226.500 525.300 227.400 ;
        RECT 512.100 219.600 517.800 220.500 ;
        RECT 516.000 218.700 517.800 219.600 ;
        RECT 512.400 214.050 514.200 215.850 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 512.400 211.950 514.500 214.050 ;
        RECT 461.100 210.150 462.900 211.950 ;
        RECT 413.100 208.950 415.200 209.100 ;
        RECT 389.400 204.600 390.900 207.900 ;
        RECT 407.100 206.700 408.900 208.500 ;
        RECT 416.400 208.200 418.200 209.100 ;
        RECT 422.700 206.400 423.600 209.400 ;
        RECT 424.500 208.200 441.300 209.400 ;
        RECT 424.500 207.300 426.600 208.200 ;
        RECT 435.300 206.700 437.100 207.300 ;
        RECT 395.100 204.600 401.700 206.400 ;
        RECT 416.400 205.200 423.600 206.400 ;
        RECT 428.700 205.500 437.100 206.700 ;
        RECT 416.400 204.600 417.300 205.200 ;
        RECT 419.400 204.600 421.200 205.200 ;
        RECT 428.700 204.600 430.200 205.500 ;
        RECT 440.100 204.600 441.300 208.200 ;
        RECT 464.700 207.600 465.900 211.950 ;
        RECT 467.100 210.150 468.900 211.950 ;
        RECT 488.100 210.150 489.900 211.950 ;
        RECT 491.700 207.600 492.900 211.950 ;
        RECT 494.100 210.150 495.900 211.950 ;
        RECT 464.700 206.700 468.300 207.600 ;
        RECT 491.700 206.700 495.300 207.600 ;
        RECT 381.300 198.600 383.100 204.600 ;
        RECT 386.700 198.000 388.500 204.600 ;
        RECT 389.400 203.400 393.600 204.600 ;
        RECT 391.800 198.600 393.600 203.400 ;
        RECT 395.700 201.600 397.800 203.700 ;
        RECT 398.700 201.600 400.800 203.700 ;
        RECT 401.700 201.600 403.800 203.700 ;
        RECT 404.700 201.600 406.800 203.700 ;
        RECT 410.100 202.500 412.800 204.600 ;
        RECT 414.600 203.400 417.300 204.600 ;
        RECT 414.600 202.500 416.400 203.400 ;
        RECT 396.000 198.600 397.800 201.600 ;
        RECT 399.000 198.600 400.800 201.600 ;
        RECT 402.000 198.600 403.800 201.600 ;
        RECT 405.000 198.600 406.800 201.600 ;
        RECT 408.000 198.000 409.800 201.600 ;
        RECT 411.000 198.600 412.800 202.500 ;
        RECT 418.200 201.600 420.300 203.700 ;
        RECT 421.200 201.600 423.300 203.700 ;
        RECT 424.200 201.600 426.300 203.700 ;
        RECT 415.500 198.000 417.300 201.600 ;
        RECT 418.500 198.600 420.300 201.600 ;
        RECT 421.500 198.600 423.300 201.600 ;
        RECT 424.500 198.600 426.300 201.600 ;
        RECT 428.700 198.600 430.500 204.600 ;
        RECT 434.100 198.000 435.900 204.600 ;
        RECT 439.500 198.600 441.300 204.600 ;
        RECT 458.100 203.700 465.900 205.050 ;
        RECT 458.100 198.600 459.900 203.700 ;
        RECT 461.100 198.000 462.900 202.800 ;
        RECT 464.100 198.600 465.900 203.700 ;
        RECT 467.100 204.600 468.300 206.700 ;
        RECT 467.100 198.600 468.900 204.600 ;
        RECT 485.100 203.700 492.900 205.050 ;
        RECT 485.100 198.600 486.900 203.700 ;
        RECT 488.100 198.000 489.900 202.800 ;
        RECT 491.100 198.600 492.900 203.700 ;
        RECT 494.100 204.600 495.300 206.700 ;
        RECT 516.000 207.300 516.900 218.700 ;
        RECT 518.700 214.050 519.900 221.400 ;
        RECT 517.800 211.950 519.900 214.050 ;
        RECT 516.000 206.400 517.800 207.300 ;
        RECT 512.100 205.500 517.800 206.400 ;
        RECT 494.100 198.600 495.900 204.600 ;
        RECT 512.100 201.600 513.300 205.500 ;
        RECT 518.700 204.600 519.900 211.950 ;
        RECT 512.100 198.600 513.900 201.600 ;
        RECT 515.100 198.000 516.900 204.600 ;
        RECT 518.100 198.600 519.900 204.600 ;
        RECT 521.700 225.600 525.300 226.500 ;
        RECT 521.700 209.400 522.900 225.600 ;
        RECT 526.200 224.400 528.000 224.700 ;
        RECT 530.700 224.400 532.500 233.400 ;
        RECT 533.700 227.400 535.500 234.000 ;
        RECT 537.300 230.400 539.100 233.400 ;
        RECT 540.300 230.400 542.100 233.400 ;
        RECT 537.300 228.300 539.400 230.400 ;
        RECT 540.300 228.300 542.400 230.400 ;
        RECT 543.300 227.400 545.100 233.400 ;
        RECT 546.300 227.400 548.100 234.000 ;
        RECT 542.700 225.300 544.800 227.400 ;
        RECT 550.200 225.900 552.000 233.400 ;
        RECT 553.200 227.400 555.000 234.000 ;
        RECT 556.200 227.400 558.000 233.400 ;
        RECT 559.200 230.400 561.000 233.400 ;
        RECT 562.200 230.400 564.000 233.400 ;
        RECT 565.200 230.400 567.000 233.400 ;
        RECT 559.200 228.300 561.300 230.400 ;
        RECT 562.200 228.300 564.300 230.400 ;
        RECT 565.200 228.300 567.300 230.400 ;
        RECT 568.200 227.400 570.000 234.000 ;
        RECT 571.200 227.400 573.000 233.400 ;
        RECT 574.200 227.400 576.000 234.000 ;
        RECT 577.200 227.400 579.000 233.400 ;
        RECT 580.200 227.400 582.000 234.000 ;
        RECT 583.500 227.400 585.300 233.400 ;
        RECT 586.500 227.400 588.300 234.000 ;
        RECT 526.200 223.200 545.400 224.400 ;
        RECT 550.200 223.800 553.500 225.900 ;
        RECT 556.200 223.500 558.900 227.400 ;
        RECT 562.200 226.500 564.300 227.400 ;
        RECT 562.200 225.300 570.300 226.500 ;
        RECT 568.500 224.700 570.300 225.300 ;
        RECT 571.200 224.400 572.400 227.400 ;
        RECT 577.800 226.500 579.000 227.400 ;
        RECT 577.800 225.600 581.700 226.500 ;
        RECT 575.100 224.400 576.900 225.000 ;
        RECT 526.200 222.900 528.000 223.200 ;
        RECT 544.200 222.600 545.400 223.200 ;
        RECT 559.800 222.600 561.900 223.500 ;
        RECT 529.500 221.700 531.300 222.300 ;
        RECT 539.400 221.700 541.500 222.300 ;
        RECT 529.500 220.500 541.500 221.700 ;
        RECT 544.200 221.400 561.900 222.600 ;
        RECT 565.200 222.300 567.300 223.500 ;
        RECT 571.200 223.200 576.900 224.400 ;
        RECT 580.800 222.300 581.700 225.600 ;
        RECT 565.200 221.400 581.700 222.300 ;
        RECT 539.400 220.200 541.500 220.500 ;
        RECT 544.200 219.300 579.900 220.500 ;
        RECT 544.200 218.700 545.400 219.300 ;
        RECT 578.100 218.700 579.900 219.300 ;
        RECT 531.900 217.800 545.400 218.700 ;
        RECT 556.800 217.800 558.900 218.100 ;
        RECT 531.900 217.050 533.700 217.800 ;
        RECT 523.800 214.950 525.900 217.050 ;
        RECT 529.800 215.250 533.700 217.050 ;
        RECT 551.400 216.300 553.500 217.200 ;
        RECT 529.800 214.950 531.900 215.250 ;
        RECT 542.400 215.100 553.500 216.300 ;
        RECT 555.000 216.000 558.900 217.800 ;
        RECT 563.100 216.300 564.900 218.100 ;
        RECT 564.000 215.100 564.900 216.300 ;
        RECT 524.100 213.300 525.900 214.950 ;
        RECT 542.400 214.500 544.200 215.100 ;
        RECT 551.400 214.200 564.900 215.100 ;
        RECT 567.600 214.800 572.700 216.600 ;
        RECT 574.800 214.950 576.900 217.050 ;
        RECT 567.600 213.300 568.500 214.800 ;
        RECT 524.100 212.100 568.500 213.300 ;
        RECT 574.800 212.100 576.300 214.950 ;
        RECT 539.400 209.400 541.200 211.200 ;
        RECT 547.800 210.000 549.900 211.050 ;
        RECT 569.700 210.600 576.300 212.100 ;
        RECT 521.700 208.200 538.500 209.400 ;
        RECT 521.700 204.600 522.900 208.200 ;
        RECT 536.400 207.300 538.500 208.200 ;
        RECT 525.900 206.700 527.700 207.300 ;
        RECT 525.900 205.500 534.300 206.700 ;
        RECT 532.800 204.600 534.300 205.500 ;
        RECT 539.400 206.400 540.300 209.400 ;
        RECT 544.800 209.100 549.900 210.000 ;
        RECT 544.800 208.200 546.600 209.100 ;
        RECT 547.800 208.950 549.900 209.100 ;
        RECT 554.100 209.100 571.200 210.600 ;
        RECT 554.100 208.500 556.200 209.100 ;
        RECT 554.100 206.700 555.900 208.500 ;
        RECT 572.100 207.900 579.900 209.700 ;
        RECT 539.400 205.200 546.600 206.400 ;
        RECT 541.800 204.600 543.600 205.200 ;
        RECT 545.700 204.600 546.600 205.200 ;
        RECT 561.300 204.600 567.900 206.400 ;
        RECT 572.100 204.600 573.600 207.900 ;
        RECT 580.800 204.600 581.700 221.400 ;
        RECT 521.700 198.600 523.500 204.600 ;
        RECT 527.100 198.000 528.900 204.600 ;
        RECT 532.500 198.600 534.300 204.600 ;
        RECT 536.700 201.600 538.800 203.700 ;
        RECT 539.700 201.600 541.800 203.700 ;
        RECT 542.700 201.600 544.800 203.700 ;
        RECT 545.700 203.400 548.400 204.600 ;
        RECT 546.600 202.500 548.400 203.400 ;
        RECT 550.200 202.500 552.900 204.600 ;
        RECT 536.700 198.600 538.500 201.600 ;
        RECT 539.700 198.600 541.500 201.600 ;
        RECT 542.700 198.600 544.500 201.600 ;
        RECT 545.700 198.000 547.500 201.600 ;
        RECT 550.200 198.600 552.000 202.500 ;
        RECT 556.200 201.600 558.300 203.700 ;
        RECT 559.200 201.600 561.300 203.700 ;
        RECT 562.200 201.600 564.300 203.700 ;
        RECT 565.200 201.600 567.300 203.700 ;
        RECT 569.400 203.400 573.600 204.600 ;
        RECT 553.200 198.000 555.000 201.600 ;
        RECT 556.200 198.600 558.000 201.600 ;
        RECT 559.200 198.600 561.000 201.600 ;
        RECT 562.200 198.600 564.000 201.600 ;
        RECT 565.200 198.600 567.000 201.600 ;
        RECT 569.400 198.600 571.200 203.400 ;
        RECT 574.500 198.000 576.300 204.600 ;
        RECT 579.900 198.600 581.700 204.600 ;
        RECT 583.500 217.050 585.000 227.400 ;
        RECT 606.000 222.600 607.800 233.400 ;
        RECT 606.000 221.400 609.600 222.600 ;
        RECT 611.100 221.400 612.900 234.000 ;
        RECT 629.700 227.400 631.500 234.000 ;
        RECT 630.000 224.100 631.800 225.900 ;
        RECT 632.700 222.900 634.500 233.400 ;
        RECT 632.100 221.400 634.500 222.900 ;
        RECT 637.800 221.400 639.600 234.000 ;
        RECT 656.100 227.400 657.900 234.000 ;
        RECT 659.100 227.400 660.900 233.400 ;
        RECT 662.100 227.400 663.900 234.000 ;
        RECT 583.500 214.950 585.900 217.050 ;
        RECT 583.500 201.600 585.000 214.950 ;
        RECT 605.100 214.050 606.900 215.850 ;
        RECT 608.700 214.050 609.600 221.400 ;
        RECT 610.950 214.050 612.750 215.850 ;
        RECT 632.100 214.050 633.300 221.400 ;
        RECT 638.100 214.050 639.900 215.850 ;
        RECT 659.100 214.050 660.300 227.400 ;
        RECT 680.100 222.600 681.900 233.400 ;
        RECT 683.100 223.500 684.900 234.000 ;
        RECT 686.100 232.500 693.900 233.400 ;
        RECT 686.100 222.600 687.900 232.500 ;
        RECT 680.100 221.700 687.900 222.600 ;
        RECT 689.100 220.500 690.900 231.600 ;
        RECT 692.100 221.400 693.900 232.500 ;
        RECT 710.100 227.400 711.900 233.400 ;
        RECT 713.100 228.000 714.900 234.000 ;
        RECT 711.000 227.100 711.900 227.400 ;
        RECT 716.100 227.400 717.900 233.400 ;
        RECT 719.100 227.400 720.900 234.000 ;
        RECT 737.100 227.400 738.900 233.400 ;
        RECT 740.100 227.400 741.900 234.000 ;
        RECT 716.100 227.100 717.600 227.400 ;
        RECT 711.000 226.200 717.600 227.100 ;
        RECT 686.100 219.600 690.900 220.500 ;
        RECT 683.250 214.050 685.050 215.850 ;
        RECT 686.100 214.050 687.000 219.600 ;
        RECT 689.100 214.050 690.900 215.850 ;
        RECT 711.000 214.050 711.900 226.200 ;
        RECT 716.100 214.050 717.900 215.850 ;
        RECT 737.700 214.050 738.900 227.400 ;
        RECT 758.100 221.400 759.900 233.400 ;
        RECT 761.100 222.300 762.900 233.400 ;
        RECT 764.100 223.200 765.900 234.000 ;
        RECT 767.100 222.300 768.900 233.400 ;
        RECT 770.700 227.400 772.500 234.000 ;
        RECT 773.700 227.400 775.500 233.400 ;
        RECT 777.000 227.400 778.800 234.000 ;
        RECT 780.000 227.400 781.800 233.400 ;
        RECT 783.000 227.400 784.800 234.000 ;
        RECT 786.000 227.400 787.800 233.400 ;
        RECT 789.000 227.400 790.800 234.000 ;
        RECT 792.000 230.400 793.800 233.400 ;
        RECT 795.000 230.400 796.800 233.400 ;
        RECT 798.000 230.400 799.800 233.400 ;
        RECT 791.700 228.300 793.800 230.400 ;
        RECT 794.700 228.300 796.800 230.400 ;
        RECT 797.700 228.300 799.800 230.400 ;
        RECT 801.000 227.400 802.800 233.400 ;
        RECT 804.000 227.400 805.800 234.000 ;
        RECT 761.100 221.400 768.900 222.300 ;
        RECT 740.100 214.050 741.900 215.850 ;
        RECT 758.400 214.050 759.300 221.400 ;
        RECT 774.000 217.050 775.500 227.400 ;
        RECT 780.000 226.500 781.200 227.400 ;
        RECT 763.950 214.050 765.750 215.850 ;
        RECT 773.100 214.950 775.500 217.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 608.700 201.600 609.600 211.950 ;
        RECT 629.100 210.150 630.900 211.950 ;
        RECT 632.100 207.600 633.300 211.950 ;
        RECT 635.100 210.150 636.900 211.950 ;
        RECT 656.250 210.150 658.050 211.950 ;
        RECT 629.700 206.700 633.300 207.600 ;
        RECT 659.100 206.700 660.300 211.950 ;
        RECT 662.100 210.150 663.900 211.950 ;
        RECT 680.250 210.150 682.050 211.950 ;
        RECT 629.700 204.600 630.900 206.700 ;
        RECT 659.100 205.800 663.300 206.700 ;
        RECT 583.500 198.600 585.300 201.600 ;
        RECT 586.500 198.000 588.300 201.600 ;
        RECT 605.100 198.000 606.900 201.600 ;
        RECT 608.100 198.600 609.900 201.600 ;
        RECT 611.100 198.000 612.900 201.600 ;
        RECT 629.100 198.600 630.900 204.600 ;
        RECT 632.100 203.700 639.900 205.050 ;
        RECT 632.100 198.600 633.900 203.700 ;
        RECT 635.100 198.000 636.900 202.800 ;
        RECT 638.100 198.600 639.900 203.700 ;
        RECT 656.400 198.000 658.200 204.600 ;
        RECT 661.500 198.600 663.300 205.800 ;
        RECT 686.100 204.600 687.300 211.950 ;
        RECT 692.100 210.150 693.900 211.950 ;
        RECT 711.000 208.200 711.900 211.950 ;
        RECT 713.100 210.150 714.900 211.950 ;
        RECT 719.100 210.150 720.900 211.950 ;
        RECT 711.000 207.000 714.300 208.200 ;
        RECT 680.700 198.000 682.500 204.600 ;
        RECT 685.200 198.600 687.000 204.600 ;
        RECT 689.700 198.000 691.500 204.600 ;
        RECT 712.500 198.600 714.300 207.000 ;
        RECT 719.100 198.000 720.900 207.600 ;
        RECT 737.700 201.600 738.900 211.950 ;
        RECT 758.400 204.600 759.300 211.950 ;
        RECT 760.950 210.150 762.750 211.950 ;
        RECT 767.100 210.150 768.900 211.950 ;
        RECT 758.400 203.400 763.500 204.600 ;
        RECT 737.100 198.600 738.900 201.600 ;
        RECT 740.100 198.000 741.900 201.600 ;
        RECT 758.700 198.000 760.500 201.600 ;
        RECT 761.700 198.600 763.500 203.400 ;
        RECT 766.200 198.000 768.000 204.600 ;
        RECT 774.000 201.600 775.500 214.950 ;
        RECT 770.700 198.000 772.500 201.600 ;
        RECT 773.700 198.600 775.500 201.600 ;
        RECT 777.300 225.600 781.200 226.500 ;
        RECT 777.300 222.300 778.200 225.600 ;
        RECT 782.100 224.400 783.900 225.000 ;
        RECT 786.600 224.400 787.800 227.400 ;
        RECT 794.700 226.500 796.800 227.400 ;
        RECT 788.700 225.300 796.800 226.500 ;
        RECT 788.700 224.700 790.500 225.300 ;
        RECT 782.100 223.200 787.800 224.400 ;
        RECT 800.100 223.500 802.800 227.400 ;
        RECT 807.000 225.900 808.800 233.400 ;
        RECT 810.900 227.400 812.700 234.000 ;
        RECT 813.900 227.400 815.700 233.400 ;
        RECT 816.900 230.400 818.700 233.400 ;
        RECT 819.900 230.400 821.700 233.400 ;
        RECT 816.600 228.300 818.700 230.400 ;
        RECT 819.600 228.300 821.700 230.400 ;
        RECT 823.500 227.400 825.300 234.000 ;
        RECT 805.500 223.800 808.800 225.900 ;
        RECT 814.200 225.300 816.300 227.400 ;
        RECT 826.500 224.400 828.300 233.400 ;
        RECT 829.500 227.400 831.300 234.000 ;
        RECT 832.500 228.300 834.300 233.400 ;
        RECT 832.500 227.400 834.600 228.300 ;
        RECT 835.500 227.400 837.300 234.000 ;
        RECT 854.100 227.400 855.900 234.000 ;
        RECT 857.100 227.400 858.900 233.400 ;
        RECT 860.700 227.400 862.500 234.000 ;
        RECT 863.700 228.300 865.500 233.400 ;
        RECT 863.400 227.400 865.500 228.300 ;
        RECT 866.700 227.400 868.500 234.000 ;
        RECT 833.700 226.500 834.600 227.400 ;
        RECT 833.700 225.600 837.300 226.500 ;
        RECT 831.000 224.400 832.800 224.700 ;
        RECT 791.700 222.300 793.800 223.500 ;
        RECT 777.300 221.400 793.800 222.300 ;
        RECT 797.100 222.600 799.200 223.500 ;
        RECT 813.600 223.200 832.800 224.400 ;
        RECT 813.600 222.600 814.800 223.200 ;
        RECT 831.000 222.900 832.800 223.200 ;
        RECT 797.100 221.400 814.800 222.600 ;
        RECT 817.500 221.700 819.600 222.300 ;
        RECT 827.700 221.700 829.500 222.300 ;
        RECT 777.300 204.600 778.200 221.400 ;
        RECT 817.500 220.500 829.500 221.700 ;
        RECT 779.100 219.300 814.800 220.500 ;
        RECT 817.500 220.200 819.600 220.500 ;
        RECT 779.100 218.700 780.900 219.300 ;
        RECT 813.600 218.700 814.800 219.300 ;
        RECT 782.100 214.950 784.200 217.050 ;
        RECT 782.700 212.100 784.200 214.950 ;
        RECT 786.300 214.800 791.400 216.600 ;
        RECT 790.500 213.300 791.400 214.800 ;
        RECT 794.100 216.300 795.900 218.100 ;
        RECT 800.100 217.800 802.200 218.100 ;
        RECT 813.600 217.800 827.100 218.700 ;
        RECT 794.100 215.100 795.000 216.300 ;
        RECT 800.100 216.000 804.000 217.800 ;
        RECT 805.500 216.300 807.600 217.200 ;
        RECT 825.300 217.050 827.100 217.800 ;
        RECT 805.500 215.100 816.600 216.300 ;
        RECT 825.300 215.250 829.200 217.050 ;
        RECT 794.100 214.200 807.600 215.100 ;
        RECT 814.800 214.500 816.600 215.100 ;
        RECT 827.100 214.950 829.200 215.250 ;
        RECT 833.100 214.950 835.200 217.050 ;
        RECT 833.100 213.300 834.900 214.950 ;
        RECT 790.500 212.100 834.900 213.300 ;
        RECT 782.700 210.600 789.300 212.100 ;
        RECT 779.100 207.900 786.900 209.700 ;
        RECT 787.800 209.100 804.900 210.600 ;
        RECT 802.800 208.500 804.900 209.100 ;
        RECT 809.100 210.000 811.200 211.050 ;
        RECT 809.100 209.100 814.200 210.000 ;
        RECT 817.800 209.400 819.600 211.200 ;
        RECT 836.100 209.400 837.300 225.600 ;
        RECT 854.100 214.050 855.900 215.850 ;
        RECT 857.100 214.050 858.300 227.400 ;
        RECT 863.400 226.500 864.300 227.400 ;
        RECT 860.700 225.600 864.300 226.500 ;
        RECT 853.950 211.950 856.050 214.050 ;
        RECT 856.950 211.950 859.050 214.050 ;
        RECT 809.100 208.950 811.200 209.100 ;
        RECT 785.400 204.600 786.900 207.900 ;
        RECT 803.100 206.700 804.900 208.500 ;
        RECT 812.400 208.200 814.200 209.100 ;
        RECT 818.700 206.400 819.600 209.400 ;
        RECT 820.500 208.200 837.300 209.400 ;
        RECT 820.500 207.300 822.600 208.200 ;
        RECT 831.300 206.700 833.100 207.300 ;
        RECT 791.100 204.600 797.700 206.400 ;
        RECT 812.400 205.200 819.600 206.400 ;
        RECT 824.700 205.500 833.100 206.700 ;
        RECT 812.400 204.600 813.300 205.200 ;
        RECT 815.400 204.600 817.200 205.200 ;
        RECT 824.700 204.600 826.200 205.500 ;
        RECT 836.100 204.600 837.300 208.200 ;
        RECT 844.950 207.450 847.050 208.050 ;
        RECT 853.950 207.450 856.050 208.050 ;
        RECT 844.950 206.550 856.050 207.450 ;
        RECT 844.950 205.950 847.050 206.550 ;
        RECT 853.950 205.950 856.050 206.550 ;
        RECT 777.300 198.600 779.100 204.600 ;
        RECT 782.700 198.000 784.500 204.600 ;
        RECT 785.400 203.400 789.600 204.600 ;
        RECT 787.800 198.600 789.600 203.400 ;
        RECT 791.700 201.600 793.800 203.700 ;
        RECT 794.700 201.600 796.800 203.700 ;
        RECT 797.700 201.600 799.800 203.700 ;
        RECT 800.700 201.600 802.800 203.700 ;
        RECT 806.100 202.500 808.800 204.600 ;
        RECT 810.600 203.400 813.300 204.600 ;
        RECT 810.600 202.500 812.400 203.400 ;
        RECT 792.000 198.600 793.800 201.600 ;
        RECT 795.000 198.600 796.800 201.600 ;
        RECT 798.000 198.600 799.800 201.600 ;
        RECT 801.000 198.600 802.800 201.600 ;
        RECT 804.000 198.000 805.800 201.600 ;
        RECT 807.000 198.600 808.800 202.500 ;
        RECT 814.200 201.600 816.300 203.700 ;
        RECT 817.200 201.600 819.300 203.700 ;
        RECT 820.200 201.600 822.300 203.700 ;
        RECT 811.500 198.000 813.300 201.600 ;
        RECT 814.500 198.600 816.300 201.600 ;
        RECT 817.500 198.600 819.300 201.600 ;
        RECT 820.500 198.600 822.300 201.600 ;
        RECT 824.700 198.600 826.500 204.600 ;
        RECT 830.100 198.000 831.900 204.600 ;
        RECT 835.500 198.600 837.300 204.600 ;
        RECT 857.100 201.600 858.300 211.950 ;
        RECT 860.700 209.400 861.900 225.600 ;
        RECT 865.200 224.400 867.000 224.700 ;
        RECT 869.700 224.400 871.500 233.400 ;
        RECT 872.700 227.400 874.500 234.000 ;
        RECT 876.300 230.400 878.100 233.400 ;
        RECT 879.300 230.400 881.100 233.400 ;
        RECT 876.300 228.300 878.400 230.400 ;
        RECT 879.300 228.300 881.400 230.400 ;
        RECT 882.300 227.400 884.100 233.400 ;
        RECT 885.300 227.400 887.100 234.000 ;
        RECT 881.700 225.300 883.800 227.400 ;
        RECT 889.200 225.900 891.000 233.400 ;
        RECT 892.200 227.400 894.000 234.000 ;
        RECT 895.200 227.400 897.000 233.400 ;
        RECT 898.200 230.400 900.000 233.400 ;
        RECT 901.200 230.400 903.000 233.400 ;
        RECT 904.200 230.400 906.000 233.400 ;
        RECT 898.200 228.300 900.300 230.400 ;
        RECT 901.200 228.300 903.300 230.400 ;
        RECT 904.200 228.300 906.300 230.400 ;
        RECT 907.200 227.400 909.000 234.000 ;
        RECT 910.200 227.400 912.000 233.400 ;
        RECT 913.200 227.400 915.000 234.000 ;
        RECT 916.200 227.400 918.000 233.400 ;
        RECT 919.200 227.400 921.000 234.000 ;
        RECT 922.500 227.400 924.300 233.400 ;
        RECT 925.500 227.400 927.300 234.000 ;
        RECT 944.700 227.400 946.500 234.000 ;
        RECT 865.200 223.200 884.400 224.400 ;
        RECT 889.200 223.800 892.500 225.900 ;
        RECT 895.200 223.500 897.900 227.400 ;
        RECT 901.200 226.500 903.300 227.400 ;
        RECT 901.200 225.300 909.300 226.500 ;
        RECT 907.500 224.700 909.300 225.300 ;
        RECT 910.200 224.400 911.400 227.400 ;
        RECT 916.800 226.500 918.000 227.400 ;
        RECT 916.800 225.600 920.700 226.500 ;
        RECT 914.100 224.400 915.900 225.000 ;
        RECT 865.200 222.900 867.000 223.200 ;
        RECT 883.200 222.600 884.400 223.200 ;
        RECT 898.800 222.600 900.900 223.500 ;
        RECT 868.500 221.700 870.300 222.300 ;
        RECT 878.400 221.700 880.500 222.300 ;
        RECT 868.500 220.500 880.500 221.700 ;
        RECT 883.200 221.400 900.900 222.600 ;
        RECT 904.200 222.300 906.300 223.500 ;
        RECT 910.200 223.200 915.900 224.400 ;
        RECT 919.800 222.300 920.700 225.600 ;
        RECT 904.200 221.400 920.700 222.300 ;
        RECT 878.400 220.200 880.500 220.500 ;
        RECT 883.200 219.300 918.900 220.500 ;
        RECT 883.200 218.700 884.400 219.300 ;
        RECT 917.100 218.700 918.900 219.300 ;
        RECT 870.900 217.800 884.400 218.700 ;
        RECT 895.800 217.800 897.900 218.100 ;
        RECT 870.900 217.050 872.700 217.800 ;
        RECT 862.800 214.950 864.900 217.050 ;
        RECT 868.800 215.250 872.700 217.050 ;
        RECT 890.400 216.300 892.500 217.200 ;
        RECT 868.800 214.950 870.900 215.250 ;
        RECT 881.400 215.100 892.500 216.300 ;
        RECT 894.000 216.000 897.900 217.800 ;
        RECT 902.100 216.300 903.900 218.100 ;
        RECT 903.000 215.100 903.900 216.300 ;
        RECT 863.100 213.300 864.900 214.950 ;
        RECT 881.400 214.500 883.200 215.100 ;
        RECT 890.400 214.200 903.900 215.100 ;
        RECT 906.600 214.800 911.700 216.600 ;
        RECT 913.800 214.950 915.900 217.050 ;
        RECT 906.600 213.300 907.500 214.800 ;
        RECT 863.100 212.100 907.500 213.300 ;
        RECT 913.800 212.100 915.300 214.950 ;
        RECT 878.400 209.400 880.200 211.200 ;
        RECT 886.800 210.000 888.900 211.050 ;
        RECT 908.700 210.600 915.300 212.100 ;
        RECT 860.700 208.200 877.500 209.400 ;
        RECT 860.700 204.600 861.900 208.200 ;
        RECT 875.400 207.300 877.500 208.200 ;
        RECT 864.900 206.700 866.700 207.300 ;
        RECT 864.900 205.500 873.300 206.700 ;
        RECT 871.800 204.600 873.300 205.500 ;
        RECT 878.400 206.400 879.300 209.400 ;
        RECT 883.800 209.100 888.900 210.000 ;
        RECT 883.800 208.200 885.600 209.100 ;
        RECT 886.800 208.950 888.900 209.100 ;
        RECT 893.100 209.100 910.200 210.600 ;
        RECT 893.100 208.500 895.200 209.100 ;
        RECT 893.100 206.700 894.900 208.500 ;
        RECT 911.100 207.900 918.900 209.700 ;
        RECT 878.400 205.200 885.600 206.400 ;
        RECT 880.800 204.600 882.600 205.200 ;
        RECT 884.700 204.600 885.600 205.200 ;
        RECT 900.300 204.600 906.900 206.400 ;
        RECT 911.100 204.600 912.600 207.900 ;
        RECT 919.800 204.600 920.700 221.400 ;
        RECT 854.100 198.000 855.900 201.600 ;
        RECT 857.100 198.600 858.900 201.600 ;
        RECT 860.700 198.600 862.500 204.600 ;
        RECT 866.100 198.000 867.900 204.600 ;
        RECT 871.500 198.600 873.300 204.600 ;
        RECT 875.700 201.600 877.800 203.700 ;
        RECT 878.700 201.600 880.800 203.700 ;
        RECT 881.700 201.600 883.800 203.700 ;
        RECT 884.700 203.400 887.400 204.600 ;
        RECT 885.600 202.500 887.400 203.400 ;
        RECT 889.200 202.500 891.900 204.600 ;
        RECT 875.700 198.600 877.500 201.600 ;
        RECT 878.700 198.600 880.500 201.600 ;
        RECT 881.700 198.600 883.500 201.600 ;
        RECT 884.700 198.000 886.500 201.600 ;
        RECT 889.200 198.600 891.000 202.500 ;
        RECT 895.200 201.600 897.300 203.700 ;
        RECT 898.200 201.600 900.300 203.700 ;
        RECT 901.200 201.600 903.300 203.700 ;
        RECT 904.200 201.600 906.300 203.700 ;
        RECT 908.400 203.400 912.600 204.600 ;
        RECT 892.200 198.000 894.000 201.600 ;
        RECT 895.200 198.600 897.000 201.600 ;
        RECT 898.200 198.600 900.000 201.600 ;
        RECT 901.200 198.600 903.000 201.600 ;
        RECT 904.200 198.600 906.000 201.600 ;
        RECT 908.400 198.600 910.200 203.400 ;
        RECT 913.500 198.000 915.300 204.600 ;
        RECT 918.900 198.600 920.700 204.600 ;
        RECT 922.500 217.050 924.000 227.400 ;
        RECT 945.000 224.100 946.800 225.900 ;
        RECT 947.700 222.900 949.500 233.400 ;
        RECT 947.100 221.400 949.500 222.900 ;
        RECT 952.800 221.400 954.600 234.000 ;
        RECT 971.100 227.400 972.900 234.000 ;
        RECT 974.100 227.400 975.900 233.400 ;
        RECT 922.500 214.950 924.900 217.050 ;
        RECT 922.500 201.600 924.000 214.950 ;
        RECT 947.100 214.050 948.300 221.400 ;
        RECT 949.950 219.450 952.050 220.200 ;
        RECT 958.950 219.450 961.050 220.050 ;
        RECT 949.950 218.550 961.050 219.450 ;
        RECT 949.950 218.100 952.050 218.550 ;
        RECT 958.950 217.950 961.050 218.550 ;
        RECT 953.100 214.050 954.900 215.850 ;
        RECT 971.100 214.050 972.900 215.850 ;
        RECT 974.100 214.050 975.300 227.400 ;
        RECT 992.100 221.400 993.900 234.000 ;
        RECT 997.200 222.600 999.000 233.400 ;
        RECT 1016.100 227.400 1017.900 234.000 ;
        RECT 1019.100 227.400 1020.900 233.400 ;
        RECT 1022.100 227.400 1023.900 234.000 ;
        RECT 995.400 221.400 999.000 222.600 ;
        RECT 992.250 214.050 994.050 215.850 ;
        RECT 995.400 214.050 996.300 221.400 ;
        RECT 998.100 214.050 999.900 215.850 ;
        RECT 1019.100 214.050 1020.300 227.400 ;
        RECT 943.950 211.950 946.050 214.050 ;
        RECT 946.950 211.950 949.050 214.050 ;
        RECT 949.950 211.950 952.050 214.050 ;
        RECT 952.950 211.950 955.050 214.050 ;
        RECT 970.950 211.950 973.050 214.050 ;
        RECT 973.950 211.950 976.050 214.050 ;
        RECT 991.950 211.950 994.050 214.050 ;
        RECT 994.950 211.950 997.050 214.050 ;
        RECT 997.950 211.950 1000.050 214.050 ;
        RECT 1015.950 211.950 1018.050 214.050 ;
        RECT 1018.950 211.950 1021.050 214.050 ;
        RECT 1021.950 211.950 1024.050 214.050 ;
        RECT 944.100 210.150 945.900 211.950 ;
        RECT 947.100 207.600 948.300 211.950 ;
        RECT 950.100 210.150 951.900 211.950 ;
        RECT 944.700 206.700 948.300 207.600 ;
        RECT 944.700 204.600 945.900 206.700 ;
        RECT 922.500 198.600 924.300 201.600 ;
        RECT 925.500 198.000 927.300 201.600 ;
        RECT 944.100 198.600 945.900 204.600 ;
        RECT 947.100 203.700 954.900 205.050 ;
        RECT 947.100 198.600 948.900 203.700 ;
        RECT 950.100 198.000 951.900 202.800 ;
        RECT 953.100 198.600 954.900 203.700 ;
        RECT 974.100 201.600 975.300 211.950 ;
        RECT 995.400 201.600 996.300 211.950 ;
        RECT 1016.250 210.150 1018.050 211.950 ;
        RECT 1019.100 206.700 1020.300 211.950 ;
        RECT 1022.100 210.150 1023.900 211.950 ;
        RECT 1019.100 205.800 1023.300 206.700 ;
        RECT 971.100 198.000 972.900 201.600 ;
        RECT 974.100 198.600 975.900 201.600 ;
        RECT 992.100 198.000 993.900 201.600 ;
        RECT 995.100 198.600 996.900 201.600 ;
        RECT 998.100 198.000 999.900 201.600 ;
        RECT 1016.400 198.000 1018.200 204.600 ;
        RECT 1021.500 198.600 1023.300 205.800 ;
        RECT 17.100 188.400 18.900 195.000 ;
        RECT 20.100 188.400 21.900 194.400 ;
        RECT 38.100 189.300 39.900 194.400 ;
        RECT 41.100 190.200 42.900 195.000 ;
        RECT 44.100 189.300 45.900 194.400 ;
        RECT 17.100 181.050 18.900 182.850 ;
        RECT 20.100 181.050 21.300 188.400 ;
        RECT 38.100 187.950 45.900 189.300 ;
        RECT 47.100 188.400 48.900 194.400 ;
        RECT 65.400 188.400 67.200 195.000 ;
        RECT 47.100 186.300 48.300 188.400 ;
        RECT 70.500 187.200 72.300 194.400 ;
        RECT 89.100 191.400 90.900 195.000 ;
        RECT 92.100 191.400 93.900 194.400 ;
        RECT 95.100 191.400 96.900 195.000 ;
        RECT 44.700 185.400 48.300 186.300 ;
        RECT 68.100 186.300 72.300 187.200 ;
        RECT 41.100 181.050 42.900 182.850 ;
        RECT 44.700 181.050 45.900 185.400 ;
        RECT 47.100 181.050 48.900 182.850 ;
        RECT 65.250 181.050 67.050 182.850 ;
        RECT 68.100 181.050 69.300 186.300 ;
        RECT 71.100 181.050 72.900 182.850 ;
        RECT 92.400 181.050 93.300 191.400 ;
        RECT 113.700 187.200 115.500 194.400 ;
        RECT 118.800 188.400 120.600 195.000 ;
        RECT 137.700 187.200 139.500 194.400 ;
        RECT 142.800 188.400 144.600 195.000 ;
        RECT 161.100 194.400 162.300 195.000 ;
        RECT 161.100 191.400 162.900 194.400 ;
        RECT 164.100 191.400 165.900 194.400 ;
        RECT 164.400 187.200 165.300 191.400 ;
        RECT 167.100 189.000 168.900 195.000 ;
        RECT 170.100 188.400 171.900 194.400 ;
        RECT 188.400 188.400 190.200 195.000 ;
        RECT 113.700 186.300 117.900 187.200 ;
        RECT 137.700 186.300 141.900 187.200 ;
        RECT 164.400 186.300 169.800 187.200 ;
        RECT 113.100 181.050 114.900 182.850 ;
        RECT 116.700 181.050 117.900 186.300 ;
        RECT 118.950 181.050 120.750 182.850 ;
        RECT 137.100 181.050 138.900 182.850 ;
        RECT 140.700 181.050 141.900 186.300 ;
        RECT 167.700 185.400 169.800 186.300 ;
        RECT 142.950 181.050 144.750 182.850 ;
        RECT 161.400 181.050 163.200 182.850 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 70.950 178.950 73.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 161.100 178.950 163.200 181.050 ;
        RECT 164.400 178.950 166.500 181.050 ;
        RECT 20.100 171.600 21.300 178.950 ;
        RECT 38.100 177.150 39.900 178.950 ;
        RECT 44.700 171.600 45.900 178.950 ;
        RECT 17.100 159.000 18.900 171.600 ;
        RECT 20.100 159.600 21.900 171.600 ;
        RECT 38.400 159.000 40.200 171.600 ;
        RECT 43.500 170.100 45.900 171.600 ;
        RECT 43.500 159.600 45.300 170.100 ;
        RECT 46.200 167.100 48.000 168.900 ;
        RECT 68.100 165.600 69.300 178.950 ;
        RECT 89.250 177.150 91.050 178.950 ;
        RECT 92.400 171.600 93.300 178.950 ;
        RECT 95.100 177.150 96.900 178.950 ;
        RECT 46.500 159.000 48.300 165.600 ;
        RECT 65.100 159.000 66.900 165.600 ;
        RECT 68.100 159.600 69.900 165.600 ;
        RECT 71.100 159.000 72.900 165.600 ;
        RECT 89.100 159.000 90.900 171.600 ;
        RECT 92.400 170.400 96.000 171.600 ;
        RECT 94.200 159.600 96.000 170.400 ;
        RECT 116.700 165.600 117.900 178.950 ;
        RECT 121.950 174.450 124.050 175.050 ;
        RECT 130.950 174.450 133.050 175.050 ;
        RECT 136.950 174.450 139.050 175.050 ;
        RECT 121.950 173.550 139.050 174.450 ;
        RECT 121.950 172.950 124.050 173.550 ;
        RECT 130.950 172.950 133.050 173.550 ;
        RECT 136.950 172.950 139.050 173.550 ;
        RECT 140.700 165.600 141.900 178.950 ;
        RECT 165.000 177.150 166.800 178.950 ;
        RECT 142.950 174.450 145.050 175.050 ;
        RECT 154.950 174.450 157.050 175.050 ;
        RECT 167.700 174.900 168.600 185.400 ;
        RECT 171.000 181.050 171.900 188.400 ;
        RECT 193.500 187.200 195.300 194.400 ;
        RECT 191.100 186.300 195.300 187.200 ;
        RECT 188.250 181.050 190.050 182.850 ;
        RECT 191.100 181.050 192.300 186.300 ;
        RECT 214.500 186.000 216.300 194.400 ;
        RECT 213.000 184.800 216.300 186.000 ;
        RECT 221.100 185.400 222.900 195.000 ;
        RECT 239.400 188.400 241.200 195.000 ;
        RECT 244.500 187.200 246.300 194.400 ;
        RECT 265.500 188.400 267.300 195.000 ;
        RECT 270.000 188.400 271.800 194.400 ;
        RECT 274.500 188.400 276.300 195.000 ;
        RECT 293.700 191.400 295.500 195.000 ;
        RECT 296.700 189.600 298.500 194.400 ;
        RECT 293.400 188.400 298.500 189.600 ;
        RECT 301.200 188.400 303.000 195.000 ;
        RECT 320.100 188.400 321.900 194.400 ;
        RECT 242.100 186.300 246.300 187.200 ;
        RECT 194.100 181.050 195.900 182.850 ;
        RECT 213.000 181.050 213.900 184.800 ;
        RECT 215.100 181.050 216.900 182.850 ;
        RECT 221.100 181.050 222.900 182.850 ;
        RECT 239.250 181.050 241.050 182.850 ;
        RECT 242.100 181.050 243.300 186.300 ;
        RECT 245.100 181.050 246.900 182.850 ;
        RECT 263.100 181.050 264.900 182.850 ;
        RECT 269.700 181.050 270.900 188.400 ;
        RECT 274.950 181.050 276.750 182.850 ;
        RECT 293.400 181.050 294.300 188.400 ;
        RECT 320.700 186.300 321.900 188.400 ;
        RECT 323.100 189.300 324.900 194.400 ;
        RECT 326.100 190.200 327.900 195.000 ;
        RECT 329.100 189.300 330.900 194.400 ;
        RECT 323.100 187.950 330.900 189.300 ;
        RECT 347.100 188.400 348.900 194.400 ;
        RECT 347.700 186.300 348.900 188.400 ;
        RECT 350.100 189.300 351.900 194.400 ;
        RECT 353.100 190.200 354.900 195.000 ;
        RECT 356.100 189.300 357.900 194.400 ;
        RECT 374.100 191.400 375.900 194.400 ;
        RECT 377.100 191.400 378.900 195.000 ;
        RECT 350.100 187.950 357.900 189.300 ;
        RECT 320.700 185.400 324.300 186.300 ;
        RECT 347.700 185.400 351.300 186.300 ;
        RECT 295.950 181.050 297.750 182.850 ;
        RECT 302.100 181.050 303.900 182.850 ;
        RECT 320.100 181.050 321.900 182.850 ;
        RECT 323.100 181.050 324.300 185.400 ;
        RECT 326.100 181.050 327.900 182.850 ;
        RECT 347.100 181.050 348.900 182.850 ;
        RECT 350.100 181.050 351.300 185.400 ;
        RECT 358.950 183.450 363.000 184.050 ;
        RECT 353.100 181.050 354.900 182.850 ;
        RECT 358.950 181.950 363.450 183.450 ;
        RECT 169.800 178.950 171.900 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 142.950 173.550 157.050 174.450 ;
        RECT 167.100 174.300 168.900 174.900 ;
        RECT 142.950 172.950 145.050 173.550 ;
        RECT 154.950 172.950 157.050 173.550 ;
        RECT 161.100 173.100 168.900 174.300 ;
        RECT 161.100 171.600 162.300 173.100 ;
        RECT 169.800 171.600 171.000 178.950 ;
        RECT 175.950 174.450 178.050 175.050 ;
        RECT 187.950 174.450 190.050 175.050 ;
        RECT 175.950 173.550 190.050 174.450 ;
        RECT 175.950 172.950 178.050 173.550 ;
        RECT 187.950 172.950 190.050 173.550 ;
        RECT 113.100 159.000 114.900 165.600 ;
        RECT 116.100 159.600 117.900 165.600 ;
        RECT 119.100 159.000 120.900 165.600 ;
        RECT 137.100 159.000 138.900 165.600 ;
        RECT 140.100 159.600 141.900 165.600 ;
        RECT 143.100 159.000 144.900 165.600 ;
        RECT 161.100 159.600 162.900 171.600 ;
        RECT 165.600 159.000 167.400 171.600 ;
        RECT 168.600 170.100 171.000 171.600 ;
        RECT 168.600 159.600 170.400 170.100 ;
        RECT 191.100 165.600 192.300 178.950 ;
        RECT 213.000 166.800 213.900 178.950 ;
        RECT 218.100 177.150 219.900 178.950 ;
        RECT 213.000 165.900 219.600 166.800 ;
        RECT 213.000 165.600 213.900 165.900 ;
        RECT 188.100 159.000 189.900 165.600 ;
        RECT 191.100 159.600 192.900 165.600 ;
        RECT 194.100 159.000 195.900 165.600 ;
        RECT 212.100 159.600 213.900 165.600 ;
        RECT 218.100 165.600 219.600 165.900 ;
        RECT 242.100 165.600 243.300 178.950 ;
        RECT 266.100 177.150 267.900 178.950 ;
        RECT 270.000 173.400 270.900 178.950 ;
        RECT 271.950 177.150 273.750 178.950 ;
        RECT 266.100 172.500 270.900 173.400 ;
        RECT 215.100 159.000 216.900 165.000 ;
        RECT 218.100 159.600 219.900 165.600 ;
        RECT 221.100 159.000 222.900 165.600 ;
        RECT 239.100 159.000 240.900 165.600 ;
        RECT 242.100 159.600 243.900 165.600 ;
        RECT 245.100 159.000 246.900 165.600 ;
        RECT 263.100 160.500 264.900 171.600 ;
        RECT 266.100 161.400 267.900 172.500 ;
        RECT 293.400 171.600 294.300 178.950 ;
        RECT 298.950 177.150 300.750 178.950 ;
        RECT 295.950 174.450 298.050 175.050 ;
        RECT 307.950 174.450 310.050 175.050 ;
        RECT 295.950 173.550 310.050 174.450 ;
        RECT 295.950 172.950 298.050 173.550 ;
        RECT 307.950 172.950 310.050 173.550 ;
        RECT 323.100 171.600 324.300 178.950 ;
        RECT 329.100 177.150 330.900 178.950 ;
        RECT 350.100 171.600 351.300 178.950 ;
        RECT 356.100 177.150 357.900 178.950 ;
        RECT 362.550 178.050 363.450 181.950 ;
        RECT 374.700 181.050 375.900 191.400 ;
        RECT 395.100 189.300 396.900 194.400 ;
        RECT 398.100 190.200 399.900 195.000 ;
        RECT 401.100 189.300 402.900 194.400 ;
        RECT 395.100 187.950 402.900 189.300 ;
        RECT 404.100 188.400 405.900 194.400 ;
        RECT 423.000 188.400 424.800 195.000 ;
        RECT 427.500 189.600 429.300 194.400 ;
        RECT 430.500 191.400 432.300 195.000 ;
        RECT 449.100 191.400 450.900 195.000 ;
        RECT 452.100 191.400 453.900 194.400 ;
        RECT 455.100 191.400 456.900 195.000 ;
        RECT 427.500 188.400 432.600 189.600 ;
        RECT 404.100 186.300 405.300 188.400 ;
        RECT 401.700 185.400 405.300 186.300 ;
        RECT 398.100 181.050 399.900 182.850 ;
        RECT 401.700 181.050 402.900 185.400 ;
        RECT 404.100 181.050 405.900 182.850 ;
        RECT 422.100 181.050 423.900 182.850 ;
        RECT 428.250 181.050 430.050 182.850 ;
        RECT 431.700 181.050 432.600 188.400 ;
        RECT 433.950 183.450 438.000 184.050 ;
        RECT 433.950 181.950 438.450 183.450 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 397.950 178.950 400.050 181.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 358.950 176.550 363.450 178.050 ;
        RECT 358.950 175.950 363.000 176.550 ;
        RECT 269.100 170.400 276.900 171.300 ;
        RECT 269.100 160.500 270.900 170.400 ;
        RECT 263.100 159.600 270.900 160.500 ;
        RECT 272.100 159.000 273.900 169.500 ;
        RECT 275.100 159.600 276.900 170.400 ;
        RECT 293.100 159.600 294.900 171.600 ;
        RECT 296.100 170.700 303.900 171.600 ;
        RECT 296.100 159.600 297.900 170.700 ;
        RECT 299.100 159.000 300.900 169.800 ;
        RECT 302.100 159.600 303.900 170.700 ;
        RECT 323.100 170.100 325.500 171.600 ;
        RECT 321.000 167.100 322.800 168.900 ;
        RECT 320.700 159.000 322.500 165.600 ;
        RECT 323.700 159.600 325.500 170.100 ;
        RECT 328.800 159.000 330.600 171.600 ;
        RECT 350.100 170.100 352.500 171.600 ;
        RECT 348.000 167.100 349.800 168.900 ;
        RECT 347.700 159.000 349.500 165.600 ;
        RECT 350.700 159.600 352.500 170.100 ;
        RECT 355.800 159.000 357.600 171.600 ;
        RECT 374.700 165.600 375.900 178.950 ;
        RECT 377.100 177.150 378.900 178.950 ;
        RECT 395.100 177.150 396.900 178.950 ;
        RECT 376.950 174.450 379.050 175.050 ;
        RECT 382.950 174.450 385.050 175.050 ;
        RECT 397.950 174.450 400.050 175.050 ;
        RECT 376.950 173.550 400.050 174.450 ;
        RECT 376.950 172.950 379.050 173.550 ;
        RECT 382.950 172.950 385.050 173.550 ;
        RECT 397.950 172.950 400.050 173.550 ;
        RECT 401.700 171.600 402.900 178.950 ;
        RECT 425.250 177.150 427.050 178.950 ;
        RECT 409.950 174.450 412.050 175.050 ;
        RECT 421.950 174.450 424.050 175.050 ;
        RECT 409.950 173.550 424.050 174.450 ;
        RECT 409.950 172.950 412.050 173.550 ;
        RECT 421.950 172.950 424.050 173.550 ;
        RECT 431.700 171.600 432.600 178.950 ;
        RECT 437.550 177.450 438.450 181.950 ;
        RECT 452.400 181.050 453.300 191.400 ;
        RECT 458.700 188.400 460.500 194.400 ;
        RECT 464.100 188.400 465.900 195.000 ;
        RECT 469.500 188.400 471.300 194.400 ;
        RECT 473.700 191.400 475.500 194.400 ;
        RECT 476.700 191.400 478.500 194.400 ;
        RECT 479.700 191.400 481.500 194.400 ;
        RECT 482.700 191.400 484.500 195.000 ;
        RECT 473.700 189.300 475.800 191.400 ;
        RECT 476.700 189.300 478.800 191.400 ;
        RECT 479.700 189.300 481.800 191.400 ;
        RECT 487.200 190.500 489.000 194.400 ;
        RECT 490.200 191.400 492.000 195.000 ;
        RECT 493.200 191.400 495.000 194.400 ;
        RECT 496.200 191.400 498.000 194.400 ;
        RECT 499.200 191.400 501.000 194.400 ;
        RECT 502.200 191.400 504.000 194.400 ;
        RECT 483.600 189.600 485.400 190.500 ;
        RECT 482.700 188.400 485.400 189.600 ;
        RECT 487.200 188.400 489.900 190.500 ;
        RECT 493.200 189.300 495.300 191.400 ;
        RECT 496.200 189.300 498.300 191.400 ;
        RECT 499.200 189.300 501.300 191.400 ;
        RECT 502.200 189.300 504.300 191.400 ;
        RECT 506.400 189.600 508.200 194.400 ;
        RECT 506.400 188.400 510.600 189.600 ;
        RECT 511.500 188.400 513.300 195.000 ;
        RECT 516.900 188.400 518.700 194.400 ;
        RECT 458.700 184.800 459.900 188.400 ;
        RECT 469.800 187.500 471.300 188.400 ;
        RECT 478.800 187.800 480.600 188.400 ;
        RECT 482.700 187.800 483.600 188.400 ;
        RECT 462.900 186.300 471.300 187.500 ;
        RECT 476.400 186.600 483.600 187.800 ;
        RECT 498.300 186.600 504.900 188.400 ;
        RECT 462.900 185.700 464.700 186.300 ;
        RECT 473.400 184.800 475.500 185.700 ;
        RECT 458.700 183.600 475.500 184.800 ;
        RECT 476.400 183.600 477.300 186.600 ;
        RECT 481.800 183.900 483.600 184.800 ;
        RECT 491.100 184.500 492.900 186.300 ;
        RECT 509.100 185.100 510.600 188.400 ;
        RECT 484.800 183.900 486.900 184.050 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 445.950 177.450 448.050 178.050 ;
        RECT 437.550 176.550 448.050 177.450 ;
        RECT 449.250 177.150 451.050 178.950 ;
        RECT 445.950 175.950 448.050 176.550 ;
        RECT 452.400 171.600 453.300 178.950 ;
        RECT 455.100 177.150 456.900 178.950 ;
        RECT 374.100 159.600 375.900 165.600 ;
        RECT 377.100 159.000 378.900 165.600 ;
        RECT 395.400 159.000 397.200 171.600 ;
        RECT 400.500 170.100 402.900 171.600 ;
        RECT 422.100 170.700 429.900 171.600 ;
        RECT 400.500 159.600 402.300 170.100 ;
        RECT 403.200 167.100 405.000 168.900 ;
        RECT 403.500 159.000 405.300 165.600 ;
        RECT 422.100 159.600 423.900 170.700 ;
        RECT 425.100 159.000 426.900 169.800 ;
        RECT 428.100 159.600 429.900 170.700 ;
        RECT 431.100 159.600 432.900 171.600 ;
        RECT 449.100 159.000 450.900 171.600 ;
        RECT 452.400 170.400 456.000 171.600 ;
        RECT 454.200 159.600 456.000 170.400 ;
        RECT 458.700 167.400 459.900 183.600 ;
        RECT 476.400 181.800 478.200 183.600 ;
        RECT 481.800 183.000 486.900 183.900 ;
        RECT 484.800 181.950 486.900 183.000 ;
        RECT 491.100 183.900 493.200 184.500 ;
        RECT 491.100 182.400 508.200 183.900 ;
        RECT 509.100 183.300 516.900 185.100 ;
        RECT 506.700 180.900 513.300 182.400 ;
        RECT 461.100 179.700 505.500 180.900 ;
        RECT 461.100 178.050 462.900 179.700 ;
        RECT 460.800 175.950 462.900 178.050 ;
        RECT 466.800 177.750 468.900 178.050 ;
        RECT 479.400 177.900 481.200 178.500 ;
        RECT 488.400 177.900 501.900 178.800 ;
        RECT 466.800 175.950 470.700 177.750 ;
        RECT 479.400 176.700 490.500 177.900 ;
        RECT 468.900 175.200 470.700 175.950 ;
        RECT 488.400 175.800 490.500 176.700 ;
        RECT 492.000 175.200 495.900 177.000 ;
        RECT 501.000 176.700 501.900 177.900 ;
        RECT 468.900 174.300 482.400 175.200 ;
        RECT 493.800 174.900 495.900 175.200 ;
        RECT 500.100 174.900 501.900 176.700 ;
        RECT 504.600 178.200 505.500 179.700 ;
        RECT 504.600 176.400 509.700 178.200 ;
        RECT 511.800 178.050 513.300 180.900 ;
        RECT 511.800 175.950 513.900 178.050 ;
        RECT 481.200 173.700 482.400 174.300 ;
        RECT 515.100 173.700 516.900 174.300 ;
        RECT 476.400 172.500 478.500 172.800 ;
        RECT 481.200 172.500 516.900 173.700 ;
        RECT 466.500 171.300 478.500 172.500 ;
        RECT 517.800 171.600 518.700 188.400 ;
        RECT 466.500 170.700 468.300 171.300 ;
        RECT 476.400 170.700 478.500 171.300 ;
        RECT 481.200 170.400 498.900 171.600 ;
        RECT 463.200 169.800 465.000 170.100 ;
        RECT 481.200 169.800 482.400 170.400 ;
        RECT 463.200 168.600 482.400 169.800 ;
        RECT 496.800 169.500 498.900 170.400 ;
        RECT 502.200 170.700 518.700 171.600 ;
        RECT 502.200 169.500 504.300 170.700 ;
        RECT 463.200 168.300 465.000 168.600 ;
        RECT 458.700 166.500 462.300 167.400 ;
        RECT 461.400 165.600 462.300 166.500 ;
        RECT 458.700 159.000 460.500 165.600 ;
        RECT 461.400 164.700 463.500 165.600 ;
        RECT 461.700 159.600 463.500 164.700 ;
        RECT 464.700 159.000 466.500 165.600 ;
        RECT 467.700 159.600 469.500 168.600 ;
        RECT 479.700 165.600 481.800 167.700 ;
        RECT 487.200 167.100 490.500 169.200 ;
        RECT 470.700 159.000 472.500 165.600 ;
        RECT 474.300 162.600 476.400 164.700 ;
        RECT 477.300 162.600 479.400 164.700 ;
        RECT 474.300 159.600 476.100 162.600 ;
        RECT 477.300 159.600 479.100 162.600 ;
        RECT 480.300 159.600 482.100 165.600 ;
        RECT 483.300 159.000 485.100 165.600 ;
        RECT 487.200 159.600 489.000 167.100 ;
        RECT 493.200 165.600 495.900 169.500 ;
        RECT 508.200 168.600 513.900 169.800 ;
        RECT 505.500 167.700 507.300 168.300 ;
        RECT 499.200 166.500 507.300 167.700 ;
        RECT 499.200 165.600 501.300 166.500 ;
        RECT 508.200 165.600 509.400 168.600 ;
        RECT 512.100 168.000 513.900 168.600 ;
        RECT 517.800 167.400 518.700 170.700 ;
        RECT 514.800 166.500 518.700 167.400 ;
        RECT 520.500 191.400 522.300 194.400 ;
        RECT 523.500 191.400 525.300 195.000 ;
        RECT 520.500 178.050 522.000 191.400 ;
        RECT 542.100 188.400 543.900 195.000 ;
        RECT 545.100 187.500 546.900 194.400 ;
        RECT 548.100 188.400 549.900 195.000 ;
        RECT 551.100 187.500 552.900 194.400 ;
        RECT 554.100 188.400 555.900 195.000 ;
        RECT 557.100 187.500 558.900 194.400 ;
        RECT 560.100 188.400 561.900 195.000 ;
        RECT 563.100 187.500 564.900 194.400 ;
        RECT 566.100 188.400 567.900 195.000 ;
        RECT 544.050 186.300 546.900 187.500 ;
        RECT 549.000 186.300 552.900 187.500 ;
        RECT 555.000 186.300 558.900 187.500 ;
        RECT 561.000 186.300 564.900 187.500 ;
        RECT 544.050 181.050 545.100 186.300 ;
        RECT 549.000 185.400 550.200 186.300 ;
        RECT 555.000 185.400 556.200 186.300 ;
        RECT 561.000 185.400 562.200 186.300 ;
        RECT 586.500 186.000 588.300 194.400 ;
        RECT 546.000 184.200 550.200 185.400 ;
        RECT 546.000 183.600 547.800 184.200 ;
        RECT 544.050 178.950 547.200 181.050 ;
        RECT 520.500 175.950 522.900 178.050 ;
        RECT 514.800 165.600 516.000 166.500 ;
        RECT 520.500 165.600 522.000 175.950 ;
        RECT 544.050 173.700 545.100 178.950 ;
        RECT 549.000 173.700 550.200 184.200 ;
        RECT 552.000 184.200 556.200 185.400 ;
        RECT 552.000 183.600 553.800 184.200 ;
        RECT 555.000 173.700 556.200 184.200 ;
        RECT 558.000 184.200 562.200 185.400 ;
        RECT 558.000 183.600 559.800 184.200 ;
        RECT 561.000 173.700 562.200 184.200 ;
        RECT 585.000 184.800 588.300 186.000 ;
        RECT 593.100 185.400 594.900 195.000 ;
        RECT 611.100 191.400 612.900 195.000 ;
        RECT 614.100 191.400 615.900 194.400 ;
        RECT 617.100 191.400 618.900 195.000 ;
        RECT 563.400 181.050 565.200 182.850 ;
        RECT 585.000 181.050 585.900 184.800 ;
        RECT 587.100 181.050 588.900 182.850 ;
        RECT 593.100 181.050 594.900 182.850 ;
        RECT 614.400 181.050 615.300 191.400 ;
        RECT 637.500 186.000 639.300 194.400 ;
        RECT 636.000 184.800 639.300 186.000 ;
        RECT 644.100 185.400 645.900 195.000 ;
        RECT 662.100 188.400 663.900 195.000 ;
        RECT 665.100 188.400 666.900 194.400 ;
        RECT 636.000 181.050 636.900 184.800 ;
        RECT 638.100 181.050 639.900 182.850 ;
        RECT 644.100 181.050 645.900 182.850 ;
        RECT 662.100 181.050 663.900 182.850 ;
        RECT 665.100 181.050 666.300 188.400 ;
        RECT 685.500 186.000 687.300 194.400 ;
        RECT 684.000 184.800 687.300 186.000 ;
        RECT 692.100 185.400 693.900 195.000 ;
        RECT 710.100 191.400 711.900 194.400 ;
        RECT 713.100 191.400 714.900 195.000 ;
        RECT 684.000 181.050 684.900 184.800 ;
        RECT 686.100 181.050 687.900 182.850 ;
        RECT 692.100 181.050 693.900 182.850 ;
        RECT 710.700 181.050 711.900 191.400 ;
        RECT 731.100 188.400 732.900 194.400 ;
        RECT 734.100 189.300 735.900 195.000 ;
        RECT 738.600 188.400 740.400 194.400 ;
        RECT 743.100 189.300 744.900 195.000 ;
        RECT 746.100 188.400 747.900 194.400 ;
        RECT 731.700 186.600 732.900 188.400 ;
        RECT 738.900 186.900 740.100 188.400 ;
        RECT 743.100 187.500 747.900 188.400 ;
        RECT 764.100 189.300 765.900 194.400 ;
        RECT 767.100 190.200 768.900 195.000 ;
        RECT 770.100 189.300 771.900 194.400 ;
        RECT 764.100 187.950 771.900 189.300 ;
        RECT 773.100 188.400 774.900 194.400 ;
        RECT 791.100 191.400 792.900 194.400 ;
        RECT 794.100 191.400 795.900 195.000 ;
        RECT 812.100 191.400 813.900 195.000 ;
        RECT 815.100 191.400 816.900 194.400 ;
        RECT 818.100 191.400 819.900 195.000 ;
        RECT 821.700 191.400 823.500 195.000 ;
        RECT 824.700 191.400 826.500 194.400 ;
        RECT 731.700 185.700 738.000 186.600 ;
        RECT 735.900 183.600 738.000 185.700 ;
        RECT 731.400 181.050 733.200 182.850 ;
        RECT 736.200 181.800 738.000 183.600 ;
        RECT 738.900 184.800 741.900 186.900 ;
        RECT 743.100 186.300 745.200 187.500 ;
        RECT 773.100 186.300 774.300 188.400 ;
        RECT 770.700 185.400 774.300 186.300 ;
        RECT 563.100 178.950 565.200 181.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 691.950 178.950 694.050 181.050 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 731.100 180.300 733.200 181.050 ;
        RECT 731.100 178.950 738.000 180.300 ;
        RECT 544.050 172.500 546.900 173.700 ;
        RECT 549.000 172.500 552.900 173.700 ;
        RECT 555.000 172.500 558.900 173.700 ;
        RECT 561.000 172.500 564.900 173.700 ;
        RECT 490.200 159.000 492.000 165.600 ;
        RECT 493.200 159.600 495.000 165.600 ;
        RECT 496.200 162.600 498.300 164.700 ;
        RECT 499.200 162.600 501.300 164.700 ;
        RECT 502.200 162.600 504.300 164.700 ;
        RECT 496.200 159.600 498.000 162.600 ;
        RECT 499.200 159.600 501.000 162.600 ;
        RECT 502.200 159.600 504.000 162.600 ;
        RECT 505.200 159.000 507.000 165.600 ;
        RECT 508.200 159.600 510.000 165.600 ;
        RECT 511.200 159.000 513.000 165.600 ;
        RECT 514.200 159.600 516.000 165.600 ;
        RECT 517.200 159.000 519.000 165.600 ;
        RECT 520.500 159.600 522.300 165.600 ;
        RECT 523.500 159.000 525.300 165.600 ;
        RECT 542.100 159.000 543.900 171.600 ;
        RECT 545.100 159.600 546.900 172.500 ;
        RECT 548.100 159.000 549.900 171.600 ;
        RECT 551.100 159.600 552.900 172.500 ;
        RECT 554.100 159.000 555.900 171.600 ;
        RECT 557.100 159.600 558.900 172.500 ;
        RECT 560.100 159.000 561.900 171.600 ;
        RECT 563.100 159.600 564.900 172.500 ;
        RECT 566.100 159.000 567.900 171.600 ;
        RECT 585.000 166.800 585.900 178.950 ;
        RECT 590.100 177.150 591.900 178.950 ;
        RECT 611.250 177.150 613.050 178.950 ;
        RECT 614.400 171.600 615.300 178.950 ;
        RECT 617.100 177.150 618.900 178.950 ;
        RECT 585.000 165.900 591.600 166.800 ;
        RECT 585.000 165.600 585.900 165.900 ;
        RECT 584.100 159.600 585.900 165.600 ;
        RECT 590.100 165.600 591.600 165.900 ;
        RECT 587.100 159.000 588.900 165.000 ;
        RECT 590.100 159.600 591.900 165.600 ;
        RECT 593.100 159.000 594.900 165.600 ;
        RECT 611.100 159.000 612.900 171.600 ;
        RECT 614.400 170.400 618.000 171.600 ;
        RECT 616.200 159.600 618.000 170.400 ;
        RECT 636.000 166.800 636.900 178.950 ;
        RECT 641.100 177.150 642.900 178.950 ;
        RECT 665.100 171.600 666.300 178.950 ;
        RECT 636.000 165.900 642.600 166.800 ;
        RECT 636.000 165.600 636.900 165.900 ;
        RECT 635.100 159.600 636.900 165.600 ;
        RECT 641.100 165.600 642.600 165.900 ;
        RECT 638.100 159.000 639.900 165.000 ;
        RECT 641.100 159.600 642.900 165.600 ;
        RECT 644.100 159.000 645.900 165.600 ;
        RECT 662.100 159.000 663.900 171.600 ;
        RECT 665.100 159.600 666.900 171.600 ;
        RECT 684.000 166.800 684.900 178.950 ;
        RECT 689.100 177.150 690.900 178.950 ;
        RECT 684.000 165.900 690.600 166.800 ;
        RECT 684.000 165.600 684.900 165.900 ;
        RECT 683.100 159.600 684.900 165.600 ;
        RECT 689.100 165.600 690.600 165.900 ;
        RECT 710.700 165.600 711.900 178.950 ;
        RECT 713.100 177.150 714.900 178.950 ;
        RECT 736.200 178.500 738.000 178.950 ;
        RECT 738.900 179.100 740.100 184.800 ;
        RECT 741.000 181.800 743.100 183.900 ;
        RECT 741.300 180.000 743.100 181.800 ;
        RECT 767.100 181.050 768.900 182.850 ;
        RECT 770.700 181.050 771.900 185.400 ;
        RECT 773.100 181.050 774.900 182.850 ;
        RECT 791.700 181.050 792.900 191.400 ;
        RECT 815.400 181.050 816.300 191.400 ;
        RECT 738.900 178.200 741.300 179.100 ;
        RECT 739.800 178.050 741.300 178.200 ;
        RECT 745.800 178.950 747.900 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 769.950 178.950 772.050 181.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 735.000 175.500 738.900 177.300 ;
        RECT 736.800 175.200 738.900 175.500 ;
        RECT 739.800 175.950 741.900 178.050 ;
        RECT 745.800 177.150 747.600 178.950 ;
        RECT 764.100 177.150 765.900 178.950 ;
        RECT 739.800 174.000 740.700 175.950 ;
        RECT 733.500 171.600 735.600 173.700 ;
        RECT 739.200 172.950 740.700 174.000 ;
        RECT 739.200 171.600 740.400 172.950 ;
        RECT 731.100 170.700 735.600 171.600 ;
        RECT 686.100 159.000 687.900 165.000 ;
        RECT 689.100 159.600 690.900 165.600 ;
        RECT 692.100 159.000 693.900 165.600 ;
        RECT 710.100 159.600 711.900 165.600 ;
        RECT 713.100 159.000 714.900 165.600 ;
        RECT 731.100 159.600 732.900 170.700 ;
        RECT 734.100 159.000 735.900 169.500 ;
        RECT 738.600 159.600 740.400 171.600 ;
        RECT 743.100 171.600 745.200 172.500 ;
        RECT 770.700 171.600 771.900 178.950 ;
        RECT 743.100 170.400 747.900 171.600 ;
        RECT 743.100 159.000 744.900 169.500 ;
        RECT 746.100 159.600 747.900 170.400 ;
        RECT 764.400 159.000 766.200 171.600 ;
        RECT 769.500 170.100 771.900 171.600 ;
        RECT 769.500 159.600 771.300 170.100 ;
        RECT 772.200 167.100 774.000 168.900 ;
        RECT 791.700 165.600 792.900 178.950 ;
        RECT 794.100 177.150 795.900 178.950 ;
        RECT 812.250 177.150 814.050 178.950 ;
        RECT 815.400 171.600 816.300 178.950 ;
        RECT 818.100 177.150 819.900 178.950 ;
        RECT 825.000 178.050 826.500 191.400 ;
        RECT 824.100 175.950 826.500 178.050 ;
        RECT 772.500 159.000 774.300 165.600 ;
        RECT 791.100 159.600 792.900 165.600 ;
        RECT 794.100 159.000 795.900 165.600 ;
        RECT 812.100 159.000 813.900 171.600 ;
        RECT 815.400 170.400 819.000 171.600 ;
        RECT 817.200 159.600 819.000 170.400 ;
        RECT 825.000 165.600 826.500 175.950 ;
        RECT 828.300 188.400 830.100 194.400 ;
        RECT 833.700 188.400 835.500 195.000 ;
        RECT 838.800 189.600 840.600 194.400 ;
        RECT 843.000 191.400 844.800 194.400 ;
        RECT 846.000 191.400 847.800 194.400 ;
        RECT 849.000 191.400 850.800 194.400 ;
        RECT 852.000 191.400 853.800 194.400 ;
        RECT 855.000 191.400 856.800 195.000 ;
        RECT 836.400 188.400 840.600 189.600 ;
        RECT 842.700 189.300 844.800 191.400 ;
        RECT 845.700 189.300 847.800 191.400 ;
        RECT 848.700 189.300 850.800 191.400 ;
        RECT 851.700 189.300 853.800 191.400 ;
        RECT 858.000 190.500 859.800 194.400 ;
        RECT 862.500 191.400 864.300 195.000 ;
        RECT 865.500 191.400 867.300 194.400 ;
        RECT 868.500 191.400 870.300 194.400 ;
        RECT 871.500 191.400 873.300 194.400 ;
        RECT 857.100 188.400 859.800 190.500 ;
        RECT 861.600 189.600 863.400 190.500 ;
        RECT 861.600 188.400 864.300 189.600 ;
        RECT 865.200 189.300 867.300 191.400 ;
        RECT 868.200 189.300 870.300 191.400 ;
        RECT 871.200 189.300 873.300 191.400 ;
        RECT 875.700 188.400 877.500 194.400 ;
        RECT 881.100 188.400 882.900 195.000 ;
        RECT 886.500 188.400 888.300 194.400 ;
        RECT 828.300 171.600 829.200 188.400 ;
        RECT 836.400 185.100 837.900 188.400 ;
        RECT 842.100 186.600 848.700 188.400 ;
        RECT 863.400 187.800 864.300 188.400 ;
        RECT 866.400 187.800 868.200 188.400 ;
        RECT 863.400 186.600 870.600 187.800 ;
        RECT 830.100 183.300 837.900 185.100 ;
        RECT 854.100 184.500 855.900 186.300 ;
        RECT 853.800 183.900 855.900 184.500 ;
        RECT 838.800 182.400 855.900 183.900 ;
        RECT 860.100 183.900 862.200 184.050 ;
        RECT 863.400 183.900 865.200 184.800 ;
        RECT 860.100 183.000 865.200 183.900 ;
        RECT 869.700 183.600 870.600 186.600 ;
        RECT 875.700 187.500 877.200 188.400 ;
        RECT 875.700 186.300 884.100 187.500 ;
        RECT 882.300 185.700 884.100 186.300 ;
        RECT 871.500 184.800 873.600 185.700 ;
        RECT 887.100 184.800 888.300 188.400 ;
        RECT 905.100 190.200 906.900 193.200 ;
        RECT 908.100 192.600 909.300 195.000 ;
        RECT 917.100 193.200 918.300 195.000 ;
        RECT 905.100 186.900 906.000 190.200 ;
        RECT 908.100 187.800 909.900 192.600 ;
        RECT 912.600 188.700 914.400 193.200 ;
        RECT 912.600 187.800 914.700 188.700 ;
        RECT 905.100 186.000 912.300 186.900 ;
        RECT 871.500 183.600 888.300 184.800 ;
        RECT 833.700 180.900 840.300 182.400 ;
        RECT 860.100 181.950 862.200 183.000 ;
        RECT 868.800 181.800 870.600 183.600 ;
        RECT 833.700 178.050 835.200 180.900 ;
        RECT 841.500 179.700 885.900 180.900 ;
        RECT 841.500 178.200 842.400 179.700 ;
        RECT 833.100 175.950 835.200 178.050 ;
        RECT 837.300 176.400 842.400 178.200 ;
        RECT 845.100 177.900 858.600 178.800 ;
        RECT 865.800 177.900 867.600 178.500 ;
        RECT 884.100 178.050 885.900 179.700 ;
        RECT 845.100 176.700 846.000 177.900 ;
        RECT 845.100 174.900 846.900 176.700 ;
        RECT 851.100 175.200 855.000 177.000 ;
        RECT 856.500 176.700 867.600 177.900 ;
        RECT 878.100 177.750 880.200 178.050 ;
        RECT 856.500 175.800 858.600 176.700 ;
        RECT 876.300 175.950 880.200 177.750 ;
        RECT 884.100 175.950 886.200 178.050 ;
        RECT 876.300 175.200 878.100 175.950 ;
        RECT 851.100 174.900 853.200 175.200 ;
        RECT 864.600 174.300 878.100 175.200 ;
        RECT 830.100 173.700 831.900 174.300 ;
        RECT 864.600 173.700 865.800 174.300 ;
        RECT 830.100 172.500 865.800 173.700 ;
        RECT 868.500 172.500 870.600 172.800 ;
        RECT 828.300 170.700 844.800 171.600 ;
        RECT 828.300 167.400 829.200 170.700 ;
        RECT 833.100 168.600 838.800 169.800 ;
        RECT 842.700 169.500 844.800 170.700 ;
        RECT 848.100 170.400 865.800 171.600 ;
        RECT 868.500 171.300 880.500 172.500 ;
        RECT 868.500 170.700 870.600 171.300 ;
        RECT 878.700 170.700 880.500 171.300 ;
        RECT 848.100 169.500 850.200 170.400 ;
        RECT 864.600 169.800 865.800 170.400 ;
        RECT 882.000 169.800 883.800 170.100 ;
        RECT 833.100 168.000 834.900 168.600 ;
        RECT 828.300 166.500 832.200 167.400 ;
        RECT 831.000 165.600 832.200 166.500 ;
        RECT 837.600 165.600 838.800 168.600 ;
        RECT 839.700 167.700 841.500 168.300 ;
        RECT 839.700 166.500 847.800 167.700 ;
        RECT 845.700 165.600 847.800 166.500 ;
        RECT 851.100 165.600 853.800 169.500 ;
        RECT 856.500 167.100 859.800 169.200 ;
        RECT 864.600 168.600 883.800 169.800 ;
        RECT 821.700 159.000 823.500 165.600 ;
        RECT 824.700 159.600 826.500 165.600 ;
        RECT 828.000 159.000 829.800 165.600 ;
        RECT 831.000 159.600 832.800 165.600 ;
        RECT 834.000 159.000 835.800 165.600 ;
        RECT 837.000 159.600 838.800 165.600 ;
        RECT 840.000 159.000 841.800 165.600 ;
        RECT 842.700 162.600 844.800 164.700 ;
        RECT 845.700 162.600 847.800 164.700 ;
        RECT 848.700 162.600 850.800 164.700 ;
        RECT 843.000 159.600 844.800 162.600 ;
        RECT 846.000 159.600 847.800 162.600 ;
        RECT 849.000 159.600 850.800 162.600 ;
        RECT 852.000 159.600 853.800 165.600 ;
        RECT 855.000 159.000 856.800 165.600 ;
        RECT 858.000 159.600 859.800 167.100 ;
        RECT 865.200 165.600 867.300 167.700 ;
        RECT 861.900 159.000 863.700 165.600 ;
        RECT 864.900 159.600 866.700 165.600 ;
        RECT 867.600 162.600 869.700 164.700 ;
        RECT 870.600 162.600 872.700 164.700 ;
        RECT 867.900 159.600 869.700 162.600 ;
        RECT 870.900 159.600 872.700 162.600 ;
        RECT 874.500 159.000 876.300 165.600 ;
        RECT 877.500 159.600 879.300 168.600 ;
        RECT 882.000 168.300 883.800 168.600 ;
        RECT 887.100 167.400 888.300 183.600 ;
        RECT 905.100 181.050 906.900 182.850 ;
        RECT 905.100 178.950 907.200 181.050 ;
        RECT 908.100 178.950 910.200 181.050 ;
        RECT 911.100 178.950 912.300 186.000 ;
        RECT 913.800 181.050 914.700 187.800 ;
        RECT 917.100 187.200 918.900 193.200 ;
        RECT 935.100 188.400 936.900 194.400 ;
        RECT 938.100 189.300 939.900 195.000 ;
        RECT 942.600 188.400 944.400 194.400 ;
        RECT 947.100 189.300 948.900 195.000 ;
        RECT 950.100 188.400 951.900 194.400 ;
        RECT 968.100 191.400 969.900 195.000 ;
        RECT 971.100 191.400 972.900 194.400 ;
        RECT 974.100 191.400 975.900 195.000 ;
        RECT 992.100 191.400 993.900 194.400 ;
        RECT 995.100 191.400 996.900 195.000 ;
        RECT 935.100 187.500 939.900 188.400 ;
        RECT 937.800 186.300 939.900 187.500 ;
        RECT 942.900 186.900 944.100 188.400 ;
        RECT 941.100 184.800 944.100 186.900 ;
        RECT 950.100 186.600 951.300 188.400 ;
        RECT 939.900 181.800 942.000 183.900 ;
        RECT 913.800 178.950 915.900 181.050 ;
        RECT 916.800 178.950 918.900 181.050 ;
        RECT 935.100 178.950 937.200 181.050 ;
        RECT 939.900 180.000 941.700 181.800 ;
        RECT 942.900 179.100 944.100 184.800 ;
        RECT 945.000 185.700 951.300 186.600 ;
        RECT 945.000 183.600 947.100 185.700 ;
        RECT 945.000 181.800 946.800 183.600 ;
        RECT 949.800 181.050 951.600 182.850 ;
        RECT 971.400 181.050 972.300 191.400 ;
        RECT 992.700 181.050 993.900 191.400 ;
        RECT 1014.000 188.400 1015.800 195.000 ;
        RECT 1018.500 189.600 1020.300 194.400 ;
        RECT 1021.500 191.400 1023.300 195.000 ;
        RECT 1018.500 188.400 1023.600 189.600 ;
        RECT 994.950 186.450 997.050 187.050 ;
        RECT 1003.950 186.450 1006.050 187.050 ;
        RECT 994.950 185.550 1006.050 186.450 ;
        RECT 994.950 184.950 997.050 185.550 ;
        RECT 1003.950 184.950 1006.050 185.550 ;
        RECT 1013.100 181.050 1014.900 182.850 ;
        RECT 1019.250 181.050 1021.050 182.850 ;
        RECT 1022.700 181.050 1023.600 188.400 ;
        RECT 949.800 180.300 951.900 181.050 ;
        RECT 892.950 177.450 895.050 178.050 ;
        RECT 901.950 177.450 904.050 178.050 ;
        RECT 892.950 176.550 904.050 177.450 ;
        RECT 908.100 177.150 909.900 178.950 ;
        RECT 911.100 177.150 912.900 178.950 ;
        RECT 892.950 175.950 895.050 176.550 ;
        RECT 901.950 175.950 904.050 176.550 ;
        RECT 911.700 172.800 912.900 177.150 ;
        RECT 884.700 166.500 888.300 167.400 ;
        RECT 905.100 171.900 912.900 172.800 ;
        RECT 905.100 166.800 906.000 171.900 ;
        RECT 913.800 171.000 914.700 178.950 ;
        RECT 916.800 177.150 918.600 178.950 ;
        RECT 935.400 177.150 937.200 178.950 ;
        RECT 941.700 178.200 944.100 179.100 ;
        RECT 945.000 178.950 951.900 180.300 ;
        RECT 967.950 178.950 970.050 181.050 ;
        RECT 970.950 178.950 973.050 181.050 ;
        RECT 973.950 178.950 976.050 181.050 ;
        RECT 991.950 178.950 994.050 181.050 ;
        RECT 994.950 178.950 997.050 181.050 ;
        RECT 1012.950 178.950 1015.050 181.050 ;
        RECT 1015.950 178.950 1018.050 181.050 ;
        RECT 1018.950 178.950 1021.050 181.050 ;
        RECT 1021.950 178.950 1024.050 181.050 ;
        RECT 945.000 178.500 946.800 178.950 ;
        RECT 941.700 178.050 943.200 178.200 ;
        RECT 941.100 175.950 943.200 178.050 ;
        RECT 942.300 174.000 943.200 175.950 ;
        RECT 944.100 175.500 948.000 177.300 ;
        RECT 968.250 177.150 970.050 178.950 ;
        RECT 944.100 175.200 946.200 175.500 ;
        RECT 942.300 172.950 943.800 174.000 ;
        RECT 937.800 171.600 939.900 172.500 ;
        RECT 884.700 165.600 885.600 166.500 ;
        RECT 880.500 159.000 882.300 165.600 ;
        RECT 883.500 164.700 885.600 165.600 ;
        RECT 883.500 159.600 885.300 164.700 ;
        RECT 886.500 159.000 888.300 165.600 ;
        RECT 905.100 160.800 906.900 166.800 ;
        RECT 908.100 159.000 909.900 171.000 ;
        RECT 912.600 170.100 914.700 171.000 ;
        RECT 912.600 159.600 914.400 170.100 ;
        RECT 917.100 159.000 918.900 171.600 ;
        RECT 935.100 170.400 939.900 171.600 ;
        RECT 942.600 171.600 943.800 172.950 ;
        RECT 947.400 171.600 949.500 173.700 ;
        RECT 971.400 171.600 972.300 178.950 ;
        RECT 974.100 177.150 975.900 178.950 ;
        RECT 935.100 159.600 936.900 170.400 ;
        RECT 938.100 159.000 939.900 169.500 ;
        RECT 942.600 159.600 944.400 171.600 ;
        RECT 947.400 170.700 951.900 171.600 ;
        RECT 947.100 159.000 948.900 169.500 ;
        RECT 950.100 159.600 951.900 170.700 ;
        RECT 968.100 159.000 969.900 171.600 ;
        RECT 971.400 170.400 975.000 171.600 ;
        RECT 973.200 159.600 975.000 170.400 ;
        RECT 992.700 165.600 993.900 178.950 ;
        RECT 995.100 177.150 996.900 178.950 ;
        RECT 1016.250 177.150 1018.050 178.950 ;
        RECT 1022.700 171.600 1023.600 178.950 ;
        RECT 1013.100 170.700 1020.900 171.600 ;
        RECT 992.100 159.600 993.900 165.600 ;
        RECT 995.100 159.000 996.900 165.600 ;
        RECT 1013.100 159.600 1014.900 170.700 ;
        RECT 1016.100 159.000 1017.900 169.800 ;
        RECT 1019.100 159.600 1020.900 170.700 ;
        RECT 1022.100 159.600 1023.900 171.600 ;
        RECT 17.100 143.400 18.900 156.000 ;
        RECT 21.600 143.400 24.900 155.400 ;
        RECT 27.600 143.400 29.400 156.000 ;
        RECT 47.100 149.400 48.900 156.000 ;
        RECT 50.100 149.400 51.900 155.400 ;
        RECT 53.100 149.400 54.900 156.000 ;
        RECT 71.700 149.400 73.500 156.000 ;
        RECT 17.100 136.050 18.900 137.850 ;
        RECT 22.950 136.050 24.000 143.400 ;
        RECT 25.950 141.450 28.050 142.050 ;
        RECT 46.950 141.450 49.050 142.050 ;
        RECT 25.950 140.550 49.050 141.450 ;
        RECT 25.950 139.950 28.050 140.550 ;
        RECT 46.950 139.950 49.050 140.550 ;
        RECT 28.950 136.050 30.750 137.850 ;
        RECT 50.700 136.050 51.900 149.400 ;
        RECT 72.000 146.100 73.800 147.900 ;
        RECT 74.700 144.900 76.500 155.400 ;
        RECT 74.100 143.400 76.500 144.900 ;
        RECT 79.800 143.400 81.600 156.000 ;
        RECT 98.100 149.400 99.900 156.000 ;
        RECT 101.100 149.400 102.900 155.400 ;
        RECT 104.100 149.400 105.900 156.000 ;
        RECT 74.100 136.050 75.300 143.400 ;
        RECT 80.100 136.050 81.900 137.850 ;
        RECT 101.700 136.050 102.900 149.400 ;
        RECT 122.100 143.400 123.900 155.400 ;
        RECT 125.100 144.000 126.900 156.000 ;
        RECT 128.100 149.400 129.900 155.400 ;
        RECT 131.100 149.400 132.900 156.000 ;
        RECT 106.950 138.450 109.050 139.050 ;
        RECT 115.950 138.450 118.050 139.050 ;
        RECT 106.950 137.550 118.050 138.450 ;
        RECT 106.950 136.950 109.050 137.550 ;
        RECT 115.950 136.950 118.050 137.550 ;
        RECT 122.700 136.050 123.600 143.400 ;
        RECT 126.000 136.050 127.800 137.850 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 20.250 132.150 22.050 133.950 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 28.950 133.950 31.050 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 122.100 133.950 124.200 136.050 ;
        RECT 125.400 133.950 127.500 136.050 ;
        RECT 22.950 129.300 24.000 133.950 ;
        RECT 25.950 132.150 27.750 133.950 ;
        RECT 47.100 132.150 48.900 133.950 ;
        RECT 22.950 128.100 27.300 129.300 ;
        RECT 50.700 128.700 51.900 133.950 ;
        RECT 52.950 132.150 54.750 133.950 ;
        RECT 71.100 132.150 72.900 133.950 ;
        RECT 74.100 129.600 75.300 133.950 ;
        RECT 77.100 132.150 78.900 133.950 ;
        RECT 98.100 132.150 99.900 133.950 ;
        RECT 17.100 126.000 24.900 126.900 ;
        RECT 26.400 126.600 27.300 128.100 ;
        RECT 47.700 127.800 51.900 128.700 ;
        RECT 71.700 128.700 75.300 129.600 ;
        RECT 101.700 128.700 102.900 133.950 ;
        RECT 103.950 132.150 105.750 133.950 ;
        RECT 17.100 120.600 18.900 126.000 ;
        RECT 20.100 120.000 21.900 125.100 ;
        RECT 23.100 121.500 24.900 126.000 ;
        RECT 26.100 122.400 27.900 126.600 ;
        RECT 29.100 121.500 30.900 126.600 ;
        RECT 23.100 120.600 30.900 121.500 ;
        RECT 47.700 120.600 49.500 127.800 ;
        RECT 71.700 126.600 72.900 128.700 ;
        RECT 98.700 127.800 102.900 128.700 ;
        RECT 52.800 120.000 54.600 126.600 ;
        RECT 71.100 120.600 72.900 126.600 ;
        RECT 74.100 125.700 81.900 127.050 ;
        RECT 74.100 120.600 75.900 125.700 ;
        RECT 77.100 120.000 78.900 124.800 ;
        RECT 80.100 120.600 81.900 125.700 ;
        RECT 98.700 120.600 100.500 127.800 ;
        RECT 122.700 126.600 123.600 133.950 ;
        RECT 129.000 129.300 129.900 149.400 ;
        RECT 149.100 144.600 150.900 155.400 ;
        RECT 152.100 145.500 153.900 156.000 ;
        RECT 149.100 143.400 153.900 144.600 ;
        RECT 151.800 142.500 153.900 143.400 ;
        RECT 156.600 143.400 158.400 155.400 ;
        RECT 161.100 145.500 162.900 156.000 ;
        RECT 164.100 144.300 165.900 155.400 ;
        RECT 182.700 149.400 184.500 156.000 ;
        RECT 183.000 146.100 184.800 147.900 ;
        RECT 185.700 144.900 187.500 155.400 ;
        RECT 161.400 143.400 165.900 144.300 ;
        RECT 185.100 143.400 187.500 144.900 ;
        RECT 190.800 143.400 192.600 156.000 ;
        RECT 210.000 144.600 211.800 155.400 ;
        RECT 210.000 143.400 213.600 144.600 ;
        RECT 215.100 143.400 216.900 156.000 ;
        RECT 233.100 143.400 234.900 156.000 ;
        RECT 238.200 144.600 240.000 155.400 ;
        RECT 257.100 149.400 258.900 156.000 ;
        RECT 260.100 149.400 261.900 155.400 ;
        RECT 263.100 150.000 264.900 156.000 ;
        RECT 260.400 149.100 261.900 149.400 ;
        RECT 266.100 149.400 267.900 155.400 ;
        RECT 284.100 149.400 285.900 156.000 ;
        RECT 287.100 149.400 288.900 155.400 ;
        RECT 290.100 149.400 291.900 156.000 ;
        RECT 266.100 149.100 267.000 149.400 ;
        RECT 260.400 148.200 267.000 149.100 ;
        RECT 236.400 143.400 240.000 144.600 ;
        RECT 156.600 142.050 157.800 143.400 ;
        RECT 156.300 141.000 157.800 142.050 ;
        RECT 161.400 141.300 163.500 143.400 ;
        RECT 156.300 139.050 157.200 141.000 ;
        RECT 149.400 136.050 151.200 137.850 ;
        RECT 155.100 136.950 157.200 139.050 ;
        RECT 158.100 139.500 160.200 139.800 ;
        RECT 158.100 137.700 162.000 139.500 ;
        RECT 130.800 133.950 132.900 136.050 ;
        RECT 149.100 133.950 151.200 136.050 ;
        RECT 155.700 136.800 157.200 136.950 ;
        RECT 155.700 135.900 158.100 136.800 ;
        RECT 130.950 132.150 132.750 133.950 ;
        RECT 153.900 133.200 155.700 135.000 ;
        RECT 153.900 131.100 156.000 133.200 ;
        RECT 156.900 130.200 158.100 135.900 ;
        RECT 159.000 136.050 160.800 136.500 ;
        RECT 185.100 136.050 186.300 143.400 ;
        RECT 191.100 136.050 192.900 137.850 ;
        RECT 209.100 136.050 210.900 137.850 ;
        RECT 212.700 136.050 213.600 143.400 ;
        RECT 214.950 136.050 216.750 137.850 ;
        RECT 233.250 136.050 235.050 137.850 ;
        RECT 236.400 136.050 237.300 143.400 ;
        RECT 239.100 136.050 240.900 137.850 ;
        RECT 260.100 136.050 261.900 137.850 ;
        RECT 266.100 136.050 267.000 148.200 ;
        RECT 287.100 136.050 288.300 149.400 ;
        RECT 308.100 143.400 309.900 156.000 ;
        RECT 313.200 144.600 315.000 155.400 ;
        RECT 311.400 143.400 315.000 144.600 ;
        RECT 332.400 143.400 334.200 156.000 ;
        RECT 337.500 144.900 339.300 155.400 ;
        RECT 340.500 149.400 342.300 156.000 ;
        RECT 340.200 146.100 342.000 147.900 ;
        RECT 337.500 143.400 339.900 144.900 ;
        RECT 359.100 143.400 360.900 155.400 ;
        RECT 362.100 143.400 363.900 156.000 ;
        RECT 380.100 143.400 381.900 155.400 ;
        RECT 383.100 145.200 384.900 156.000 ;
        RECT 386.100 149.400 387.900 155.400 ;
        RECT 308.250 136.050 310.050 137.850 ;
        RECT 311.400 136.050 312.300 143.400 ;
        RECT 314.100 136.050 315.900 137.850 ;
        RECT 332.100 136.050 333.900 137.850 ;
        RECT 338.700 136.050 339.900 143.400 ;
        RECT 359.700 136.050 360.900 143.400 ;
        RECT 380.100 136.050 381.300 143.400 ;
        RECT 386.700 142.500 387.900 149.400 ;
        RECT 404.100 143.400 405.900 156.000 ;
        RECT 409.200 144.600 411.000 155.400 ;
        RECT 428.100 149.400 429.900 155.400 ;
        RECT 431.100 149.400 432.900 156.000 ;
        RECT 407.400 143.400 411.000 144.600 ;
        RECT 382.200 141.600 387.900 142.500 ;
        RECT 382.200 140.700 384.000 141.600 ;
        RECT 159.000 134.700 165.900 136.050 ;
        RECT 163.800 133.950 165.900 134.700 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 184.950 133.950 187.050 136.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 190.950 133.950 193.050 136.050 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 232.950 133.950 235.050 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 380.100 133.950 382.200 136.050 ;
        RECT 124.500 128.400 132.900 129.300 ;
        RECT 124.500 127.500 126.300 128.400 ;
        RECT 103.800 120.000 105.600 126.600 ;
        RECT 122.700 124.800 125.400 126.600 ;
        RECT 123.600 120.600 125.400 124.800 ;
        RECT 126.600 120.000 128.400 126.600 ;
        RECT 131.100 120.600 132.900 128.400 ;
        RECT 151.800 127.500 153.900 128.700 ;
        RECT 155.100 128.100 158.100 130.200 ;
        RECT 159.000 131.400 160.800 133.200 ;
        RECT 163.800 132.150 165.600 133.950 ;
        RECT 182.100 132.150 183.900 133.950 ;
        RECT 159.000 129.300 161.100 131.400 ;
        RECT 185.100 129.600 186.300 133.950 ;
        RECT 188.100 132.150 189.900 133.950 ;
        RECT 159.000 128.400 165.300 129.300 ;
        RECT 149.100 126.600 153.900 127.500 ;
        RECT 156.900 126.600 158.100 128.100 ;
        RECT 164.100 126.600 165.300 128.400 ;
        RECT 182.700 128.700 186.300 129.600 ;
        RECT 182.700 126.600 183.900 128.700 ;
        RECT 149.100 120.600 150.900 126.600 ;
        RECT 152.100 120.000 153.900 125.700 ;
        RECT 156.600 120.600 158.400 126.600 ;
        RECT 161.100 120.000 162.900 125.700 ;
        RECT 164.100 120.600 165.900 126.600 ;
        RECT 182.100 120.600 183.900 126.600 ;
        RECT 185.100 125.700 192.900 127.050 ;
        RECT 185.100 120.600 186.900 125.700 ;
        RECT 188.100 120.000 189.900 124.800 ;
        RECT 191.100 120.600 192.900 125.700 ;
        RECT 202.950 126.450 205.050 127.050 ;
        RECT 208.950 126.450 211.050 127.050 ;
        RECT 202.950 125.550 211.050 126.450 ;
        RECT 202.950 124.950 205.050 125.550 ;
        RECT 208.950 124.950 211.050 125.550 ;
        RECT 212.700 123.600 213.600 133.950 ;
        RECT 236.400 123.600 237.300 133.950 ;
        RECT 257.100 132.150 258.900 133.950 ;
        RECT 263.100 132.150 264.900 133.950 ;
        RECT 266.100 130.200 267.000 133.950 ;
        RECT 284.250 132.150 286.050 133.950 ;
        RECT 238.950 129.450 241.050 130.050 ;
        RECT 250.950 129.450 253.050 130.050 ;
        RECT 238.950 128.550 253.050 129.450 ;
        RECT 238.950 127.950 241.050 128.550 ;
        RECT 250.950 127.950 253.050 128.550 ;
        RECT 209.100 120.000 210.900 123.600 ;
        RECT 212.100 120.600 213.900 123.600 ;
        RECT 215.100 120.000 216.900 123.600 ;
        RECT 233.100 120.000 234.900 123.600 ;
        RECT 236.100 120.600 237.900 123.600 ;
        RECT 239.100 120.000 240.900 123.600 ;
        RECT 257.100 120.000 258.900 129.600 ;
        RECT 263.700 129.000 267.000 130.200 ;
        RECT 263.700 120.600 265.500 129.000 ;
        RECT 287.100 128.700 288.300 133.950 ;
        RECT 290.100 132.150 291.900 133.950 ;
        RECT 287.100 127.800 291.300 128.700 ;
        RECT 284.400 120.000 286.200 126.600 ;
        RECT 289.500 120.600 291.300 127.800 ;
        RECT 311.400 123.600 312.300 133.950 ;
        RECT 335.100 132.150 336.900 133.950 ;
        RECT 338.700 129.600 339.900 133.950 ;
        RECT 341.100 132.150 342.900 133.950 ;
        RECT 338.700 128.700 342.300 129.600 ;
        RECT 332.100 125.700 339.900 127.050 ;
        RECT 308.100 120.000 309.900 123.600 ;
        RECT 311.100 120.600 312.900 123.600 ;
        RECT 314.100 120.000 315.900 123.600 ;
        RECT 332.100 120.600 333.900 125.700 ;
        RECT 335.100 120.000 336.900 124.800 ;
        RECT 338.100 120.600 339.900 125.700 ;
        RECT 341.100 126.600 342.300 128.700 ;
        RECT 359.700 126.600 360.900 133.950 ;
        RECT 362.100 132.150 363.900 133.950 ;
        RECT 380.100 126.600 381.300 133.950 ;
        RECT 383.100 129.300 384.000 140.700 ;
        RECT 385.800 136.050 387.600 137.850 ;
        RECT 404.250 136.050 406.050 137.850 ;
        RECT 407.400 136.050 408.300 143.400 ;
        RECT 410.100 136.050 411.900 137.850 ;
        RECT 428.700 136.050 429.900 149.400 ;
        RECT 449.100 143.400 450.900 156.000 ;
        RECT 454.200 144.600 456.000 155.400 ;
        RECT 452.400 143.400 456.000 144.600 ;
        RECT 470.100 143.400 471.900 155.400 ;
        RECT 473.100 144.300 474.900 155.400 ;
        RECT 476.100 145.200 477.900 156.000 ;
        RECT 479.100 144.300 480.900 155.400 ;
        RECT 473.100 143.400 480.900 144.300 ;
        RECT 497.100 144.600 498.900 155.400 ;
        RECT 500.100 145.500 502.200 156.000 ;
        RECT 497.100 143.400 502.200 144.600 ;
        RECT 504.600 144.300 506.400 155.400 ;
        RECT 509.100 145.500 510.900 156.000 ;
        RECT 512.100 144.300 513.900 155.400 ;
        RECT 431.100 136.050 432.900 137.850 ;
        RECT 449.250 136.050 451.050 137.850 ;
        RECT 452.400 136.050 453.300 143.400 ;
        RECT 455.100 136.050 456.900 137.850 ;
        RECT 470.400 136.050 471.300 143.400 ;
        RECT 500.100 142.500 502.200 143.400 ;
        RECT 503.100 143.400 506.400 144.300 ;
        RECT 503.100 139.050 504.300 143.400 ;
        RECT 509.100 143.100 513.900 144.300 ;
        RECT 530.400 143.400 532.200 156.000 ;
        RECT 535.500 144.900 537.300 155.400 ;
        RECT 538.500 149.400 540.300 156.000 ;
        RECT 538.200 146.100 540.000 147.900 ;
        RECT 535.500 143.400 537.900 144.900 ;
        RECT 557.100 144.300 558.900 155.400 ;
        RECT 560.100 145.500 561.900 156.000 ;
        RECT 557.100 143.400 561.600 144.300 ;
        RECT 564.600 143.400 566.400 155.400 ;
        RECT 569.100 145.500 570.900 156.000 ;
        RECT 572.100 144.600 573.900 155.400 ;
        RECT 590.100 149.400 591.900 156.000 ;
        RECT 593.100 149.400 594.900 155.400 ;
        RECT 611.100 149.400 612.900 155.400 ;
        RECT 614.100 150.000 615.900 156.000 ;
        RECT 509.100 142.200 511.200 143.100 ;
        RECT 505.800 141.300 511.200 142.200 ;
        RECT 514.950 141.450 517.050 142.050 ;
        RECT 520.950 141.450 523.050 142.050 ;
        RECT 505.800 139.500 507.600 141.300 ;
        RECT 514.950 140.550 523.050 141.450 ;
        RECT 514.950 139.950 517.050 140.550 ;
        RECT 520.950 139.950 523.050 140.550 ;
        RECT 502.800 138.300 504.900 139.050 ;
        RECT 475.950 136.050 477.750 137.850 ;
        RECT 497.400 136.050 499.200 137.850 ;
        RECT 502.800 136.950 505.800 138.300 ;
        RECT 385.500 133.950 387.600 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 406.950 133.950 409.050 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 497.100 133.950 499.200 136.050 ;
        RECT 502.200 134.100 504.000 135.900 ;
        RECT 382.200 128.400 384.000 129.300 ;
        RECT 382.200 127.500 387.900 128.400 ;
        RECT 341.100 120.600 342.900 126.600 ;
        RECT 359.100 120.600 360.900 126.600 ;
        RECT 362.100 120.000 363.900 126.600 ;
        RECT 380.100 120.600 381.900 126.600 ;
        RECT 383.100 120.000 384.900 126.600 ;
        RECT 386.700 123.600 387.900 127.500 ;
        RECT 388.950 126.450 391.050 127.050 ;
        RECT 397.950 126.450 400.050 127.050 ;
        RECT 388.950 125.550 400.050 126.450 ;
        RECT 388.950 124.950 391.050 125.550 ;
        RECT 397.950 124.950 400.050 125.550 ;
        RECT 407.400 123.600 408.300 133.950 ;
        RECT 428.700 123.600 429.900 133.950 ;
        RECT 452.400 123.600 453.300 133.950 ;
        RECT 470.400 126.600 471.300 133.950 ;
        RECT 472.950 132.150 474.750 133.950 ;
        RECT 479.100 132.150 480.900 133.950 ;
        RECT 501.900 132.000 504.000 134.100 ;
        RECT 504.900 130.200 505.800 136.950 ;
        RECT 507.300 136.200 509.100 138.000 ;
        RECT 507.000 134.100 509.100 136.200 ;
        RECT 530.100 136.050 531.900 137.850 ;
        RECT 536.700 136.050 537.900 143.400 ;
        RECT 559.500 141.300 561.600 143.400 ;
        RECT 565.200 142.050 566.400 143.400 ;
        RECT 569.100 143.400 573.900 144.600 ;
        RECT 569.100 142.500 571.200 143.400 ;
        RECT 565.200 141.000 566.700 142.050 ;
        RECT 562.800 139.500 564.900 139.800 ;
        RECT 561.000 137.700 564.900 139.500 ;
        RECT 565.800 139.050 566.700 141.000 ;
        RECT 565.800 136.950 567.900 139.050 ;
        RECT 565.800 136.800 567.300 136.950 ;
        RECT 562.200 136.050 564.000 136.500 ;
        RECT 511.800 133.800 513.900 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 557.100 134.700 564.000 136.050 ;
        RECT 564.900 135.900 567.300 136.800 ;
        RECT 571.800 136.050 573.600 137.850 ;
        RECT 590.100 136.050 591.900 137.850 ;
        RECT 593.100 136.050 594.300 149.400 ;
        RECT 612.000 149.100 612.900 149.400 ;
        RECT 617.100 149.400 618.900 155.400 ;
        RECT 620.100 149.400 621.900 156.000 ;
        RECT 617.100 149.100 618.600 149.400 ;
        RECT 612.000 148.200 618.600 149.100 ;
        RECT 612.000 136.050 612.900 148.200 ;
        RECT 628.950 147.450 631.050 148.050 ;
        RECT 634.950 147.450 637.050 148.050 ;
        RECT 628.950 146.550 637.050 147.450 ;
        RECT 628.950 145.950 631.050 146.550 ;
        RECT 634.950 145.950 637.050 146.550 ;
        RECT 638.100 144.300 639.900 155.400 ;
        RECT 641.100 145.500 642.900 156.000 ;
        RECT 638.100 143.400 642.600 144.300 ;
        RECT 645.600 143.400 647.400 155.400 ;
        RECT 650.100 145.500 651.900 156.000 ;
        RECT 653.100 144.600 654.900 155.400 ;
        RECT 671.100 149.400 672.900 156.000 ;
        RECT 674.100 149.400 675.900 155.400 ;
        RECT 677.100 149.400 678.900 156.000 ;
        RECT 640.500 141.300 642.600 143.400 ;
        RECT 646.200 142.050 647.400 143.400 ;
        RECT 650.100 143.400 654.900 144.600 ;
        RECT 664.950 144.450 667.050 145.050 ;
        RECT 670.950 144.450 673.050 145.050 ;
        RECT 664.950 143.550 673.050 144.450 ;
        RECT 650.100 142.500 652.200 143.400 ;
        RECT 664.950 142.950 667.050 143.550 ;
        RECT 670.950 142.950 673.050 143.550 ;
        RECT 646.200 141.000 647.700 142.050 ;
        RECT 643.800 139.500 645.900 139.800 ;
        RECT 617.100 136.050 618.900 137.850 ;
        RECT 642.000 137.700 645.900 139.500 ;
        RECT 646.800 139.050 647.700 141.000 ;
        RECT 646.800 136.950 648.900 139.050 ;
        RECT 646.800 136.800 648.300 136.950 ;
        RECT 643.200 136.050 645.000 136.500 ;
        RECT 557.100 133.950 559.200 134.700 ;
        RECT 511.800 133.200 513.600 133.800 ;
        RECT 507.000 132.000 513.600 133.200 ;
        RECT 533.100 132.150 534.900 133.950 ;
        RECT 507.000 131.100 509.100 132.000 ;
        RECT 499.500 127.500 501.600 129.900 ;
        RECT 502.800 128.100 505.800 130.200 ;
        RECT 506.700 129.300 508.500 131.100 ;
        RECT 536.700 129.600 537.900 133.950 ;
        RECT 539.100 132.150 540.900 133.950 ;
        RECT 557.400 132.150 559.200 133.950 ;
        RECT 562.200 131.400 564.000 133.200 ;
        RECT 497.100 126.600 501.600 127.500 ;
        RECT 470.400 125.400 475.500 126.600 ;
        RECT 386.100 120.600 387.900 123.600 ;
        RECT 404.100 120.000 405.900 123.600 ;
        RECT 407.100 120.600 408.900 123.600 ;
        RECT 410.100 120.000 411.900 123.600 ;
        RECT 428.100 120.600 429.900 123.600 ;
        RECT 431.100 120.000 432.900 123.600 ;
        RECT 449.100 120.000 450.900 123.600 ;
        RECT 452.100 120.600 453.900 123.600 ;
        RECT 455.100 120.000 456.900 123.600 ;
        RECT 470.700 120.000 472.500 123.600 ;
        RECT 473.700 120.600 475.500 125.400 ;
        RECT 478.200 120.000 480.000 126.600 ;
        RECT 497.100 120.600 498.900 126.600 ;
        RECT 504.900 126.000 505.800 128.100 ;
        RECT 509.400 129.000 511.500 129.600 ;
        RECT 509.400 127.500 513.900 129.000 ;
        RECT 536.700 128.700 540.300 129.600 ;
        RECT 561.900 129.300 564.000 131.400 ;
        RECT 512.400 126.600 513.900 127.500 ;
        RECT 500.400 120.000 502.200 125.700 ;
        RECT 504.900 120.600 506.700 126.000 ;
        RECT 509.100 120.000 510.900 125.700 ;
        RECT 512.100 120.600 513.900 126.600 ;
        RECT 530.100 125.700 537.900 127.050 ;
        RECT 530.100 120.600 531.900 125.700 ;
        RECT 533.100 120.000 534.900 124.800 ;
        RECT 536.100 120.600 537.900 125.700 ;
        RECT 539.100 126.600 540.300 128.700 ;
        RECT 557.700 128.400 564.000 129.300 ;
        RECT 564.900 130.200 566.100 135.900 ;
        RECT 567.300 133.200 569.100 135.000 ;
        RECT 571.800 133.950 573.900 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 638.100 134.700 645.000 136.050 ;
        RECT 645.900 135.900 648.300 136.800 ;
        RECT 652.800 136.050 654.600 137.850 ;
        RECT 674.100 136.050 675.300 149.400 ;
        RECT 676.950 144.450 679.050 145.050 ;
        RECT 688.950 144.450 691.050 145.050 ;
        RECT 676.950 143.550 691.050 144.450 ;
        RECT 676.950 142.950 679.050 143.550 ;
        RECT 688.950 142.950 691.050 143.550 ;
        RECT 695.100 144.600 696.900 155.400 ;
        RECT 698.100 145.500 700.200 156.000 ;
        RECT 695.100 143.400 700.200 144.600 ;
        RECT 702.600 144.300 704.400 155.400 ;
        RECT 707.100 145.500 708.900 156.000 ;
        RECT 710.100 144.300 711.900 155.400 ;
        RECT 698.100 142.500 700.200 143.400 ;
        RECT 701.100 143.400 704.400 144.300 ;
        RECT 679.950 141.450 682.050 142.050 ;
        RECT 691.950 141.450 694.050 142.050 ;
        RECT 679.950 140.550 694.050 141.450 ;
        RECT 679.950 139.950 682.050 140.550 ;
        RECT 691.950 139.950 694.050 140.550 ;
        RECT 701.100 139.050 702.300 143.400 ;
        RECT 707.100 143.100 711.900 144.300 ;
        RECT 728.400 143.400 730.200 156.000 ;
        RECT 733.500 144.900 735.300 155.400 ;
        RECT 736.500 149.400 738.300 156.000 ;
        RECT 736.200 146.100 738.000 147.900 ;
        RECT 733.500 143.400 735.900 144.900 ;
        RECT 755.100 143.400 756.900 156.000 ;
        RECT 707.100 142.200 709.200 143.100 ;
        RECT 703.800 141.300 709.200 142.200 ;
        RECT 703.800 139.500 705.600 141.300 ;
        RECT 700.800 138.300 702.900 139.050 ;
        RECT 695.400 136.050 697.200 137.850 ;
        RECT 700.800 136.950 703.800 138.300 ;
        RECT 638.100 133.950 640.200 134.700 ;
        RECT 567.000 131.100 569.100 133.200 ;
        RECT 557.700 126.600 558.900 128.400 ;
        RECT 564.900 128.100 567.900 130.200 ;
        RECT 574.950 129.450 577.050 130.050 ;
        RECT 583.950 129.450 586.050 130.050 ;
        RECT 589.950 129.450 592.050 130.050 ;
        RECT 564.900 126.600 566.100 128.100 ;
        RECT 569.100 127.500 571.200 128.700 ;
        RECT 574.950 128.550 592.050 129.450 ;
        RECT 574.950 127.950 577.050 128.550 ;
        RECT 583.950 127.950 586.050 128.550 ;
        RECT 589.950 127.950 592.050 128.550 ;
        RECT 569.100 126.600 573.900 127.500 ;
        RECT 539.100 120.600 540.900 126.600 ;
        RECT 557.100 120.600 558.900 126.600 ;
        RECT 560.100 120.000 561.900 125.700 ;
        RECT 564.600 120.600 566.400 126.600 ;
        RECT 569.100 120.000 570.900 125.700 ;
        RECT 572.100 120.600 573.900 126.600 ;
        RECT 593.100 123.600 594.300 133.950 ;
        RECT 612.000 130.200 612.900 133.950 ;
        RECT 614.100 132.150 615.900 133.950 ;
        RECT 620.100 132.150 621.900 133.950 ;
        RECT 638.400 132.150 640.200 133.950 ;
        RECT 643.200 131.400 645.000 133.200 ;
        RECT 612.000 129.000 615.300 130.200 ;
        RECT 590.100 120.000 591.900 123.600 ;
        RECT 593.100 120.600 594.900 123.600 ;
        RECT 613.500 120.600 615.300 129.000 ;
        RECT 620.100 120.000 621.900 129.600 ;
        RECT 642.900 129.300 645.000 131.400 ;
        RECT 638.700 128.400 645.000 129.300 ;
        RECT 645.900 130.200 647.100 135.900 ;
        RECT 648.300 133.200 650.100 135.000 ;
        RECT 652.800 133.950 654.900 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 695.100 133.950 697.200 136.050 ;
        RECT 700.200 134.100 702.000 135.900 ;
        RECT 648.000 131.100 650.100 133.200 ;
        RECT 671.250 132.150 673.050 133.950 ;
        RECT 638.700 126.600 639.900 128.400 ;
        RECT 645.900 128.100 648.900 130.200 ;
        RECT 658.950 129.450 661.050 130.050 ;
        RECT 670.950 129.450 673.050 130.050 ;
        RECT 645.900 126.600 647.100 128.100 ;
        RECT 650.100 127.500 652.200 128.700 ;
        RECT 658.950 128.550 673.050 129.450 ;
        RECT 658.950 127.950 661.050 128.550 ;
        RECT 670.950 127.950 673.050 128.550 ;
        RECT 674.100 128.700 675.300 133.950 ;
        RECT 677.100 132.150 678.900 133.950 ;
        RECT 699.900 132.000 702.000 134.100 ;
        RECT 702.900 130.200 703.800 136.950 ;
        RECT 705.300 136.200 707.100 138.000 ;
        RECT 705.000 134.100 707.100 136.200 ;
        RECT 728.100 136.050 729.900 137.850 ;
        RECT 734.700 136.050 735.900 143.400 ;
        RECT 758.100 142.500 759.900 155.400 ;
        RECT 761.100 143.400 762.900 156.000 ;
        RECT 764.100 142.500 765.900 155.400 ;
        RECT 767.100 143.400 768.900 156.000 ;
        RECT 770.100 142.500 771.900 155.400 ;
        RECT 773.100 143.400 774.900 156.000 ;
        RECT 776.100 142.500 777.900 155.400 ;
        RECT 779.100 143.400 780.900 156.000 ;
        RECT 797.100 149.400 798.900 156.000 ;
        RECT 800.100 149.400 801.900 155.400 ;
        RECT 803.100 149.400 804.900 156.000 ;
        RECT 821.700 149.400 823.500 156.000 ;
        RECT 758.100 141.300 762.000 142.500 ;
        RECT 764.100 141.300 768.000 142.500 ;
        RECT 770.100 141.300 774.000 142.500 ;
        RECT 776.100 141.300 778.950 142.500 ;
        RECT 709.800 133.800 711.900 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 757.800 133.950 759.900 136.050 ;
        RECT 709.800 133.200 711.600 133.800 ;
        RECT 705.000 132.000 711.600 133.200 ;
        RECT 731.100 132.150 732.900 133.950 ;
        RECT 705.000 131.100 707.100 132.000 ;
        RECT 674.100 127.800 678.300 128.700 ;
        RECT 650.100 126.600 654.900 127.500 ;
        RECT 638.100 120.600 639.900 126.600 ;
        RECT 641.100 120.000 642.900 125.700 ;
        RECT 645.600 120.600 647.400 126.600 ;
        RECT 650.100 120.000 651.900 125.700 ;
        RECT 653.100 120.600 654.900 126.600 ;
        RECT 671.400 120.000 673.200 126.600 ;
        RECT 676.500 120.600 678.300 127.800 ;
        RECT 697.500 127.500 699.600 129.900 ;
        RECT 700.800 128.100 703.800 130.200 ;
        RECT 704.700 129.300 706.500 131.100 ;
        RECT 734.700 129.600 735.900 133.950 ;
        RECT 737.100 132.150 738.900 133.950 ;
        RECT 757.800 132.150 759.600 133.950 ;
        RECT 760.800 130.800 762.000 141.300 ;
        RECT 763.200 130.800 765.000 131.400 ;
        RECT 760.800 129.600 765.000 130.800 ;
        RECT 766.800 130.800 768.000 141.300 ;
        RECT 769.200 130.800 771.000 131.400 ;
        RECT 766.800 129.600 771.000 130.800 ;
        RECT 772.800 130.800 774.000 141.300 ;
        RECT 777.900 136.050 778.950 141.300 ;
        RECT 800.100 136.050 801.300 149.400 ;
        RECT 822.000 146.100 823.800 147.900 ;
        RECT 824.700 144.900 826.500 155.400 ;
        RECT 824.100 143.400 826.500 144.900 ;
        RECT 829.800 143.400 831.600 156.000 ;
        RECT 848.100 144.600 849.900 155.400 ;
        RECT 851.100 145.500 852.900 156.000 ;
        RECT 848.100 143.400 852.900 144.600 ;
        RECT 824.100 136.050 825.300 143.400 ;
        RECT 850.800 142.500 852.900 143.400 ;
        RECT 855.600 143.400 857.400 155.400 ;
        RECT 860.100 145.500 861.900 156.000 ;
        RECT 863.100 144.300 864.900 155.400 ;
        RECT 881.100 149.400 882.900 156.000 ;
        RECT 884.100 149.400 885.900 155.400 ;
        RECT 887.100 149.400 888.900 156.000 ;
        RECT 905.100 149.400 906.900 156.000 ;
        RECT 908.100 149.400 909.900 155.400 ;
        RECT 860.400 143.400 864.900 144.300 ;
        RECT 855.600 142.050 856.800 143.400 ;
        RECT 826.950 141.450 829.050 142.050 ;
        RECT 838.950 141.450 841.050 142.050 ;
        RECT 826.950 140.550 841.050 141.450 ;
        RECT 826.950 139.950 829.050 140.550 ;
        RECT 838.950 139.950 841.050 140.550 ;
        RECT 855.300 141.000 856.800 142.050 ;
        RECT 860.400 141.300 862.500 143.400 ;
        RECT 855.300 139.050 856.200 141.000 ;
        RECT 830.100 136.050 831.900 137.850 ;
        RECT 848.400 136.050 850.200 137.850 ;
        RECT 854.100 136.950 856.200 139.050 ;
        RECT 857.100 139.500 859.200 139.800 ;
        RECT 857.100 137.700 861.000 139.500 ;
        RECT 775.800 133.950 778.950 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 826.950 133.950 829.050 136.050 ;
        RECT 829.950 133.950 832.050 136.050 ;
        RECT 848.100 133.950 850.200 136.050 ;
        RECT 854.700 136.800 856.200 136.950 ;
        RECT 854.700 135.900 857.100 136.800 ;
        RECT 775.200 130.800 777.000 131.400 ;
        RECT 772.800 129.600 777.000 130.800 ;
        RECT 695.100 126.600 699.600 127.500 ;
        RECT 695.100 120.600 696.900 126.600 ;
        RECT 702.900 126.000 703.800 128.100 ;
        RECT 707.400 129.000 709.500 129.600 ;
        RECT 707.400 127.500 711.900 129.000 ;
        RECT 734.700 128.700 738.300 129.600 ;
        RECT 760.800 128.700 762.000 129.600 ;
        RECT 766.800 128.700 768.000 129.600 ;
        RECT 772.800 128.700 774.000 129.600 ;
        RECT 777.900 128.700 778.950 133.950 ;
        RECT 797.250 132.150 799.050 133.950 ;
        RECT 710.400 126.600 711.900 127.500 ;
        RECT 698.400 120.000 700.200 125.700 ;
        RECT 702.900 120.600 704.700 126.000 ;
        RECT 707.100 120.000 708.900 125.700 ;
        RECT 710.100 120.600 711.900 126.600 ;
        RECT 728.100 125.700 735.900 127.050 ;
        RECT 728.100 120.600 729.900 125.700 ;
        RECT 731.100 120.000 732.900 124.800 ;
        RECT 734.100 120.600 735.900 125.700 ;
        RECT 737.100 126.600 738.300 128.700 ;
        RECT 758.100 127.500 762.000 128.700 ;
        RECT 764.100 127.500 768.000 128.700 ;
        RECT 770.100 127.500 774.000 128.700 ;
        RECT 776.100 127.500 778.950 128.700 ;
        RECT 800.100 128.700 801.300 133.950 ;
        RECT 803.100 132.150 804.900 133.950 ;
        RECT 821.100 132.150 822.900 133.950 ;
        RECT 824.100 129.600 825.300 133.950 ;
        RECT 827.100 132.150 828.900 133.950 ;
        RECT 852.900 133.200 854.700 135.000 ;
        RECT 852.900 131.100 855.000 133.200 ;
        RECT 855.900 130.200 857.100 135.900 ;
        RECT 858.000 136.050 859.800 136.500 ;
        RECT 884.100 136.050 885.300 149.400 ;
        RECT 905.100 136.050 906.900 137.850 ;
        RECT 908.100 136.050 909.300 149.400 ;
        RECT 926.100 144.600 927.900 155.400 ;
        RECT 929.100 145.500 930.900 156.000 ;
        RECT 926.100 143.400 930.900 144.600 ;
        RECT 928.800 142.500 930.900 143.400 ;
        RECT 933.600 143.400 935.400 155.400 ;
        RECT 938.100 145.500 939.900 156.000 ;
        RECT 941.100 144.300 942.900 155.400 ;
        RECT 938.400 143.400 942.900 144.300 ;
        RECT 943.950 144.450 946.050 145.050 ;
        RECT 952.950 144.450 955.050 145.050 ;
        RECT 943.950 143.550 955.050 144.450 ;
        RECT 933.600 142.050 934.800 143.400 ;
        RECT 933.300 141.000 934.800 142.050 ;
        RECT 938.400 141.300 940.500 143.400 ;
        RECT 943.950 142.950 946.050 143.550 ;
        RECT 952.950 142.950 955.050 143.550 ;
        RECT 959.100 143.400 960.900 155.400 ;
        RECT 962.100 143.400 963.900 156.000 ;
        RECT 980.100 144.600 981.900 155.400 ;
        RECT 983.100 145.500 984.900 156.000 ;
        RECT 980.100 143.400 984.900 144.600 ;
        RECT 933.300 139.050 934.200 141.000 ;
        RECT 926.400 136.050 928.200 137.850 ;
        RECT 932.100 136.950 934.200 139.050 ;
        RECT 935.100 139.500 937.200 139.800 ;
        RECT 935.100 137.700 939.000 139.500 ;
        RECT 943.950 138.450 946.050 139.050 ;
        RECT 955.950 138.450 958.050 139.050 ;
        RECT 943.950 137.550 958.050 138.450 ;
        RECT 943.950 136.950 946.050 137.550 ;
        RECT 955.950 136.950 958.050 137.550 ;
        RECT 858.000 134.700 864.900 136.050 ;
        RECT 862.800 133.950 864.900 134.700 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 926.100 133.950 928.200 136.050 ;
        RECT 932.700 136.800 934.200 136.950 ;
        RECT 932.700 135.900 935.100 136.800 ;
        RECT 821.700 128.700 825.300 129.600 ;
        RECT 800.100 127.800 804.300 128.700 ;
        RECT 737.100 120.600 738.900 126.600 ;
        RECT 755.100 120.000 756.900 126.600 ;
        RECT 758.100 120.600 759.900 127.500 ;
        RECT 761.100 120.000 762.900 126.600 ;
        RECT 764.100 120.600 765.900 127.500 ;
        RECT 767.100 120.000 768.900 126.600 ;
        RECT 770.100 120.600 771.900 127.500 ;
        RECT 773.100 120.000 774.900 126.600 ;
        RECT 776.100 120.600 777.900 127.500 ;
        RECT 779.100 120.000 780.900 126.600 ;
        RECT 797.400 120.000 799.200 126.600 ;
        RECT 802.500 120.600 804.300 127.800 ;
        RECT 821.700 126.600 822.900 128.700 ;
        RECT 850.800 127.500 852.900 128.700 ;
        RECT 854.100 128.100 857.100 130.200 ;
        RECT 858.000 131.400 859.800 133.200 ;
        RECT 862.800 132.150 864.600 133.950 ;
        RECT 881.250 132.150 883.050 133.950 ;
        RECT 858.000 129.300 860.100 131.400 ;
        RECT 858.000 128.400 864.300 129.300 ;
        RECT 821.100 120.600 822.900 126.600 ;
        RECT 824.100 125.700 831.900 127.050 ;
        RECT 824.100 120.600 825.900 125.700 ;
        RECT 827.100 120.000 828.900 124.800 ;
        RECT 830.100 120.600 831.900 125.700 ;
        RECT 848.100 126.600 852.900 127.500 ;
        RECT 855.900 126.600 857.100 128.100 ;
        RECT 863.100 126.600 864.300 128.400 ;
        RECT 884.100 128.700 885.300 133.950 ;
        RECT 887.100 132.150 888.900 133.950 ;
        RECT 884.100 127.800 888.300 128.700 ;
        RECT 848.100 120.600 849.900 126.600 ;
        RECT 851.100 120.000 852.900 125.700 ;
        RECT 855.600 120.600 857.400 126.600 ;
        RECT 860.100 120.000 861.900 125.700 ;
        RECT 863.100 120.600 864.900 126.600 ;
        RECT 881.400 120.000 883.200 126.600 ;
        RECT 886.500 120.600 888.300 127.800 ;
        RECT 908.100 123.600 909.300 133.950 ;
        RECT 930.900 133.200 932.700 135.000 ;
        RECT 930.900 131.100 933.000 133.200 ;
        RECT 933.900 130.200 935.100 135.900 ;
        RECT 936.000 136.050 937.800 136.500 ;
        RECT 959.700 136.050 960.900 143.400 ;
        RECT 982.800 142.500 984.900 143.400 ;
        RECT 987.600 143.400 989.400 155.400 ;
        RECT 992.100 145.500 993.900 156.000 ;
        RECT 995.100 144.300 996.900 155.400 ;
        RECT 1013.700 149.400 1015.500 156.000 ;
        RECT 1014.000 146.100 1015.800 147.900 ;
        RECT 1016.700 144.900 1018.500 155.400 ;
        RECT 992.400 143.400 996.900 144.300 ;
        RECT 1016.100 143.400 1018.500 144.900 ;
        RECT 1021.800 143.400 1023.600 156.000 ;
        RECT 987.600 142.050 988.800 143.400 ;
        RECT 987.300 141.000 988.800 142.050 ;
        RECT 992.400 141.300 994.500 143.400 ;
        RECT 987.300 139.050 988.200 141.000 ;
        RECT 980.400 136.050 982.200 137.850 ;
        RECT 986.100 136.950 988.200 139.050 ;
        RECT 989.100 139.500 991.200 139.800 ;
        RECT 989.100 137.700 993.000 139.500 ;
        RECT 936.000 134.700 942.900 136.050 ;
        RECT 940.800 133.950 942.900 134.700 ;
        RECT 958.950 133.950 961.050 136.050 ;
        RECT 961.950 133.950 964.050 136.050 ;
        RECT 980.100 133.950 982.200 136.050 ;
        RECT 986.700 136.800 988.200 136.950 ;
        RECT 986.700 135.900 989.100 136.800 ;
        RECT 928.800 127.500 930.900 128.700 ;
        RECT 932.100 128.100 935.100 130.200 ;
        RECT 936.000 131.400 937.800 133.200 ;
        RECT 940.800 132.150 942.600 133.950 ;
        RECT 936.000 129.300 938.100 131.400 ;
        RECT 936.000 128.400 942.300 129.300 ;
        RECT 926.100 126.600 930.900 127.500 ;
        RECT 933.900 126.600 935.100 128.100 ;
        RECT 941.100 126.600 942.300 128.400 ;
        RECT 959.700 126.600 960.900 133.950 ;
        RECT 962.100 132.150 963.900 133.950 ;
        RECT 984.900 133.200 986.700 135.000 ;
        RECT 984.900 131.100 987.000 133.200 ;
        RECT 987.900 130.200 989.100 135.900 ;
        RECT 990.000 136.050 991.800 136.500 ;
        RECT 1016.100 136.050 1017.300 143.400 ;
        RECT 1022.100 136.050 1023.900 137.850 ;
        RECT 990.000 134.700 996.900 136.050 ;
        RECT 994.800 133.950 996.900 134.700 ;
        RECT 1012.950 133.950 1015.050 136.050 ;
        RECT 1015.950 133.950 1018.050 136.050 ;
        RECT 1018.950 133.950 1021.050 136.050 ;
        RECT 1021.950 133.950 1024.050 136.050 ;
        RECT 982.800 127.500 984.900 128.700 ;
        RECT 986.100 128.100 989.100 130.200 ;
        RECT 990.000 131.400 991.800 133.200 ;
        RECT 994.800 132.150 996.600 133.950 ;
        RECT 1013.100 132.150 1014.900 133.950 ;
        RECT 990.000 129.300 992.100 131.400 ;
        RECT 1016.100 129.600 1017.300 133.950 ;
        RECT 1019.100 132.150 1020.900 133.950 ;
        RECT 990.000 128.400 996.300 129.300 ;
        RECT 980.100 126.600 984.900 127.500 ;
        RECT 987.900 126.600 989.100 128.100 ;
        RECT 995.100 126.600 996.300 128.400 ;
        RECT 1013.700 128.700 1017.300 129.600 ;
        RECT 1013.700 126.600 1014.900 128.700 ;
        RECT 905.100 120.000 906.900 123.600 ;
        RECT 908.100 120.600 909.900 123.600 ;
        RECT 926.100 120.600 927.900 126.600 ;
        RECT 929.100 120.000 930.900 125.700 ;
        RECT 933.600 120.600 935.400 126.600 ;
        RECT 938.100 120.000 939.900 125.700 ;
        RECT 941.100 120.600 942.900 126.600 ;
        RECT 959.100 120.600 960.900 126.600 ;
        RECT 962.100 120.000 963.900 126.600 ;
        RECT 980.100 120.600 981.900 126.600 ;
        RECT 983.100 120.000 984.900 125.700 ;
        RECT 987.600 120.600 989.400 126.600 ;
        RECT 992.100 120.000 993.900 125.700 ;
        RECT 995.100 120.600 996.900 126.600 ;
        RECT 1013.100 120.600 1014.900 126.600 ;
        RECT 1016.100 125.700 1023.900 127.050 ;
        RECT 1016.100 120.600 1017.900 125.700 ;
        RECT 1019.100 120.000 1020.900 124.800 ;
        RECT 1022.100 120.600 1023.900 125.700 ;
        RECT 17.100 113.400 18.900 117.000 ;
        RECT 20.100 113.400 21.900 116.400 ;
        RECT 23.100 113.400 24.900 117.000 ;
        RECT 20.700 103.050 21.600 113.400 ;
        RECT 41.100 110.400 42.900 116.400 ;
        RECT 41.700 108.300 42.900 110.400 ;
        RECT 44.100 111.300 45.900 116.400 ;
        RECT 47.100 112.200 48.900 117.000 ;
        RECT 50.100 111.300 51.900 116.400 ;
        RECT 68.100 113.400 69.900 117.000 ;
        RECT 71.100 113.400 72.900 116.400 ;
        RECT 74.100 113.400 75.900 117.000 ;
        RECT 44.100 109.950 51.900 111.300 ;
        RECT 41.700 107.400 45.300 108.300 ;
        RECT 41.100 103.050 42.900 104.850 ;
        RECT 44.100 103.050 45.300 107.400 ;
        RECT 47.100 103.050 48.900 104.850 ;
        RECT 71.400 103.050 72.300 113.400 ;
        RECT 93.000 110.400 94.800 117.000 ;
        RECT 97.500 111.600 99.300 116.400 ;
        RECT 100.500 113.400 102.300 117.000 ;
        RECT 97.500 110.400 102.600 111.600 ;
        RECT 119.100 110.400 120.900 116.400 ;
        RECT 122.100 111.300 123.900 117.000 ;
        RECT 126.600 110.400 128.400 116.400 ;
        RECT 131.100 111.300 132.900 117.000 ;
        RECT 134.100 110.400 135.900 116.400 ;
        RECT 92.100 103.050 93.900 104.850 ;
        RECT 98.250 103.050 100.050 104.850 ;
        RECT 101.700 103.050 102.600 110.400 ;
        RECT 119.700 108.600 120.900 110.400 ;
        RECT 126.900 108.900 128.100 110.400 ;
        RECT 131.100 109.500 135.900 110.400 ;
        RECT 152.100 110.400 153.900 116.400 ;
        RECT 155.100 111.300 156.900 117.000 ;
        RECT 159.600 110.400 161.400 116.400 ;
        RECT 164.100 111.300 165.900 117.000 ;
        RECT 167.100 110.400 168.900 116.400 ;
        RECT 152.100 109.500 156.900 110.400 ;
        RECT 119.700 107.700 126.000 108.600 ;
        RECT 123.900 105.600 126.000 107.700 ;
        RECT 119.400 103.050 121.200 104.850 ;
        RECT 124.200 103.800 126.000 105.600 ;
        RECT 126.900 106.800 129.900 108.900 ;
        RECT 131.100 108.300 133.200 109.500 ;
        RECT 154.800 108.300 156.900 109.500 ;
        RECT 159.900 108.900 161.100 110.400 ;
        RECT 158.100 106.800 161.100 108.900 ;
        RECT 167.100 108.600 168.300 110.400 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 119.100 102.300 121.200 103.050 ;
        RECT 119.100 100.950 126.000 102.300 ;
        RECT 17.100 99.150 18.900 100.950 ;
        RECT 20.700 93.600 21.600 100.950 ;
        RECT 22.950 99.150 24.750 100.950 ;
        RECT 44.100 93.600 45.300 100.950 ;
        RECT 50.100 99.150 51.900 100.950 ;
        RECT 68.250 99.150 70.050 100.950 ;
        RECT 71.400 93.600 72.300 100.950 ;
        RECT 74.100 99.150 75.900 100.950 ;
        RECT 95.250 99.150 97.050 100.950 ;
        RECT 82.950 96.450 85.050 97.050 ;
        RECT 97.950 96.450 100.050 97.050 ;
        RECT 82.950 95.550 100.050 96.450 ;
        RECT 82.950 94.950 85.050 95.550 ;
        RECT 97.950 94.950 100.050 95.550 ;
        RECT 101.700 93.600 102.600 100.950 ;
        RECT 124.200 100.500 126.000 100.950 ;
        RECT 126.900 101.100 128.100 106.800 ;
        RECT 129.000 103.800 131.100 105.900 ;
        RECT 129.300 102.000 131.100 103.800 ;
        RECT 156.900 103.800 159.000 105.900 ;
        RECT 126.900 100.200 129.300 101.100 ;
        RECT 127.800 100.050 129.300 100.200 ;
        RECT 133.800 100.950 135.900 103.050 ;
        RECT 152.100 100.950 154.200 103.050 ;
        RECT 156.900 102.000 158.700 103.800 ;
        RECT 159.900 101.100 161.100 106.800 ;
        RECT 162.000 107.700 168.300 108.600 ;
        RECT 185.700 109.200 187.500 116.400 ;
        RECT 190.800 110.400 192.600 117.000 ;
        RECT 185.700 108.300 189.900 109.200 ;
        RECT 162.000 105.600 164.100 107.700 ;
        RECT 162.000 103.800 163.800 105.600 ;
        RECT 166.800 103.050 168.600 104.850 ;
        RECT 185.100 103.050 186.900 104.850 ;
        RECT 188.700 103.050 189.900 108.300 ;
        RECT 209.100 107.400 210.900 117.000 ;
        RECT 215.700 108.000 217.500 116.400 ;
        RECT 236.700 113.400 238.500 117.000 ;
        RECT 239.700 111.600 241.500 116.400 ;
        RECT 236.400 110.400 241.500 111.600 ;
        RECT 244.200 110.400 246.000 117.000 ;
        RECT 215.700 106.800 219.000 108.000 ;
        RECT 190.950 103.050 192.750 104.850 ;
        RECT 209.100 103.050 210.900 104.850 ;
        RECT 215.100 103.050 216.900 104.850 ;
        RECT 218.100 103.050 219.000 106.800 ;
        RECT 236.400 103.050 237.300 110.400 ;
        RECT 263.100 107.400 264.900 117.000 ;
        RECT 269.700 108.000 271.500 116.400 ;
        RECT 290.100 110.400 291.900 117.000 ;
        RECT 293.100 110.400 294.900 116.400 ;
        RECT 296.700 113.400 298.500 117.000 ;
        RECT 299.700 113.400 301.500 116.400 ;
        RECT 269.700 106.800 273.000 108.000 ;
        RECT 238.950 103.050 240.750 104.850 ;
        RECT 245.100 103.050 246.900 104.850 ;
        RECT 263.100 103.050 264.900 104.850 ;
        RECT 269.100 103.050 270.900 104.850 ;
        RECT 272.100 103.050 273.000 106.800 ;
        RECT 290.100 103.050 291.900 104.850 ;
        RECT 293.100 103.050 294.300 110.400 ;
        RECT 166.800 102.300 168.900 103.050 ;
        RECT 123.000 97.500 126.900 99.300 ;
        RECT 124.800 97.200 126.900 97.500 ;
        RECT 127.800 97.950 129.900 100.050 ;
        RECT 133.800 99.150 135.600 100.950 ;
        RECT 152.400 99.150 154.200 100.950 ;
        RECT 158.700 100.200 161.100 101.100 ;
        RECT 162.000 100.950 168.900 102.300 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 162.000 100.500 163.800 100.950 ;
        RECT 158.700 100.050 160.200 100.200 ;
        RECT 158.100 97.950 160.200 100.050 ;
        RECT 127.800 96.000 128.700 97.950 ;
        RECT 121.500 93.600 123.600 95.700 ;
        RECT 127.200 94.950 128.700 96.000 ;
        RECT 159.300 96.000 160.200 97.950 ;
        RECT 161.100 97.500 165.000 99.300 ;
        RECT 161.100 97.200 163.200 97.500 ;
        RECT 159.300 94.950 160.800 96.000 ;
        RECT 127.200 93.600 128.400 94.950 ;
        RECT 18.000 92.400 21.600 93.600 ;
        RECT 18.000 81.600 19.800 92.400 ;
        RECT 23.100 81.000 24.900 93.600 ;
        RECT 44.100 92.100 46.500 93.600 ;
        RECT 42.000 89.100 43.800 90.900 ;
        RECT 41.700 81.000 43.500 87.600 ;
        RECT 44.700 81.600 46.500 92.100 ;
        RECT 49.800 81.000 51.600 93.600 ;
        RECT 68.100 81.000 69.900 93.600 ;
        RECT 71.400 92.400 75.000 93.600 ;
        RECT 73.200 81.600 75.000 92.400 ;
        RECT 92.100 92.700 99.900 93.600 ;
        RECT 92.100 81.600 93.900 92.700 ;
        RECT 95.100 81.000 96.900 91.800 ;
        RECT 98.100 81.600 99.900 92.700 ;
        RECT 101.100 81.600 102.900 93.600 ;
        RECT 119.100 92.700 123.600 93.600 ;
        RECT 119.100 81.600 120.900 92.700 ;
        RECT 122.100 81.000 123.900 91.500 ;
        RECT 126.600 81.600 128.400 93.600 ;
        RECT 131.100 93.600 133.200 94.500 ;
        RECT 154.800 93.600 156.900 94.500 ;
        RECT 131.100 92.400 135.900 93.600 ;
        RECT 131.100 81.000 132.900 91.500 ;
        RECT 134.100 81.600 135.900 92.400 ;
        RECT 152.100 92.400 156.900 93.600 ;
        RECT 159.600 93.600 160.800 94.950 ;
        RECT 164.400 93.600 166.500 95.700 ;
        RECT 152.100 81.600 153.900 92.400 ;
        RECT 155.100 81.000 156.900 91.500 ;
        RECT 159.600 81.600 161.400 93.600 ;
        RECT 164.400 92.700 168.900 93.600 ;
        RECT 164.100 81.000 165.900 91.500 ;
        RECT 167.100 81.600 168.900 92.700 ;
        RECT 188.700 87.600 189.900 100.950 ;
        RECT 212.100 99.150 213.900 100.950 ;
        RECT 218.100 88.800 219.000 100.950 ;
        RECT 236.400 93.600 237.300 100.950 ;
        RECT 241.950 99.150 243.750 100.950 ;
        RECT 266.100 99.150 267.900 100.950 ;
        RECT 259.950 96.450 262.050 97.050 ;
        RECT 268.950 96.450 271.050 97.050 ;
        RECT 259.950 95.550 271.050 96.450 ;
        RECT 259.950 94.950 262.050 95.550 ;
        RECT 268.950 94.950 271.050 95.550 ;
        RECT 212.400 87.900 219.000 88.800 ;
        RECT 212.400 87.600 213.900 87.900 ;
        RECT 185.100 81.000 186.900 87.600 ;
        RECT 188.100 81.600 189.900 87.600 ;
        RECT 191.100 81.000 192.900 87.600 ;
        RECT 209.100 81.000 210.900 87.600 ;
        RECT 212.100 81.600 213.900 87.600 ;
        RECT 218.100 87.600 219.000 87.900 ;
        RECT 215.100 81.000 216.900 87.000 ;
        RECT 218.100 81.600 219.900 87.600 ;
        RECT 236.100 81.600 237.900 93.600 ;
        RECT 239.100 92.700 246.900 93.600 ;
        RECT 239.100 81.600 240.900 92.700 ;
        RECT 242.100 81.000 243.900 91.800 ;
        RECT 245.100 81.600 246.900 92.700 ;
        RECT 272.100 88.800 273.000 100.950 ;
        RECT 293.100 93.600 294.300 100.950 ;
        RECT 300.000 100.050 301.500 113.400 ;
        RECT 299.100 97.950 301.500 100.050 ;
        RECT 266.400 87.900 273.000 88.800 ;
        RECT 266.400 87.600 267.900 87.900 ;
        RECT 263.100 81.000 264.900 87.600 ;
        RECT 266.100 81.600 267.900 87.600 ;
        RECT 272.100 87.600 273.000 87.900 ;
        RECT 269.100 81.000 270.900 87.000 ;
        RECT 272.100 81.600 273.900 87.600 ;
        RECT 290.100 81.000 291.900 93.600 ;
        RECT 293.100 81.600 294.900 93.600 ;
        RECT 300.000 87.600 301.500 97.950 ;
        RECT 303.300 110.400 305.100 116.400 ;
        RECT 308.700 110.400 310.500 117.000 ;
        RECT 313.800 111.600 315.600 116.400 ;
        RECT 318.000 113.400 319.800 116.400 ;
        RECT 321.000 113.400 322.800 116.400 ;
        RECT 324.000 113.400 325.800 116.400 ;
        RECT 327.000 113.400 328.800 116.400 ;
        RECT 330.000 113.400 331.800 117.000 ;
        RECT 311.400 110.400 315.600 111.600 ;
        RECT 317.700 111.300 319.800 113.400 ;
        RECT 320.700 111.300 322.800 113.400 ;
        RECT 323.700 111.300 325.800 113.400 ;
        RECT 326.700 111.300 328.800 113.400 ;
        RECT 333.000 112.500 334.800 116.400 ;
        RECT 337.500 113.400 339.300 117.000 ;
        RECT 340.500 113.400 342.300 116.400 ;
        RECT 343.500 113.400 345.300 116.400 ;
        RECT 346.500 113.400 348.300 116.400 ;
        RECT 332.100 110.400 334.800 112.500 ;
        RECT 336.600 111.600 338.400 112.500 ;
        RECT 336.600 110.400 339.300 111.600 ;
        RECT 340.200 111.300 342.300 113.400 ;
        RECT 343.200 111.300 345.300 113.400 ;
        RECT 346.200 111.300 348.300 113.400 ;
        RECT 350.700 110.400 352.500 116.400 ;
        RECT 356.100 110.400 357.900 117.000 ;
        RECT 361.500 110.400 363.300 116.400 ;
        RECT 303.300 93.600 304.200 110.400 ;
        RECT 311.400 107.100 312.900 110.400 ;
        RECT 317.100 108.600 323.700 110.400 ;
        RECT 338.400 109.800 339.300 110.400 ;
        RECT 341.400 109.800 343.200 110.400 ;
        RECT 338.400 108.600 345.600 109.800 ;
        RECT 305.100 105.300 312.900 107.100 ;
        RECT 329.100 106.500 330.900 108.300 ;
        RECT 328.800 105.900 330.900 106.500 ;
        RECT 313.800 104.400 330.900 105.900 ;
        RECT 335.100 105.900 337.200 106.050 ;
        RECT 338.400 105.900 340.200 106.800 ;
        RECT 335.100 105.000 340.200 105.900 ;
        RECT 344.700 105.600 345.600 108.600 ;
        RECT 350.700 109.500 352.200 110.400 ;
        RECT 350.700 108.300 359.100 109.500 ;
        RECT 357.300 107.700 359.100 108.300 ;
        RECT 346.500 106.800 348.600 107.700 ;
        RECT 362.100 106.800 363.300 110.400 ;
        RECT 380.100 111.000 381.900 116.400 ;
        RECT 383.100 111.900 384.900 117.000 ;
        RECT 386.100 115.500 393.900 116.400 ;
        RECT 386.100 111.000 387.900 115.500 ;
        RECT 380.100 110.100 387.900 111.000 ;
        RECT 389.100 110.400 390.900 114.600 ;
        RECT 392.100 110.400 393.900 115.500 ;
        RECT 410.100 110.400 411.900 116.400 ;
        RECT 413.100 110.400 414.900 117.000 ;
        RECT 431.100 113.400 432.900 117.000 ;
        RECT 434.100 113.400 435.900 116.400 ;
        RECT 437.100 113.400 438.900 117.000 ;
        RECT 389.400 108.900 390.300 110.400 ;
        RECT 346.500 105.600 363.300 106.800 ;
        RECT 308.700 102.900 315.300 104.400 ;
        RECT 335.100 103.950 337.200 105.000 ;
        RECT 343.800 103.800 345.600 105.600 ;
        RECT 308.700 100.050 310.200 102.900 ;
        RECT 316.500 101.700 360.900 102.900 ;
        RECT 316.500 100.200 317.400 101.700 ;
        RECT 308.100 97.950 310.200 100.050 ;
        RECT 312.300 98.400 317.400 100.200 ;
        RECT 320.100 99.900 333.600 100.800 ;
        RECT 340.800 99.900 342.600 100.500 ;
        RECT 359.100 100.050 360.900 101.700 ;
        RECT 320.100 98.700 321.000 99.900 ;
        RECT 320.100 96.900 321.900 98.700 ;
        RECT 326.100 97.200 330.000 99.000 ;
        RECT 331.500 98.700 342.600 99.900 ;
        RECT 353.100 99.750 355.200 100.050 ;
        RECT 331.500 97.800 333.600 98.700 ;
        RECT 351.300 97.950 355.200 99.750 ;
        RECT 359.100 97.950 361.200 100.050 ;
        RECT 351.300 97.200 353.100 97.950 ;
        RECT 326.100 96.900 328.200 97.200 ;
        RECT 339.600 96.300 353.100 97.200 ;
        RECT 305.100 95.700 306.900 96.300 ;
        RECT 339.600 95.700 340.800 96.300 ;
        RECT 305.100 94.500 340.800 95.700 ;
        RECT 343.500 94.500 345.600 94.800 ;
        RECT 303.300 92.700 319.800 93.600 ;
        RECT 303.300 89.400 304.200 92.700 ;
        RECT 308.100 90.600 313.800 91.800 ;
        RECT 317.700 91.500 319.800 92.700 ;
        RECT 323.100 92.400 340.800 93.600 ;
        RECT 343.500 93.300 355.500 94.500 ;
        RECT 343.500 92.700 345.600 93.300 ;
        RECT 353.700 92.700 355.500 93.300 ;
        RECT 323.100 91.500 325.200 92.400 ;
        RECT 339.600 91.800 340.800 92.400 ;
        RECT 357.000 91.800 358.800 92.100 ;
        RECT 308.100 90.000 309.900 90.600 ;
        RECT 303.300 88.500 307.200 89.400 ;
        RECT 306.000 87.600 307.200 88.500 ;
        RECT 312.600 87.600 313.800 90.600 ;
        RECT 314.700 89.700 316.500 90.300 ;
        RECT 314.700 88.500 322.800 89.700 ;
        RECT 320.700 87.600 322.800 88.500 ;
        RECT 326.100 87.600 328.800 91.500 ;
        RECT 331.500 89.100 334.800 91.200 ;
        RECT 339.600 90.600 358.800 91.800 ;
        RECT 296.700 81.000 298.500 87.600 ;
        RECT 299.700 81.600 301.500 87.600 ;
        RECT 303.000 81.000 304.800 87.600 ;
        RECT 306.000 81.600 307.800 87.600 ;
        RECT 309.000 81.000 310.800 87.600 ;
        RECT 312.000 81.600 313.800 87.600 ;
        RECT 315.000 81.000 316.800 87.600 ;
        RECT 317.700 84.600 319.800 86.700 ;
        RECT 320.700 84.600 322.800 86.700 ;
        RECT 323.700 84.600 325.800 86.700 ;
        RECT 318.000 81.600 319.800 84.600 ;
        RECT 321.000 81.600 322.800 84.600 ;
        RECT 324.000 81.600 325.800 84.600 ;
        RECT 327.000 81.600 328.800 87.600 ;
        RECT 330.000 81.000 331.800 87.600 ;
        RECT 333.000 81.600 334.800 89.100 ;
        RECT 340.200 87.600 342.300 89.700 ;
        RECT 336.900 81.000 338.700 87.600 ;
        RECT 339.900 81.600 341.700 87.600 ;
        RECT 342.600 84.600 344.700 86.700 ;
        RECT 345.600 84.600 347.700 86.700 ;
        RECT 342.900 81.600 344.700 84.600 ;
        RECT 345.900 81.600 347.700 84.600 ;
        RECT 349.500 81.000 351.300 87.600 ;
        RECT 352.500 81.600 354.300 90.600 ;
        RECT 357.000 90.300 358.800 90.600 ;
        RECT 362.100 89.400 363.300 105.600 ;
        RECT 385.950 107.700 390.300 108.900 ;
        RECT 383.250 103.050 385.050 104.850 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 103.050 387.000 107.700 ;
        RECT 388.950 103.050 390.750 104.850 ;
        RECT 410.700 103.050 411.900 110.400 ;
        RECT 413.100 103.050 414.900 104.850 ;
        RECT 434.400 103.050 435.300 113.400 ;
        RECT 455.400 110.400 457.200 117.000 ;
        RECT 460.500 109.200 462.300 116.400 ;
        RECT 479.100 111.000 480.900 116.400 ;
        RECT 482.100 111.900 483.900 117.000 ;
        RECT 485.100 115.500 492.900 116.400 ;
        RECT 485.100 111.000 486.900 115.500 ;
        RECT 479.100 110.100 486.900 111.000 ;
        RECT 488.100 110.400 489.900 114.600 ;
        RECT 491.100 110.400 492.900 115.500 ;
        RECT 458.100 108.300 462.300 109.200 ;
        RECT 488.400 108.900 489.300 110.400 ;
        RECT 455.250 103.050 457.050 104.850 ;
        RECT 458.100 103.050 459.300 108.300 ;
        RECT 484.950 107.700 489.300 108.900 ;
        RECT 511.500 108.000 513.300 116.400 ;
        RECT 461.100 103.050 462.900 104.850 ;
        RECT 482.250 103.050 484.050 104.850 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 103.050 486.000 107.700 ;
        RECT 510.000 106.800 513.300 108.000 ;
        RECT 518.100 107.400 519.900 117.000 ;
        RECT 537.000 110.400 538.800 117.000 ;
        RECT 541.500 111.600 543.300 116.400 ;
        RECT 544.500 113.400 546.300 117.000 ;
        RECT 541.500 110.400 546.600 111.600 ;
        RECT 487.950 103.050 489.750 104.850 ;
        RECT 510.000 103.050 510.900 106.800 ;
        RECT 512.100 103.050 513.900 104.850 ;
        RECT 518.100 103.050 519.900 104.850 ;
        RECT 536.100 103.050 537.900 104.850 ;
        RECT 542.250 103.050 544.050 104.850 ;
        RECT 545.700 103.050 546.600 110.400 ;
        RECT 563.100 107.400 564.900 117.000 ;
        RECT 569.700 108.000 571.500 116.400 ;
        RECT 590.400 110.400 592.200 117.000 ;
        RECT 595.500 109.200 597.300 116.400 ;
        RECT 593.100 108.300 597.300 109.200 ;
        RECT 614.700 109.200 616.500 116.400 ;
        RECT 619.800 110.400 621.600 117.000 ;
        RECT 638.100 110.400 639.900 116.400 ;
        RECT 641.100 111.300 642.900 117.000 ;
        RECT 645.600 110.400 647.400 116.400 ;
        RECT 650.100 111.300 651.900 117.000 ;
        RECT 653.100 110.400 654.900 116.400 ;
        RECT 671.100 110.400 672.900 116.400 ;
        RECT 614.700 108.300 618.900 109.200 ;
        RECT 569.700 106.800 573.000 108.000 ;
        RECT 563.100 103.050 564.900 104.850 ;
        RECT 569.100 103.050 570.900 104.850 ;
        RECT 572.100 103.050 573.000 106.800 ;
        RECT 590.250 103.050 592.050 104.850 ;
        RECT 593.100 103.050 594.300 108.300 ;
        RECT 596.100 103.050 597.900 104.850 ;
        RECT 614.100 103.050 615.900 104.850 ;
        RECT 617.700 103.050 618.900 108.300 ;
        RECT 638.700 108.600 639.900 110.400 ;
        RECT 645.900 108.900 647.100 110.400 ;
        RECT 650.100 109.500 654.900 110.400 ;
        RECT 638.700 107.700 645.000 108.600 ;
        RECT 642.900 105.600 645.000 107.700 ;
        RECT 619.950 103.050 621.750 104.850 ;
        RECT 638.400 103.050 640.200 104.850 ;
        RECT 643.200 103.800 645.000 105.600 ;
        RECT 645.900 106.800 648.900 108.900 ;
        RECT 650.100 108.300 652.200 109.500 ;
        RECT 671.700 108.300 672.900 110.400 ;
        RECT 674.100 111.300 675.900 116.400 ;
        RECT 677.100 112.200 678.900 117.000 ;
        RECT 680.100 111.300 681.900 116.400 ;
        RECT 674.100 109.950 681.900 111.300 ;
        RECT 671.700 107.400 675.300 108.300 ;
        RECT 698.100 107.400 699.900 117.000 ;
        RECT 704.700 108.000 706.500 116.400 ;
        RECT 710.700 113.400 712.500 117.000 ;
        RECT 713.700 113.400 715.500 116.400 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 544.950 100.950 547.050 103.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 565.950 100.950 568.050 103.050 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 589.950 100.950 592.050 103.050 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 638.100 102.300 640.200 103.050 ;
        RECT 638.100 100.950 645.000 102.300 ;
        RECT 380.100 99.150 381.900 100.950 ;
        RECT 385.950 93.600 387.000 100.950 ;
        RECT 391.950 99.150 393.750 100.950 ;
        RECT 410.700 93.600 411.900 100.950 ;
        RECT 431.250 99.150 433.050 100.950 ;
        RECT 434.400 93.600 435.300 100.950 ;
        RECT 437.100 99.150 438.900 100.950 ;
        RECT 359.700 88.500 363.300 89.400 ;
        RECT 359.700 87.600 360.600 88.500 ;
        RECT 355.500 81.000 357.300 87.600 ;
        RECT 358.500 86.700 360.600 87.600 ;
        RECT 358.500 81.600 360.300 86.700 ;
        RECT 361.500 81.000 363.300 87.600 ;
        RECT 380.100 81.000 381.900 93.600 ;
        RECT 384.600 81.600 387.900 93.600 ;
        RECT 390.600 81.000 392.400 93.600 ;
        RECT 410.100 81.600 411.900 93.600 ;
        RECT 413.100 81.000 414.900 93.600 ;
        RECT 431.100 81.000 432.900 93.600 ;
        RECT 434.400 92.400 438.000 93.600 ;
        RECT 436.200 81.600 438.000 92.400 ;
        RECT 458.100 87.600 459.300 100.950 ;
        RECT 479.100 99.150 480.900 100.950 ;
        RECT 484.950 93.600 486.000 100.950 ;
        RECT 490.950 99.150 492.750 100.950 ;
        RECT 455.100 81.000 456.900 87.600 ;
        RECT 458.100 81.600 459.900 87.600 ;
        RECT 461.100 81.000 462.900 87.600 ;
        RECT 479.100 81.000 480.900 93.600 ;
        RECT 483.600 81.600 486.900 93.600 ;
        RECT 489.600 81.000 491.400 93.600 ;
        RECT 510.000 88.800 510.900 100.950 ;
        RECT 515.100 99.150 516.900 100.950 ;
        RECT 539.250 99.150 541.050 100.950 ;
        RECT 511.950 96.450 514.050 97.050 ;
        RECT 535.950 96.450 538.050 97.050 ;
        RECT 511.950 95.550 538.050 96.450 ;
        RECT 511.950 94.950 514.050 95.550 ;
        RECT 535.950 94.950 538.050 95.550 ;
        RECT 545.700 93.600 546.600 100.950 ;
        RECT 566.100 99.150 567.900 100.950 ;
        RECT 536.100 92.700 543.900 93.600 ;
        RECT 510.000 87.900 516.600 88.800 ;
        RECT 510.000 87.600 510.900 87.900 ;
        RECT 509.100 81.600 510.900 87.600 ;
        RECT 515.100 87.600 516.600 87.900 ;
        RECT 512.100 81.000 513.900 87.000 ;
        RECT 515.100 81.600 516.900 87.600 ;
        RECT 518.100 81.000 519.900 87.600 ;
        RECT 536.100 81.600 537.900 92.700 ;
        RECT 539.100 81.000 540.900 91.800 ;
        RECT 542.100 81.600 543.900 92.700 ;
        RECT 545.100 81.600 546.900 93.600 ;
        RECT 572.100 88.800 573.000 100.950 ;
        RECT 566.400 87.900 573.000 88.800 ;
        RECT 566.400 87.600 567.900 87.900 ;
        RECT 563.100 81.000 564.900 87.600 ;
        RECT 566.100 81.600 567.900 87.600 ;
        RECT 572.100 87.600 573.000 87.900 ;
        RECT 593.100 87.600 594.300 100.950 ;
        RECT 601.950 96.450 604.050 97.050 ;
        RECT 613.950 96.450 616.050 97.050 ;
        RECT 601.950 95.550 616.050 96.450 ;
        RECT 601.950 94.950 604.050 95.550 ;
        RECT 613.950 94.950 616.050 95.550 ;
        RECT 617.700 87.600 618.900 100.950 ;
        RECT 643.200 100.500 645.000 100.950 ;
        RECT 645.900 101.100 647.100 106.800 ;
        RECT 648.000 103.800 650.100 105.900 ;
        RECT 648.300 102.000 650.100 103.800 ;
        RECT 671.100 103.050 672.900 104.850 ;
        RECT 674.100 103.050 675.300 107.400 ;
        RECT 704.700 106.800 708.000 108.000 ;
        RECT 677.100 103.050 678.900 104.850 ;
        RECT 698.100 103.050 699.900 104.850 ;
        RECT 704.100 103.050 705.900 104.850 ;
        RECT 707.100 103.050 708.000 106.800 ;
        RECT 645.900 100.200 648.300 101.100 ;
        RECT 646.800 100.050 648.300 100.200 ;
        RECT 652.800 100.950 654.900 103.050 ;
        RECT 670.950 100.950 673.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 642.000 97.500 645.900 99.300 ;
        RECT 643.800 97.200 645.900 97.500 ;
        RECT 646.800 97.950 648.900 100.050 ;
        RECT 652.800 99.150 654.600 100.950 ;
        RECT 646.800 96.000 647.700 97.950 ;
        RECT 640.500 93.600 642.600 95.700 ;
        RECT 646.200 94.950 647.700 96.000 ;
        RECT 646.200 93.600 647.400 94.950 ;
        RECT 638.100 92.700 642.600 93.600 ;
        RECT 569.100 81.000 570.900 87.000 ;
        RECT 572.100 81.600 573.900 87.600 ;
        RECT 590.100 81.000 591.900 87.600 ;
        RECT 593.100 81.600 594.900 87.600 ;
        RECT 596.100 81.000 597.900 87.600 ;
        RECT 614.100 81.000 615.900 87.600 ;
        RECT 617.100 81.600 618.900 87.600 ;
        RECT 620.100 81.000 621.900 87.600 ;
        RECT 638.100 81.600 639.900 92.700 ;
        RECT 641.100 81.000 642.900 91.500 ;
        RECT 645.600 81.600 647.400 93.600 ;
        RECT 650.100 93.600 652.200 94.500 ;
        RECT 674.100 93.600 675.300 100.950 ;
        RECT 680.100 99.150 681.900 100.950 ;
        RECT 701.100 99.150 702.900 100.950 ;
        RECT 688.950 96.450 691.050 97.050 ;
        RECT 703.950 96.450 706.050 97.050 ;
        RECT 688.950 95.550 706.050 96.450 ;
        RECT 688.950 94.950 691.050 95.550 ;
        RECT 703.950 94.950 706.050 95.550 ;
        RECT 650.100 92.400 654.900 93.600 ;
        RECT 650.100 81.000 651.900 91.500 ;
        RECT 653.100 81.600 654.900 92.400 ;
        RECT 674.100 92.100 676.500 93.600 ;
        RECT 672.000 89.100 673.800 90.900 ;
        RECT 671.700 81.000 673.500 87.600 ;
        RECT 674.700 81.600 676.500 92.100 ;
        RECT 679.800 81.000 681.600 93.600 ;
        RECT 707.100 88.800 708.000 100.950 ;
        RECT 714.000 100.050 715.500 113.400 ;
        RECT 713.100 97.950 715.500 100.050 ;
        RECT 701.400 87.900 708.000 88.800 ;
        RECT 701.400 87.600 702.900 87.900 ;
        RECT 698.100 81.000 699.900 87.600 ;
        RECT 701.100 81.600 702.900 87.600 ;
        RECT 707.100 87.600 708.000 87.900 ;
        RECT 714.000 87.600 715.500 97.950 ;
        RECT 717.300 110.400 719.100 116.400 ;
        RECT 722.700 110.400 724.500 117.000 ;
        RECT 727.800 111.600 729.600 116.400 ;
        RECT 732.000 113.400 733.800 116.400 ;
        RECT 735.000 113.400 736.800 116.400 ;
        RECT 738.000 113.400 739.800 116.400 ;
        RECT 741.000 113.400 742.800 116.400 ;
        RECT 744.000 113.400 745.800 117.000 ;
        RECT 725.400 110.400 729.600 111.600 ;
        RECT 731.700 111.300 733.800 113.400 ;
        RECT 734.700 111.300 736.800 113.400 ;
        RECT 737.700 111.300 739.800 113.400 ;
        RECT 740.700 111.300 742.800 113.400 ;
        RECT 747.000 112.500 748.800 116.400 ;
        RECT 751.500 113.400 753.300 117.000 ;
        RECT 754.500 113.400 756.300 116.400 ;
        RECT 757.500 113.400 759.300 116.400 ;
        RECT 760.500 113.400 762.300 116.400 ;
        RECT 746.100 110.400 748.800 112.500 ;
        RECT 750.600 111.600 752.400 112.500 ;
        RECT 750.600 110.400 753.300 111.600 ;
        RECT 754.200 111.300 756.300 113.400 ;
        RECT 757.200 111.300 759.300 113.400 ;
        RECT 760.200 111.300 762.300 113.400 ;
        RECT 764.700 110.400 766.500 116.400 ;
        RECT 770.100 110.400 771.900 117.000 ;
        RECT 775.500 110.400 777.300 116.400 ;
        RECT 717.300 93.600 718.200 110.400 ;
        RECT 725.400 107.100 726.900 110.400 ;
        RECT 731.100 108.600 737.700 110.400 ;
        RECT 752.400 109.800 753.300 110.400 ;
        RECT 755.400 109.800 757.200 110.400 ;
        RECT 752.400 108.600 759.600 109.800 ;
        RECT 719.100 105.300 726.900 107.100 ;
        RECT 743.100 106.500 744.900 108.300 ;
        RECT 742.800 105.900 744.900 106.500 ;
        RECT 727.800 104.400 744.900 105.900 ;
        RECT 749.100 105.900 751.200 106.050 ;
        RECT 752.400 105.900 754.200 106.800 ;
        RECT 749.100 105.000 754.200 105.900 ;
        RECT 758.700 105.600 759.600 108.600 ;
        RECT 764.700 109.500 766.200 110.400 ;
        RECT 764.700 108.300 773.100 109.500 ;
        RECT 771.300 107.700 773.100 108.300 ;
        RECT 760.500 106.800 762.600 107.700 ;
        RECT 776.100 106.800 777.300 110.400 ;
        RECT 794.700 109.200 796.500 116.400 ;
        RECT 799.800 110.400 801.600 117.000 ;
        RECT 818.100 113.400 819.900 117.000 ;
        RECT 821.100 113.400 822.900 116.400 ;
        RECT 824.100 113.400 825.900 117.000 ;
        RECT 794.700 108.300 798.900 109.200 ;
        RECT 760.500 105.600 777.300 106.800 ;
        RECT 722.700 102.900 729.300 104.400 ;
        RECT 749.100 103.950 751.200 105.000 ;
        RECT 757.800 103.800 759.600 105.600 ;
        RECT 722.700 100.050 724.200 102.900 ;
        RECT 730.500 101.700 774.900 102.900 ;
        RECT 730.500 100.200 731.400 101.700 ;
        RECT 722.100 97.950 724.200 100.050 ;
        RECT 726.300 98.400 731.400 100.200 ;
        RECT 734.100 99.900 747.600 100.800 ;
        RECT 754.800 99.900 756.600 100.500 ;
        RECT 773.100 100.050 774.900 101.700 ;
        RECT 734.100 98.700 735.000 99.900 ;
        RECT 734.100 96.900 735.900 98.700 ;
        RECT 740.100 97.200 744.000 99.000 ;
        RECT 745.500 98.700 756.600 99.900 ;
        RECT 767.100 99.750 769.200 100.050 ;
        RECT 745.500 97.800 747.600 98.700 ;
        RECT 765.300 97.950 769.200 99.750 ;
        RECT 773.100 97.950 775.200 100.050 ;
        RECT 765.300 97.200 767.100 97.950 ;
        RECT 740.100 96.900 742.200 97.200 ;
        RECT 753.600 96.300 767.100 97.200 ;
        RECT 719.100 95.700 720.900 96.300 ;
        RECT 753.600 95.700 754.800 96.300 ;
        RECT 719.100 94.500 754.800 95.700 ;
        RECT 757.500 94.500 759.600 94.800 ;
        RECT 717.300 92.700 733.800 93.600 ;
        RECT 717.300 89.400 718.200 92.700 ;
        RECT 722.100 90.600 727.800 91.800 ;
        RECT 731.700 91.500 733.800 92.700 ;
        RECT 737.100 92.400 754.800 93.600 ;
        RECT 757.500 93.300 769.500 94.500 ;
        RECT 757.500 92.700 759.600 93.300 ;
        RECT 767.700 92.700 769.500 93.300 ;
        RECT 737.100 91.500 739.200 92.400 ;
        RECT 753.600 91.800 754.800 92.400 ;
        RECT 771.000 91.800 772.800 92.100 ;
        RECT 722.100 90.000 723.900 90.600 ;
        RECT 717.300 88.500 721.200 89.400 ;
        RECT 720.000 87.600 721.200 88.500 ;
        RECT 726.600 87.600 727.800 90.600 ;
        RECT 728.700 89.700 730.500 90.300 ;
        RECT 728.700 88.500 736.800 89.700 ;
        RECT 734.700 87.600 736.800 88.500 ;
        RECT 740.100 87.600 742.800 91.500 ;
        RECT 745.500 89.100 748.800 91.200 ;
        RECT 753.600 90.600 772.800 91.800 ;
        RECT 704.100 81.000 705.900 87.000 ;
        RECT 707.100 81.600 708.900 87.600 ;
        RECT 710.700 81.000 712.500 87.600 ;
        RECT 713.700 81.600 715.500 87.600 ;
        RECT 717.000 81.000 718.800 87.600 ;
        RECT 720.000 81.600 721.800 87.600 ;
        RECT 723.000 81.000 724.800 87.600 ;
        RECT 726.000 81.600 727.800 87.600 ;
        RECT 729.000 81.000 730.800 87.600 ;
        RECT 731.700 84.600 733.800 86.700 ;
        RECT 734.700 84.600 736.800 86.700 ;
        RECT 737.700 84.600 739.800 86.700 ;
        RECT 732.000 81.600 733.800 84.600 ;
        RECT 735.000 81.600 736.800 84.600 ;
        RECT 738.000 81.600 739.800 84.600 ;
        RECT 741.000 81.600 742.800 87.600 ;
        RECT 744.000 81.000 745.800 87.600 ;
        RECT 747.000 81.600 748.800 89.100 ;
        RECT 754.200 87.600 756.300 89.700 ;
        RECT 750.900 81.000 752.700 87.600 ;
        RECT 753.900 81.600 755.700 87.600 ;
        RECT 756.600 84.600 758.700 86.700 ;
        RECT 759.600 84.600 761.700 86.700 ;
        RECT 756.900 81.600 758.700 84.600 ;
        RECT 759.900 81.600 761.700 84.600 ;
        RECT 763.500 81.000 765.300 87.600 ;
        RECT 766.500 81.600 768.300 90.600 ;
        RECT 771.000 90.300 772.800 90.600 ;
        RECT 776.100 89.400 777.300 105.600 ;
        RECT 794.100 103.050 795.900 104.850 ;
        RECT 797.700 103.050 798.900 108.300 ;
        RECT 799.950 103.050 801.750 104.850 ;
        RECT 821.700 103.050 822.600 113.400 ;
        RECT 842.100 110.400 843.900 117.000 ;
        RECT 845.100 110.400 846.900 116.400 ;
        RECT 863.100 112.200 864.900 115.200 ;
        RECT 866.100 114.600 867.300 117.000 ;
        RECT 875.100 115.200 876.300 117.000 ;
        RECT 842.100 103.050 843.900 104.850 ;
        RECT 845.100 103.050 846.300 110.400 ;
        RECT 863.100 108.900 864.000 112.200 ;
        RECT 866.100 109.800 867.900 114.600 ;
        RECT 870.600 110.700 872.400 115.200 ;
        RECT 870.600 109.800 872.700 110.700 ;
        RECT 863.100 108.000 870.300 108.900 ;
        RECT 863.100 103.050 864.900 104.850 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 863.100 100.950 865.200 103.050 ;
        RECT 866.100 100.950 868.200 103.050 ;
        RECT 869.100 100.950 870.300 108.000 ;
        RECT 871.800 103.050 872.700 109.800 ;
        RECT 875.100 109.200 876.900 115.200 ;
        RECT 878.700 110.400 880.500 116.400 ;
        RECT 884.100 110.400 885.900 117.000 ;
        RECT 889.500 110.400 891.300 116.400 ;
        RECT 893.700 113.400 895.500 116.400 ;
        RECT 896.700 113.400 898.500 116.400 ;
        RECT 899.700 113.400 901.500 116.400 ;
        RECT 902.700 113.400 904.500 117.000 ;
        RECT 893.700 111.300 895.800 113.400 ;
        RECT 896.700 111.300 898.800 113.400 ;
        RECT 899.700 111.300 901.800 113.400 ;
        RECT 907.200 112.500 909.000 116.400 ;
        RECT 910.200 113.400 912.000 117.000 ;
        RECT 913.200 113.400 915.000 116.400 ;
        RECT 916.200 113.400 918.000 116.400 ;
        RECT 919.200 113.400 921.000 116.400 ;
        RECT 922.200 113.400 924.000 116.400 ;
        RECT 903.600 111.600 905.400 112.500 ;
        RECT 902.700 110.400 905.400 111.600 ;
        RECT 907.200 110.400 909.900 112.500 ;
        RECT 913.200 111.300 915.300 113.400 ;
        RECT 916.200 111.300 918.300 113.400 ;
        RECT 919.200 111.300 921.300 113.400 ;
        RECT 922.200 111.300 924.300 113.400 ;
        RECT 926.400 111.600 928.200 116.400 ;
        RECT 926.400 110.400 930.600 111.600 ;
        RECT 931.500 110.400 933.300 117.000 ;
        RECT 936.900 110.400 938.700 116.400 ;
        RECT 878.700 106.800 879.900 110.400 ;
        RECT 889.800 109.500 891.300 110.400 ;
        RECT 898.800 109.800 900.600 110.400 ;
        RECT 902.700 109.800 903.600 110.400 ;
        RECT 882.900 108.300 891.300 109.500 ;
        RECT 896.400 108.600 903.600 109.800 ;
        RECT 918.300 108.600 924.900 110.400 ;
        RECT 882.900 107.700 884.700 108.300 ;
        RECT 893.400 106.800 895.500 107.700 ;
        RECT 878.700 105.600 895.500 106.800 ;
        RECT 896.400 105.600 897.300 108.600 ;
        RECT 901.800 105.900 903.600 106.800 ;
        RECT 911.100 106.500 912.900 108.300 ;
        RECT 929.100 107.100 930.600 110.400 ;
        RECT 904.800 105.900 906.900 106.050 ;
        RECT 871.800 100.950 873.900 103.050 ;
        RECT 874.800 100.950 876.900 103.050 ;
        RECT 773.700 88.500 777.300 89.400 ;
        RECT 773.700 87.600 774.600 88.500 ;
        RECT 797.700 87.600 798.900 100.950 ;
        RECT 818.100 99.150 819.900 100.950 ;
        RECT 821.700 93.600 822.600 100.950 ;
        RECT 823.950 99.150 825.750 100.950 ;
        RECT 845.100 93.600 846.300 100.950 ;
        RECT 866.100 99.150 867.900 100.950 ;
        RECT 869.100 99.150 870.900 100.950 ;
        RECT 869.700 94.800 870.900 99.150 ;
        RECT 863.100 93.900 870.900 94.800 ;
        RECT 819.000 92.400 822.600 93.600 ;
        RECT 769.500 81.000 771.300 87.600 ;
        RECT 772.500 86.700 774.600 87.600 ;
        RECT 772.500 81.600 774.300 86.700 ;
        RECT 775.500 81.000 777.300 87.600 ;
        RECT 794.100 81.000 795.900 87.600 ;
        RECT 797.100 81.600 798.900 87.600 ;
        RECT 800.100 81.000 801.900 87.600 ;
        RECT 819.000 81.600 820.800 92.400 ;
        RECT 824.100 81.000 825.900 93.600 ;
        RECT 842.100 81.000 843.900 93.600 ;
        RECT 845.100 81.600 846.900 93.600 ;
        RECT 863.100 88.800 864.000 93.900 ;
        RECT 871.800 93.000 872.700 100.950 ;
        RECT 874.800 99.150 876.600 100.950 ;
        RECT 863.100 82.800 864.900 88.800 ;
        RECT 866.100 81.000 867.900 93.000 ;
        RECT 870.600 92.100 872.700 93.000 ;
        RECT 870.600 81.600 872.400 92.100 ;
        RECT 875.100 81.000 876.900 93.600 ;
        RECT 878.700 89.400 879.900 105.600 ;
        RECT 896.400 103.800 898.200 105.600 ;
        RECT 901.800 105.000 906.900 105.900 ;
        RECT 904.800 103.950 906.900 105.000 ;
        RECT 911.100 105.900 913.200 106.500 ;
        RECT 911.100 104.400 928.200 105.900 ;
        RECT 929.100 105.300 936.900 107.100 ;
        RECT 926.700 102.900 933.300 104.400 ;
        RECT 881.100 101.700 925.500 102.900 ;
        RECT 881.100 100.050 882.900 101.700 ;
        RECT 880.800 97.950 882.900 100.050 ;
        RECT 886.800 99.750 888.900 100.050 ;
        RECT 899.400 99.900 901.200 100.500 ;
        RECT 908.400 99.900 921.900 100.800 ;
        RECT 886.800 97.950 890.700 99.750 ;
        RECT 899.400 98.700 910.500 99.900 ;
        RECT 888.900 97.200 890.700 97.950 ;
        RECT 908.400 97.800 910.500 98.700 ;
        RECT 912.000 97.200 915.900 99.000 ;
        RECT 921.000 98.700 921.900 99.900 ;
        RECT 888.900 96.300 902.400 97.200 ;
        RECT 913.800 96.900 915.900 97.200 ;
        RECT 920.100 96.900 921.900 98.700 ;
        RECT 924.600 100.200 925.500 101.700 ;
        RECT 924.600 98.400 929.700 100.200 ;
        RECT 931.800 100.050 933.300 102.900 ;
        RECT 931.800 97.950 933.900 100.050 ;
        RECT 901.200 95.700 902.400 96.300 ;
        RECT 935.100 95.700 936.900 96.300 ;
        RECT 896.400 94.500 898.500 94.800 ;
        RECT 901.200 94.500 936.900 95.700 ;
        RECT 886.500 93.300 898.500 94.500 ;
        RECT 937.800 93.600 938.700 110.400 ;
        RECT 886.500 92.700 888.300 93.300 ;
        RECT 896.400 92.700 898.500 93.300 ;
        RECT 901.200 92.400 918.900 93.600 ;
        RECT 883.200 91.800 885.000 92.100 ;
        RECT 901.200 91.800 902.400 92.400 ;
        RECT 883.200 90.600 902.400 91.800 ;
        RECT 916.800 91.500 918.900 92.400 ;
        RECT 922.200 92.700 938.700 93.600 ;
        RECT 922.200 91.500 924.300 92.700 ;
        RECT 883.200 90.300 885.000 90.600 ;
        RECT 878.700 88.500 882.300 89.400 ;
        RECT 881.400 87.600 882.300 88.500 ;
        RECT 878.700 81.000 880.500 87.600 ;
        RECT 881.400 86.700 883.500 87.600 ;
        RECT 881.700 81.600 883.500 86.700 ;
        RECT 884.700 81.000 886.500 87.600 ;
        RECT 887.700 81.600 889.500 90.600 ;
        RECT 899.700 87.600 901.800 89.700 ;
        RECT 907.200 89.100 910.500 91.200 ;
        RECT 890.700 81.000 892.500 87.600 ;
        RECT 894.300 84.600 896.400 86.700 ;
        RECT 897.300 84.600 899.400 86.700 ;
        RECT 894.300 81.600 896.100 84.600 ;
        RECT 897.300 81.600 899.100 84.600 ;
        RECT 900.300 81.600 902.100 87.600 ;
        RECT 903.300 81.000 905.100 87.600 ;
        RECT 907.200 81.600 909.000 89.100 ;
        RECT 913.200 87.600 915.900 91.500 ;
        RECT 928.200 90.600 933.900 91.800 ;
        RECT 925.500 89.700 927.300 90.300 ;
        RECT 919.200 88.500 927.300 89.700 ;
        RECT 919.200 87.600 921.300 88.500 ;
        RECT 928.200 87.600 929.400 90.600 ;
        RECT 932.100 90.000 933.900 90.600 ;
        RECT 937.800 89.400 938.700 92.700 ;
        RECT 934.800 88.500 938.700 89.400 ;
        RECT 940.500 113.400 942.300 116.400 ;
        RECT 943.500 113.400 945.300 117.000 ;
        RECT 940.500 100.050 942.000 113.400 ;
        RECT 962.100 110.400 963.900 116.400 ;
        RECT 965.100 111.300 966.900 117.000 ;
        RECT 969.300 111.000 971.100 116.400 ;
        RECT 973.800 111.300 975.600 117.000 ;
        RECT 962.100 109.500 963.600 110.400 ;
        RECT 962.100 108.000 966.600 109.500 ;
        RECT 964.500 107.400 966.600 108.000 ;
        RECT 970.200 108.900 971.100 111.000 ;
        RECT 977.100 110.400 978.900 116.400 ;
        RECT 995.400 110.400 997.200 117.000 ;
        RECT 974.400 109.500 978.900 110.400 ;
        RECT 967.500 105.900 969.300 107.700 ;
        RECT 970.200 106.800 973.200 108.900 ;
        RECT 974.400 107.100 976.500 109.500 ;
        RECT 1000.500 109.200 1002.300 116.400 ;
        RECT 1019.100 113.400 1020.900 116.400 ;
        RECT 1022.100 113.400 1023.900 117.000 ;
        RECT 998.100 108.300 1002.300 109.200 ;
        RECT 966.900 105.000 969.000 105.900 ;
        RECT 962.400 103.800 969.000 105.000 ;
        RECT 962.400 103.200 964.200 103.800 ;
        RECT 962.100 100.950 964.200 103.200 ;
        RECT 966.900 100.800 969.000 102.900 ;
        RECT 940.500 97.950 942.900 100.050 ;
        RECT 966.900 99.000 968.700 100.800 ;
        RECT 970.200 100.050 971.100 106.800 ;
        RECT 972.000 102.900 974.100 105.000 ;
        RECT 995.250 103.050 997.050 104.850 ;
        RECT 998.100 103.050 999.300 108.300 ;
        RECT 1001.100 103.050 1002.900 104.850 ;
        RECT 1019.700 103.050 1020.900 113.400 ;
        RECT 972.000 101.100 973.800 102.900 ;
        RECT 976.800 100.950 978.900 103.050 ;
        RECT 994.950 100.950 997.050 103.050 ;
        RECT 997.950 100.950 1000.050 103.050 ;
        RECT 1000.950 100.950 1003.050 103.050 ;
        RECT 1018.950 100.950 1021.050 103.050 ;
        RECT 1021.950 100.950 1024.050 103.050 ;
        RECT 970.200 98.700 973.200 100.050 ;
        RECT 976.800 99.150 978.600 100.950 ;
        RECT 971.100 97.950 973.200 98.700 ;
        RECT 934.800 87.600 936.000 88.500 ;
        RECT 940.500 87.600 942.000 97.950 ;
        RECT 968.400 95.700 970.200 97.500 ;
        RECT 964.800 94.800 970.200 95.700 ;
        RECT 964.800 93.900 966.900 94.800 ;
        RECT 962.100 92.700 966.900 93.900 ;
        RECT 971.700 93.600 972.900 97.950 ;
        RECT 969.600 92.700 972.900 93.600 ;
        RECT 973.800 93.600 975.900 94.500 ;
        RECT 910.200 81.000 912.000 87.600 ;
        RECT 913.200 81.600 915.000 87.600 ;
        RECT 916.200 84.600 918.300 86.700 ;
        RECT 919.200 84.600 921.300 86.700 ;
        RECT 922.200 84.600 924.300 86.700 ;
        RECT 916.200 81.600 918.000 84.600 ;
        RECT 919.200 81.600 921.000 84.600 ;
        RECT 922.200 81.600 924.000 84.600 ;
        RECT 925.200 81.000 927.000 87.600 ;
        RECT 928.200 81.600 930.000 87.600 ;
        RECT 931.200 81.000 933.000 87.600 ;
        RECT 934.200 81.600 936.000 87.600 ;
        RECT 937.200 81.000 939.000 87.600 ;
        RECT 940.500 81.600 942.300 87.600 ;
        RECT 943.500 81.000 945.300 87.600 ;
        RECT 962.100 81.600 963.900 92.700 ;
        RECT 965.100 81.000 966.900 91.500 ;
        RECT 969.600 81.600 971.400 92.700 ;
        RECT 973.800 92.400 978.900 93.600 ;
        RECT 973.800 81.000 975.900 91.500 ;
        RECT 977.100 81.600 978.900 92.400 ;
        RECT 998.100 87.600 999.300 100.950 ;
        RECT 1019.700 87.600 1020.900 100.950 ;
        RECT 1022.100 99.150 1023.900 100.950 ;
        RECT 995.100 81.000 996.900 87.600 ;
        RECT 998.100 81.600 999.900 87.600 ;
        RECT 1001.100 81.000 1002.900 87.600 ;
        RECT 1019.100 81.600 1020.900 87.600 ;
        RECT 1022.100 81.000 1023.900 87.600 ;
        RECT 17.100 71.400 18.900 78.000 ;
        RECT 20.100 71.400 21.900 77.400 ;
        RECT 23.100 71.400 24.900 78.000 ;
        RECT 20.700 58.050 21.900 71.400 ;
        RECT 41.100 65.400 42.900 77.400 ;
        RECT 45.600 65.400 47.400 78.000 ;
        RECT 48.600 66.900 50.400 77.400 ;
        RECT 48.600 65.400 51.000 66.900 ;
        RECT 68.100 66.300 69.900 77.400 ;
        RECT 71.100 67.200 72.900 78.000 ;
        RECT 74.100 66.300 75.900 77.400 ;
        RECT 68.100 65.400 75.900 66.300 ;
        RECT 77.100 65.400 78.900 77.400 ;
        RECT 95.100 71.400 96.900 78.000 ;
        RECT 98.100 71.400 99.900 77.400 ;
        RECT 101.100 72.000 102.900 78.000 ;
        RECT 98.400 71.100 99.900 71.400 ;
        RECT 104.100 71.400 105.900 77.400 ;
        RECT 104.100 71.100 105.000 71.400 ;
        RECT 98.400 70.200 105.000 71.100 ;
        RECT 41.100 63.900 42.300 65.400 ;
        RECT 41.100 62.700 48.900 63.900 ;
        RECT 47.100 62.100 48.900 62.700 ;
        RECT 45.000 58.050 46.800 59.850 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 41.100 55.950 43.200 58.050 ;
        RECT 44.400 55.950 46.500 58.050 ;
        RECT 17.100 54.150 18.900 55.950 ;
        RECT 20.700 50.700 21.900 55.950 ;
        RECT 22.950 54.150 24.750 55.950 ;
        RECT 41.400 54.150 43.200 55.950 ;
        RECT 47.700 51.600 48.600 62.100 ;
        RECT 49.800 58.050 51.000 65.400 ;
        RECT 71.250 58.050 73.050 59.850 ;
        RECT 77.700 58.050 78.600 65.400 ;
        RECT 91.950 63.450 94.050 64.050 ;
        RECT 100.950 63.450 103.050 64.050 ;
        RECT 91.950 62.550 103.050 63.450 ;
        RECT 91.950 61.950 94.050 62.550 ;
        RECT 100.950 61.950 103.050 62.550 ;
        RECT 98.100 58.050 99.900 59.850 ;
        RECT 104.100 58.050 105.000 70.200 ;
        RECT 123.000 66.600 124.800 77.400 ;
        RECT 123.000 65.400 126.600 66.600 ;
        RECT 128.100 65.400 129.900 78.000 ;
        RECT 146.100 65.400 147.900 78.000 ;
        RECT 149.100 65.400 150.900 77.400 ;
        RECT 167.100 71.400 168.900 78.000 ;
        RECT 170.100 71.400 171.900 77.400 ;
        RECT 122.100 58.050 123.900 59.850 ;
        RECT 125.700 58.050 126.600 65.400 ;
        RECT 127.950 58.050 129.750 59.850 ;
        RECT 149.100 58.050 150.300 65.400 ;
        RECT 167.100 58.050 168.900 59.850 ;
        RECT 170.100 58.050 171.300 71.400 ;
        RECT 189.000 66.600 190.800 77.400 ;
        RECT 189.000 65.400 192.600 66.600 ;
        RECT 194.100 65.400 195.900 78.000 ;
        RECT 212.100 65.400 213.900 78.000 ;
        RECT 217.200 66.600 219.000 77.400 ;
        RECT 215.400 65.400 219.000 66.600 ;
        RECT 236.100 65.400 237.900 77.400 ;
        RECT 239.100 65.400 240.900 78.000 ;
        RECT 257.100 65.400 258.900 78.000 ;
        RECT 262.200 66.600 264.000 77.400 ;
        RECT 260.400 65.400 264.000 66.600 ;
        RECT 281.100 65.400 282.900 78.000 ;
        RECT 285.600 65.400 288.900 77.400 ;
        RECT 291.600 65.400 293.400 78.000 ;
        RECT 311.100 65.400 312.900 78.000 ;
        RECT 315.600 65.400 318.900 77.400 ;
        RECT 321.600 65.400 323.400 78.000 ;
        RECT 341.100 71.400 342.900 78.000 ;
        RECT 344.100 71.400 345.900 77.400 ;
        RECT 347.100 71.400 348.900 78.000 ;
        RECT 188.100 58.050 189.900 59.850 ;
        RECT 191.700 58.050 192.600 65.400 ;
        RECT 193.950 58.050 195.750 59.850 ;
        RECT 212.250 58.050 214.050 59.850 ;
        RECT 215.400 58.050 216.300 65.400 ;
        RECT 218.100 58.050 219.900 59.850 ;
        RECT 236.700 58.050 237.900 65.400 ;
        RECT 257.250 58.050 259.050 59.850 ;
        RECT 260.400 58.050 261.300 65.400 ;
        RECT 263.100 58.050 264.900 59.850 ;
        RECT 281.100 58.050 282.900 59.850 ;
        RECT 286.950 58.050 288.000 65.400 ;
        RECT 289.950 63.450 292.050 64.050 ;
        RECT 307.950 63.450 310.050 64.050 ;
        RECT 289.950 62.550 310.050 63.450 ;
        RECT 289.950 61.950 292.050 62.550 ;
        RECT 307.950 61.950 310.050 62.550 ;
        RECT 292.950 58.050 294.750 59.850 ;
        RECT 311.100 58.050 312.900 59.850 ;
        RECT 316.950 58.050 318.000 65.400 ;
        RECT 322.950 58.050 324.750 59.850 ;
        RECT 344.100 58.050 345.300 71.400 ;
        RECT 365.100 65.400 366.900 78.000 ;
        RECT 368.100 65.400 369.900 77.400 ;
        RECT 370.950 72.450 373.050 73.050 ;
        RECT 379.950 72.450 382.050 73.050 ;
        RECT 370.950 71.550 382.050 72.450 ;
        RECT 370.950 70.950 373.050 71.550 ;
        RECT 379.950 70.950 382.050 71.550 ;
        RECT 386.100 71.400 387.900 78.000 ;
        RECT 389.100 71.400 390.900 77.400 ;
        RECT 392.100 71.400 393.900 78.000 ;
        RECT 410.100 71.400 411.900 78.000 ;
        RECT 413.100 71.400 414.900 77.400 ;
        RECT 416.100 71.400 417.900 78.000 ;
        RECT 434.700 71.400 436.500 78.000 ;
        RECT 368.100 58.050 369.300 65.400 ;
        RECT 389.100 58.050 390.300 71.400 ;
        RECT 403.950 63.450 406.050 64.050 ;
        RECT 409.950 63.450 412.050 64.050 ;
        RECT 403.950 62.550 412.050 63.450 ;
        RECT 403.950 61.950 406.050 62.550 ;
        RECT 409.950 61.950 412.050 62.550 ;
        RECT 413.700 58.050 414.900 71.400 ;
        RECT 435.000 68.100 436.800 69.900 ;
        RECT 437.700 66.900 439.500 77.400 ;
        RECT 437.100 65.400 439.500 66.900 ;
        RECT 442.800 65.400 444.600 78.000 ;
        RECT 461.100 66.300 462.900 77.400 ;
        RECT 464.100 67.500 465.900 78.000 ;
        RECT 468.600 66.300 470.400 77.400 ;
        RECT 472.800 67.500 474.900 78.000 ;
        RECT 476.100 66.600 477.900 77.400 ;
        RECT 495.600 66.900 497.400 77.400 ;
        RECT 437.100 58.050 438.300 65.400 ;
        RECT 461.100 65.100 465.900 66.300 ;
        RECT 468.600 65.400 471.900 66.300 ;
        RECT 463.800 64.200 465.900 65.100 ;
        RECT 463.800 63.300 469.200 64.200 ;
        RECT 467.400 61.500 469.200 63.300 ;
        RECT 470.700 61.050 471.900 65.400 ;
        RECT 472.800 65.400 477.900 66.600 ;
        RECT 495.000 65.400 497.400 66.900 ;
        RECT 498.600 65.400 500.400 78.000 ;
        RECT 503.100 65.400 504.900 77.400 ;
        RECT 522.600 66.900 524.400 77.400 ;
        RECT 472.800 64.500 474.900 65.400 ;
        RECT 470.100 60.300 472.200 61.050 ;
        RECT 443.100 58.050 444.900 59.850 ;
        RECT 465.900 58.200 467.700 60.000 ;
        RECT 469.200 58.950 472.200 60.300 ;
        RECT 49.800 55.950 51.900 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 70.950 55.950 73.050 58.050 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 94.950 55.950 97.050 58.050 ;
        RECT 97.950 55.950 100.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 47.700 50.700 49.800 51.600 ;
        RECT 17.700 49.800 21.900 50.700 ;
        RECT 44.400 49.800 49.800 50.700 ;
        RECT 17.700 42.600 19.500 49.800 ;
        RECT 22.800 42.000 24.600 48.600 ;
        RECT 44.400 45.600 45.300 49.800 ;
        RECT 51.000 48.600 51.900 55.950 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 74.250 54.150 76.050 55.950 ;
        RECT 77.700 48.600 78.600 55.950 ;
        RECT 95.100 54.150 96.900 55.950 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 104.100 52.200 105.000 55.950 ;
        RECT 41.100 42.600 42.900 45.600 ;
        RECT 44.100 42.600 45.900 45.600 ;
        RECT 41.100 42.000 42.300 42.600 ;
        RECT 47.100 42.000 48.900 48.000 ;
        RECT 50.100 42.600 51.900 48.600 ;
        RECT 69.000 42.000 70.800 48.600 ;
        RECT 73.500 47.400 78.600 48.600 ;
        RECT 73.500 42.600 75.300 47.400 ;
        RECT 76.500 42.000 78.300 45.600 ;
        RECT 95.100 42.000 96.900 51.600 ;
        RECT 101.700 51.000 105.000 52.200 ;
        RECT 101.700 42.600 103.500 51.000 ;
        RECT 125.700 45.600 126.600 55.950 ;
        RECT 146.100 54.150 147.900 55.950 ;
        RECT 149.100 48.600 150.300 55.950 ;
        RECT 122.100 42.000 123.900 45.600 ;
        RECT 125.100 42.600 126.900 45.600 ;
        RECT 128.100 42.000 129.900 45.600 ;
        RECT 146.100 42.000 147.900 48.600 ;
        RECT 149.100 42.600 150.900 48.600 ;
        RECT 170.100 45.600 171.300 55.950 ;
        RECT 191.700 45.600 192.600 55.950 ;
        RECT 215.400 45.600 216.300 55.950 ;
        RECT 236.700 48.600 237.900 55.950 ;
        RECT 239.100 54.150 240.900 55.950 ;
        RECT 167.100 42.000 168.900 45.600 ;
        RECT 170.100 42.600 171.900 45.600 ;
        RECT 188.100 42.000 189.900 45.600 ;
        RECT 191.100 42.600 192.900 45.600 ;
        RECT 194.100 42.000 195.900 45.600 ;
        RECT 212.100 42.000 213.900 45.600 ;
        RECT 215.100 42.600 216.900 45.600 ;
        RECT 218.100 42.000 219.900 45.600 ;
        RECT 236.100 42.600 237.900 48.600 ;
        RECT 239.100 42.000 240.900 48.600 ;
        RECT 260.400 45.600 261.300 55.950 ;
        RECT 284.250 54.150 286.050 55.950 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 286.950 51.300 288.000 55.950 ;
        RECT 289.950 54.150 291.750 55.950 ;
        RECT 314.250 54.150 316.050 55.950 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 316.950 51.300 318.000 55.950 ;
        RECT 319.950 54.150 321.750 55.950 ;
        RECT 341.250 54.150 343.050 55.950 ;
        RECT 286.950 50.100 291.300 51.300 ;
        RECT 316.950 50.100 321.300 51.300 ;
        RECT 281.100 48.000 288.900 48.900 ;
        RECT 290.400 48.600 291.300 50.100 ;
        RECT 257.100 42.000 258.900 45.600 ;
        RECT 260.100 42.600 261.900 45.600 ;
        RECT 263.100 42.000 264.900 45.600 ;
        RECT 281.100 42.600 282.900 48.000 ;
        RECT 284.100 42.000 285.900 47.100 ;
        RECT 287.100 43.500 288.900 48.000 ;
        RECT 290.100 44.400 291.900 48.600 ;
        RECT 293.100 43.500 294.900 48.600 ;
        RECT 287.100 42.600 294.900 43.500 ;
        RECT 311.100 48.000 318.900 48.900 ;
        RECT 320.400 48.600 321.300 50.100 ;
        RECT 344.100 50.700 345.300 55.950 ;
        RECT 347.100 54.150 348.900 55.950 ;
        RECT 365.100 54.150 366.900 55.950 ;
        RECT 355.950 51.450 358.050 52.050 ;
        RECT 364.950 51.450 367.050 52.050 ;
        RECT 344.100 49.800 348.300 50.700 ;
        RECT 355.950 50.550 367.050 51.450 ;
        RECT 355.950 49.950 358.050 50.550 ;
        RECT 364.950 49.950 367.050 50.550 ;
        RECT 311.100 42.600 312.900 48.000 ;
        RECT 314.100 42.000 315.900 47.100 ;
        RECT 317.100 43.500 318.900 48.000 ;
        RECT 320.100 44.400 321.900 48.600 ;
        RECT 323.100 43.500 324.900 48.600 ;
        RECT 317.100 42.600 324.900 43.500 ;
        RECT 341.400 42.000 343.200 48.600 ;
        RECT 346.500 42.600 348.300 49.800 ;
        RECT 368.100 48.600 369.300 55.950 ;
        RECT 386.250 54.150 388.050 55.950 ;
        RECT 389.100 50.700 390.300 55.950 ;
        RECT 392.100 54.150 393.900 55.950 ;
        RECT 410.100 54.150 411.900 55.950 ;
        RECT 413.700 50.700 414.900 55.950 ;
        RECT 415.950 54.150 417.750 55.950 ;
        RECT 434.100 54.150 435.900 55.950 ;
        RECT 437.100 51.600 438.300 55.950 ;
        RECT 440.100 54.150 441.900 55.950 ;
        RECT 461.100 55.800 463.200 58.050 ;
        RECT 465.900 56.100 468.000 58.200 ;
        RECT 461.400 55.200 463.200 55.800 ;
        RECT 461.400 54.000 468.000 55.200 ;
        RECT 465.900 53.100 468.000 54.000 ;
        RECT 389.100 49.800 393.300 50.700 ;
        RECT 365.100 42.000 366.900 48.600 ;
        RECT 368.100 42.600 369.900 48.600 ;
        RECT 386.400 42.000 388.200 48.600 ;
        RECT 391.500 42.600 393.300 49.800 ;
        RECT 410.700 49.800 414.900 50.700 ;
        RECT 434.700 50.700 438.300 51.600 ;
        RECT 463.500 51.000 465.600 51.600 ;
        RECT 466.500 51.300 468.300 53.100 ;
        RECT 469.200 52.200 470.100 58.950 ;
        RECT 475.800 58.050 477.600 59.850 ;
        RECT 495.000 58.050 496.200 65.400 ;
        RECT 503.700 63.900 504.900 65.400 ;
        RECT 497.100 62.700 504.900 63.900 ;
        RECT 522.000 65.400 524.400 66.900 ;
        RECT 525.600 65.400 527.400 78.000 ;
        RECT 530.100 65.400 531.900 77.400 ;
        RECT 497.100 62.100 498.900 62.700 ;
        RECT 471.000 56.100 472.800 57.900 ;
        RECT 471.000 54.000 473.100 56.100 ;
        RECT 475.800 55.950 477.900 58.050 ;
        RECT 494.100 55.950 496.200 58.050 ;
        RECT 410.700 42.600 412.500 49.800 ;
        RECT 434.700 48.600 435.900 50.700 ;
        RECT 461.100 49.500 465.600 51.000 ;
        RECT 469.200 50.100 472.200 52.200 ;
        RECT 415.800 42.000 417.600 48.600 ;
        RECT 434.100 42.600 435.900 48.600 ;
        RECT 437.100 47.700 444.900 49.050 ;
        RECT 437.100 42.600 438.900 47.700 ;
        RECT 440.100 42.000 441.900 46.800 ;
        RECT 443.100 42.600 444.900 47.700 ;
        RECT 461.100 48.600 462.600 49.500 ;
        RECT 461.100 42.600 462.900 48.600 ;
        RECT 469.200 48.000 470.100 50.100 ;
        RECT 473.400 49.500 475.500 51.900 ;
        RECT 473.400 48.600 477.900 49.500 ;
        RECT 464.100 42.000 465.900 47.700 ;
        RECT 468.300 42.600 470.100 48.000 ;
        RECT 472.800 42.000 474.600 47.700 ;
        RECT 476.100 42.600 477.900 48.600 ;
        RECT 494.100 48.600 495.000 55.950 ;
        RECT 497.400 51.600 498.300 62.100 ;
        RECT 499.200 58.050 501.000 59.850 ;
        RECT 522.000 58.050 523.200 65.400 ;
        RECT 530.700 63.900 531.900 65.400 ;
        RECT 548.100 66.300 549.900 77.400 ;
        RECT 551.100 67.500 552.900 78.000 ;
        RECT 555.600 66.300 557.400 77.400 ;
        RECT 559.800 67.500 561.900 78.000 ;
        RECT 563.100 66.600 564.900 77.400 ;
        RECT 548.100 65.100 552.900 66.300 ;
        RECT 555.600 65.400 558.900 66.300 ;
        RECT 524.100 62.700 531.900 63.900 ;
        RECT 550.800 64.200 552.900 65.100 ;
        RECT 550.800 63.300 556.200 64.200 ;
        RECT 524.100 62.100 525.900 62.700 ;
        RECT 499.500 55.950 501.600 58.050 ;
        RECT 502.800 55.950 504.900 58.050 ;
        RECT 521.100 55.950 523.200 58.050 ;
        RECT 502.800 54.150 504.600 55.950 ;
        RECT 496.200 50.700 498.300 51.600 ;
        RECT 496.200 49.800 501.600 50.700 ;
        RECT 494.100 42.600 495.900 48.600 ;
        RECT 497.100 42.000 498.900 48.000 ;
        RECT 500.700 45.600 501.600 49.800 ;
        RECT 521.100 48.600 522.000 55.950 ;
        RECT 524.400 51.600 525.300 62.100 ;
        RECT 554.400 61.500 556.200 63.300 ;
        RECT 557.700 61.050 558.900 65.400 ;
        RECT 559.800 65.400 564.900 66.600 ;
        RECT 581.100 66.600 582.900 77.400 ;
        RECT 584.100 67.500 585.900 78.000 ;
        RECT 581.100 65.400 585.900 66.600 ;
        RECT 559.800 64.500 561.900 65.400 ;
        RECT 583.800 64.500 585.900 65.400 ;
        RECT 588.600 65.400 590.400 77.400 ;
        RECT 593.100 67.500 594.900 78.000 ;
        RECT 596.100 66.300 597.900 77.400 ;
        RECT 593.400 65.400 597.900 66.300 ;
        RECT 614.400 65.400 616.200 78.000 ;
        RECT 619.500 66.900 621.300 77.400 ;
        RECT 622.500 71.400 624.300 78.000 ;
        RECT 641.100 71.400 642.900 78.000 ;
        RECT 644.100 71.400 645.900 77.400 ;
        RECT 647.100 71.400 648.900 78.000 ;
        RECT 665.100 71.400 666.900 78.000 ;
        RECT 668.100 71.400 669.900 77.400 ;
        RECT 671.100 71.400 672.900 78.000 ;
        RECT 689.100 71.400 690.900 78.000 ;
        RECT 692.100 71.400 693.900 77.400 ;
        RECT 622.200 68.100 624.000 69.900 ;
        RECT 619.500 65.400 621.900 66.900 ;
        RECT 588.600 64.050 589.800 65.400 ;
        RECT 588.300 63.000 589.800 64.050 ;
        RECT 593.400 63.300 595.500 65.400 ;
        RECT 588.300 61.050 589.200 63.000 ;
        RECT 557.100 60.300 559.200 61.050 ;
        RECT 526.200 58.050 528.000 59.850 ;
        RECT 552.900 58.200 554.700 60.000 ;
        RECT 556.200 58.950 559.200 60.300 ;
        RECT 526.500 55.950 528.600 58.050 ;
        RECT 529.800 55.950 531.900 58.050 ;
        RECT 529.800 54.150 531.600 55.950 ;
        RECT 548.100 55.800 550.200 58.050 ;
        RECT 552.900 56.100 555.000 58.200 ;
        RECT 548.400 55.200 550.200 55.800 ;
        RECT 548.400 54.000 555.000 55.200 ;
        RECT 552.900 53.100 555.000 54.000 ;
        RECT 523.200 50.700 525.300 51.600 ;
        RECT 550.500 51.000 552.600 51.600 ;
        RECT 553.500 51.300 555.300 53.100 ;
        RECT 556.200 52.200 557.100 58.950 ;
        RECT 562.800 58.050 564.600 59.850 ;
        RECT 581.400 58.050 583.200 59.850 ;
        RECT 587.100 58.950 589.200 61.050 ;
        RECT 590.100 61.500 592.200 61.800 ;
        RECT 590.100 59.700 594.000 61.500 ;
        RECT 558.000 56.100 559.800 57.900 ;
        RECT 558.000 54.000 560.100 56.100 ;
        RECT 562.800 55.950 564.900 58.050 ;
        RECT 581.100 55.950 583.200 58.050 ;
        RECT 587.700 58.800 589.200 58.950 ;
        RECT 587.700 57.900 590.100 58.800 ;
        RECT 585.900 55.200 587.700 57.000 ;
        RECT 585.900 53.100 588.000 55.200 ;
        RECT 588.900 52.200 590.100 57.900 ;
        RECT 591.000 58.050 592.800 58.500 ;
        RECT 614.100 58.050 615.900 59.850 ;
        RECT 620.700 58.050 621.900 65.400 ;
        RECT 644.700 58.050 645.900 71.400 ;
        RECT 668.700 58.050 669.900 71.400 ;
        RECT 670.950 63.450 673.050 64.050 ;
        RECT 676.950 63.450 679.050 64.050 ;
        RECT 670.950 62.550 679.050 63.450 ;
        RECT 670.950 61.950 673.050 62.550 ;
        RECT 676.950 61.950 679.050 62.550 ;
        RECT 689.100 58.050 690.900 59.850 ;
        RECT 692.100 58.050 693.300 71.400 ;
        RECT 710.400 65.400 712.200 78.000 ;
        RECT 715.500 66.900 717.300 77.400 ;
        RECT 718.500 71.400 720.300 78.000 ;
        RECT 737.700 71.400 739.500 78.000 ;
        RECT 718.200 68.100 720.000 69.900 ;
        RECT 738.000 68.100 739.800 69.900 ;
        RECT 740.700 66.900 742.500 77.400 ;
        RECT 715.500 65.400 717.900 66.900 ;
        RECT 710.100 58.050 711.900 59.850 ;
        RECT 716.700 58.050 717.900 65.400 ;
        RECT 740.100 65.400 742.500 66.900 ;
        RECT 745.800 65.400 747.600 78.000 ;
        RECT 764.100 71.400 765.900 77.400 ;
        RECT 767.100 71.400 768.900 78.000 ;
        RECT 770.700 71.400 772.500 78.000 ;
        RECT 773.700 71.400 775.500 77.400 ;
        RECT 777.000 71.400 778.800 78.000 ;
        RECT 780.000 71.400 781.800 77.400 ;
        RECT 783.000 71.400 784.800 78.000 ;
        RECT 786.000 71.400 787.800 77.400 ;
        RECT 789.000 71.400 790.800 78.000 ;
        RECT 792.000 74.400 793.800 77.400 ;
        RECT 795.000 74.400 796.800 77.400 ;
        RECT 798.000 74.400 799.800 77.400 ;
        RECT 791.700 72.300 793.800 74.400 ;
        RECT 794.700 72.300 796.800 74.400 ;
        RECT 797.700 72.300 799.800 74.400 ;
        RECT 801.000 71.400 802.800 77.400 ;
        RECT 804.000 71.400 805.800 78.000 ;
        RECT 718.950 63.450 721.050 64.050 ;
        RECT 736.950 63.450 739.050 64.050 ;
        RECT 718.950 62.550 739.050 63.450 ;
        RECT 718.950 61.950 721.050 62.550 ;
        RECT 736.950 61.950 739.050 62.550 ;
        RECT 740.100 58.050 741.300 65.400 ;
        RECT 746.100 58.050 747.900 59.850 ;
        RECT 764.700 58.050 765.900 71.400 ;
        RECT 774.000 61.050 775.500 71.400 ;
        RECT 780.000 70.500 781.200 71.400 ;
        RECT 767.100 58.050 768.900 59.850 ;
        RECT 773.100 58.950 775.500 61.050 ;
        RECT 591.000 56.700 597.900 58.050 ;
        RECT 595.800 55.950 597.900 56.700 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 718.950 55.950 721.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 739.950 55.950 742.050 58.050 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 745.950 55.950 748.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 523.200 49.800 528.600 50.700 ;
        RECT 500.100 42.600 501.900 45.600 ;
        RECT 503.100 42.600 504.900 45.600 ;
        RECT 505.950 45.450 508.050 45.900 ;
        RECT 511.950 45.450 514.050 46.050 ;
        RECT 505.950 44.550 514.050 45.450 ;
        RECT 505.950 43.800 508.050 44.550 ;
        RECT 511.950 43.950 514.050 44.550 ;
        RECT 521.100 42.600 522.900 48.600 ;
        RECT 503.700 42.000 504.900 42.600 ;
        RECT 524.100 42.000 525.900 48.000 ;
        RECT 527.700 45.600 528.600 49.800 ;
        RECT 548.100 49.500 552.600 51.000 ;
        RECT 556.200 50.100 559.200 52.200 ;
        RECT 548.100 48.600 549.600 49.500 ;
        RECT 527.100 42.600 528.900 45.600 ;
        RECT 530.100 42.600 531.900 45.600 ;
        RECT 548.100 42.600 549.900 48.600 ;
        RECT 556.200 48.000 557.100 50.100 ;
        RECT 560.400 49.500 562.500 51.900 ;
        RECT 583.800 49.500 585.900 50.700 ;
        RECT 587.100 50.100 590.100 52.200 ;
        RECT 591.000 53.400 592.800 55.200 ;
        RECT 595.800 54.150 597.600 55.950 ;
        RECT 617.100 54.150 618.900 55.950 ;
        RECT 591.000 51.300 593.100 53.400 ;
        RECT 620.700 51.600 621.900 55.950 ;
        RECT 623.100 54.150 624.900 55.950 ;
        RECT 641.100 54.150 642.900 55.950 ;
        RECT 591.000 50.400 597.300 51.300 ;
        RECT 620.700 50.700 624.300 51.600 ;
        RECT 644.700 50.700 645.900 55.950 ;
        RECT 646.950 54.150 648.750 55.950 ;
        RECT 665.100 54.150 666.900 55.950 ;
        RECT 668.700 50.700 669.900 55.950 ;
        RECT 670.950 54.150 672.750 55.950 ;
        RECT 560.400 48.600 564.900 49.500 ;
        RECT 530.700 42.000 531.900 42.600 ;
        RECT 551.100 42.000 552.900 47.700 ;
        RECT 555.300 42.600 557.100 48.000 ;
        RECT 559.800 42.000 561.600 47.700 ;
        RECT 563.100 42.600 564.900 48.600 ;
        RECT 581.100 48.600 585.900 49.500 ;
        RECT 588.900 48.600 590.100 50.100 ;
        RECT 596.100 48.600 597.300 50.400 ;
        RECT 581.100 42.600 582.900 48.600 ;
        RECT 584.100 42.000 585.900 47.700 ;
        RECT 588.600 42.600 590.400 48.600 ;
        RECT 593.100 42.000 594.900 47.700 ;
        RECT 596.100 42.600 597.900 48.600 ;
        RECT 614.100 47.700 621.900 49.050 ;
        RECT 614.100 42.600 615.900 47.700 ;
        RECT 617.100 42.000 618.900 46.800 ;
        RECT 620.100 42.600 621.900 47.700 ;
        RECT 623.100 48.600 624.300 50.700 ;
        RECT 641.700 49.800 645.900 50.700 ;
        RECT 665.700 49.800 669.900 50.700 ;
        RECT 623.100 42.600 624.900 48.600 ;
        RECT 641.700 42.600 643.500 49.800 ;
        RECT 646.800 42.000 648.600 48.600 ;
        RECT 665.700 42.600 667.500 49.800 ;
        RECT 670.800 42.000 672.600 48.600 ;
        RECT 692.100 45.600 693.300 55.950 ;
        RECT 713.100 54.150 714.900 55.950 ;
        RECT 716.700 51.600 717.900 55.950 ;
        RECT 719.100 54.150 720.900 55.950 ;
        RECT 737.100 54.150 738.900 55.950 ;
        RECT 740.100 51.600 741.300 55.950 ;
        RECT 743.100 54.150 744.900 55.950 ;
        RECT 716.700 50.700 720.300 51.600 ;
        RECT 710.100 47.700 717.900 49.050 ;
        RECT 689.100 42.000 690.900 45.600 ;
        RECT 692.100 42.600 693.900 45.600 ;
        RECT 710.100 42.600 711.900 47.700 ;
        RECT 713.100 42.000 714.900 46.800 ;
        RECT 716.100 42.600 717.900 47.700 ;
        RECT 719.100 48.600 720.300 50.700 ;
        RECT 737.700 50.700 741.300 51.600 ;
        RECT 737.700 48.600 738.900 50.700 ;
        RECT 719.100 42.600 720.900 48.600 ;
        RECT 737.100 42.600 738.900 48.600 ;
        RECT 740.100 47.700 747.900 49.050 ;
        RECT 740.100 42.600 741.900 47.700 ;
        RECT 743.100 42.000 744.900 46.800 ;
        RECT 746.100 42.600 747.900 47.700 ;
        RECT 764.700 45.600 765.900 55.950 ;
        RECT 774.000 45.600 775.500 58.950 ;
        RECT 764.100 42.600 765.900 45.600 ;
        RECT 767.100 42.000 768.900 45.600 ;
        RECT 770.700 42.000 772.500 45.600 ;
        RECT 773.700 42.600 775.500 45.600 ;
        RECT 777.300 69.600 781.200 70.500 ;
        RECT 777.300 66.300 778.200 69.600 ;
        RECT 782.100 68.400 783.900 69.000 ;
        RECT 786.600 68.400 787.800 71.400 ;
        RECT 794.700 70.500 796.800 71.400 ;
        RECT 788.700 69.300 796.800 70.500 ;
        RECT 788.700 68.700 790.500 69.300 ;
        RECT 782.100 67.200 787.800 68.400 ;
        RECT 800.100 67.500 802.800 71.400 ;
        RECT 807.000 69.900 808.800 77.400 ;
        RECT 810.900 71.400 812.700 78.000 ;
        RECT 813.900 71.400 815.700 77.400 ;
        RECT 816.900 74.400 818.700 77.400 ;
        RECT 819.900 74.400 821.700 77.400 ;
        RECT 816.600 72.300 818.700 74.400 ;
        RECT 819.600 72.300 821.700 74.400 ;
        RECT 823.500 71.400 825.300 78.000 ;
        RECT 805.500 67.800 808.800 69.900 ;
        RECT 814.200 69.300 816.300 71.400 ;
        RECT 826.500 68.400 828.300 77.400 ;
        RECT 829.500 71.400 831.300 78.000 ;
        RECT 832.500 72.300 834.300 77.400 ;
        RECT 832.500 71.400 834.600 72.300 ;
        RECT 835.500 71.400 837.300 78.000 ;
        RECT 839.700 71.400 841.500 78.000 ;
        RECT 842.700 72.300 844.500 77.400 ;
        RECT 842.400 71.400 844.500 72.300 ;
        RECT 845.700 71.400 847.500 78.000 ;
        RECT 833.700 70.500 834.600 71.400 ;
        RECT 842.400 70.500 843.300 71.400 ;
        RECT 833.700 69.600 837.300 70.500 ;
        RECT 831.000 68.400 832.800 68.700 ;
        RECT 791.700 66.300 793.800 67.500 ;
        RECT 777.300 65.400 793.800 66.300 ;
        RECT 797.100 66.600 799.200 67.500 ;
        RECT 813.600 67.200 832.800 68.400 ;
        RECT 813.600 66.600 814.800 67.200 ;
        RECT 831.000 66.900 832.800 67.200 ;
        RECT 797.100 65.400 814.800 66.600 ;
        RECT 817.500 65.700 819.600 66.300 ;
        RECT 827.700 65.700 829.500 66.300 ;
        RECT 777.300 48.600 778.200 65.400 ;
        RECT 817.500 64.500 829.500 65.700 ;
        RECT 779.100 63.300 814.800 64.500 ;
        RECT 817.500 64.200 819.600 64.500 ;
        RECT 779.100 62.700 780.900 63.300 ;
        RECT 813.600 62.700 814.800 63.300 ;
        RECT 782.100 58.950 784.200 61.050 ;
        RECT 782.700 56.100 784.200 58.950 ;
        RECT 786.300 58.800 791.400 60.600 ;
        RECT 790.500 57.300 791.400 58.800 ;
        RECT 794.100 60.300 795.900 62.100 ;
        RECT 800.100 61.800 802.200 62.100 ;
        RECT 813.600 61.800 827.100 62.700 ;
        RECT 794.100 59.100 795.000 60.300 ;
        RECT 800.100 60.000 804.000 61.800 ;
        RECT 805.500 60.300 807.600 61.200 ;
        RECT 825.300 61.050 827.100 61.800 ;
        RECT 805.500 59.100 816.600 60.300 ;
        RECT 825.300 59.250 829.200 61.050 ;
        RECT 794.100 58.200 807.600 59.100 ;
        RECT 814.800 58.500 816.600 59.100 ;
        RECT 827.100 58.950 829.200 59.250 ;
        RECT 833.100 58.950 835.200 61.050 ;
        RECT 833.100 57.300 834.900 58.950 ;
        RECT 790.500 56.100 834.900 57.300 ;
        RECT 782.700 54.600 789.300 56.100 ;
        RECT 779.100 51.900 786.900 53.700 ;
        RECT 787.800 53.100 804.900 54.600 ;
        RECT 802.800 52.500 804.900 53.100 ;
        RECT 809.100 54.000 811.200 55.050 ;
        RECT 809.100 53.100 814.200 54.000 ;
        RECT 817.800 53.400 819.600 55.200 ;
        RECT 836.100 53.400 837.300 69.600 ;
        RECT 809.100 52.950 811.200 53.100 ;
        RECT 785.400 48.600 786.900 51.900 ;
        RECT 803.100 50.700 804.900 52.500 ;
        RECT 812.400 52.200 814.200 53.100 ;
        RECT 818.700 50.400 819.600 53.400 ;
        RECT 820.500 52.200 837.300 53.400 ;
        RECT 820.500 51.300 822.600 52.200 ;
        RECT 831.300 50.700 833.100 51.300 ;
        RECT 791.100 48.600 797.700 50.400 ;
        RECT 812.400 49.200 819.600 50.400 ;
        RECT 824.700 49.500 833.100 50.700 ;
        RECT 812.400 48.600 813.300 49.200 ;
        RECT 815.400 48.600 817.200 49.200 ;
        RECT 824.700 48.600 826.200 49.500 ;
        RECT 836.100 48.600 837.300 52.200 ;
        RECT 777.300 42.600 779.100 48.600 ;
        RECT 782.700 42.000 784.500 48.600 ;
        RECT 785.400 47.400 789.600 48.600 ;
        RECT 787.800 42.600 789.600 47.400 ;
        RECT 791.700 45.600 793.800 47.700 ;
        RECT 794.700 45.600 796.800 47.700 ;
        RECT 797.700 45.600 799.800 47.700 ;
        RECT 800.700 45.600 802.800 47.700 ;
        RECT 806.100 46.500 808.800 48.600 ;
        RECT 810.600 47.400 813.300 48.600 ;
        RECT 810.600 46.500 812.400 47.400 ;
        RECT 792.000 42.600 793.800 45.600 ;
        RECT 795.000 42.600 796.800 45.600 ;
        RECT 798.000 42.600 799.800 45.600 ;
        RECT 801.000 42.600 802.800 45.600 ;
        RECT 804.000 42.000 805.800 45.600 ;
        RECT 807.000 42.600 808.800 46.500 ;
        RECT 814.200 45.600 816.300 47.700 ;
        RECT 817.200 45.600 819.300 47.700 ;
        RECT 820.200 45.600 822.300 47.700 ;
        RECT 811.500 42.000 813.300 45.600 ;
        RECT 814.500 42.600 816.300 45.600 ;
        RECT 817.500 42.600 819.300 45.600 ;
        RECT 820.500 42.600 822.300 45.600 ;
        RECT 824.700 42.600 826.500 48.600 ;
        RECT 830.100 42.000 831.900 48.600 ;
        RECT 835.500 42.600 837.300 48.600 ;
        RECT 839.700 69.600 843.300 70.500 ;
        RECT 839.700 53.400 840.900 69.600 ;
        RECT 844.200 68.400 846.000 68.700 ;
        RECT 848.700 68.400 850.500 77.400 ;
        RECT 851.700 71.400 853.500 78.000 ;
        RECT 855.300 74.400 857.100 77.400 ;
        RECT 858.300 74.400 860.100 77.400 ;
        RECT 855.300 72.300 857.400 74.400 ;
        RECT 858.300 72.300 860.400 74.400 ;
        RECT 861.300 71.400 863.100 77.400 ;
        RECT 864.300 71.400 866.100 78.000 ;
        RECT 860.700 69.300 862.800 71.400 ;
        RECT 868.200 69.900 870.000 77.400 ;
        RECT 871.200 71.400 873.000 78.000 ;
        RECT 874.200 71.400 876.000 77.400 ;
        RECT 877.200 74.400 879.000 77.400 ;
        RECT 880.200 74.400 882.000 77.400 ;
        RECT 883.200 74.400 885.000 77.400 ;
        RECT 877.200 72.300 879.300 74.400 ;
        RECT 880.200 72.300 882.300 74.400 ;
        RECT 883.200 72.300 885.300 74.400 ;
        RECT 886.200 71.400 888.000 78.000 ;
        RECT 889.200 71.400 891.000 77.400 ;
        RECT 892.200 71.400 894.000 78.000 ;
        RECT 895.200 71.400 897.000 77.400 ;
        RECT 898.200 71.400 900.000 78.000 ;
        RECT 901.500 71.400 903.300 77.400 ;
        RECT 904.500 71.400 906.300 78.000 ;
        RECT 844.200 67.200 863.400 68.400 ;
        RECT 868.200 67.800 871.500 69.900 ;
        RECT 874.200 67.500 876.900 71.400 ;
        RECT 880.200 70.500 882.300 71.400 ;
        RECT 880.200 69.300 888.300 70.500 ;
        RECT 886.500 68.700 888.300 69.300 ;
        RECT 889.200 68.400 890.400 71.400 ;
        RECT 895.800 70.500 897.000 71.400 ;
        RECT 895.800 69.600 899.700 70.500 ;
        RECT 893.100 68.400 894.900 69.000 ;
        RECT 844.200 66.900 846.000 67.200 ;
        RECT 862.200 66.600 863.400 67.200 ;
        RECT 877.800 66.600 879.900 67.500 ;
        RECT 847.500 65.700 849.300 66.300 ;
        RECT 857.400 65.700 859.500 66.300 ;
        RECT 847.500 64.500 859.500 65.700 ;
        RECT 862.200 65.400 879.900 66.600 ;
        RECT 883.200 66.300 885.300 67.500 ;
        RECT 889.200 67.200 894.900 68.400 ;
        RECT 898.800 66.300 899.700 69.600 ;
        RECT 883.200 65.400 899.700 66.300 ;
        RECT 857.400 64.200 859.500 64.500 ;
        RECT 862.200 63.300 897.900 64.500 ;
        RECT 862.200 62.700 863.400 63.300 ;
        RECT 896.100 62.700 897.900 63.300 ;
        RECT 849.900 61.800 863.400 62.700 ;
        RECT 874.800 61.800 876.900 62.100 ;
        RECT 849.900 61.050 851.700 61.800 ;
        RECT 841.800 58.950 843.900 61.050 ;
        RECT 847.800 59.250 851.700 61.050 ;
        RECT 869.400 60.300 871.500 61.200 ;
        RECT 847.800 58.950 849.900 59.250 ;
        RECT 860.400 59.100 871.500 60.300 ;
        RECT 873.000 60.000 876.900 61.800 ;
        RECT 881.100 60.300 882.900 62.100 ;
        RECT 882.000 59.100 882.900 60.300 ;
        RECT 842.100 57.300 843.900 58.950 ;
        RECT 860.400 58.500 862.200 59.100 ;
        RECT 869.400 58.200 882.900 59.100 ;
        RECT 885.600 58.800 890.700 60.600 ;
        RECT 892.800 58.950 894.900 61.050 ;
        RECT 885.600 57.300 886.500 58.800 ;
        RECT 842.100 56.100 886.500 57.300 ;
        RECT 892.800 56.100 894.300 58.950 ;
        RECT 857.400 53.400 859.200 55.200 ;
        RECT 865.800 54.000 867.900 55.050 ;
        RECT 887.700 54.600 894.300 56.100 ;
        RECT 839.700 52.200 856.500 53.400 ;
        RECT 839.700 48.600 840.900 52.200 ;
        RECT 854.400 51.300 856.500 52.200 ;
        RECT 843.900 50.700 845.700 51.300 ;
        RECT 843.900 49.500 852.300 50.700 ;
        RECT 850.800 48.600 852.300 49.500 ;
        RECT 857.400 50.400 858.300 53.400 ;
        RECT 862.800 53.100 867.900 54.000 ;
        RECT 862.800 52.200 864.600 53.100 ;
        RECT 865.800 52.950 867.900 53.100 ;
        RECT 872.100 53.100 889.200 54.600 ;
        RECT 872.100 52.500 874.200 53.100 ;
        RECT 872.100 50.700 873.900 52.500 ;
        RECT 890.100 51.900 897.900 53.700 ;
        RECT 857.400 49.200 864.600 50.400 ;
        RECT 859.800 48.600 861.600 49.200 ;
        RECT 863.700 48.600 864.600 49.200 ;
        RECT 879.300 48.600 885.900 50.400 ;
        RECT 890.100 48.600 891.600 51.900 ;
        RECT 898.800 48.600 899.700 65.400 ;
        RECT 839.700 42.600 841.500 48.600 ;
        RECT 845.100 42.000 846.900 48.600 ;
        RECT 850.500 42.600 852.300 48.600 ;
        RECT 854.700 45.600 856.800 47.700 ;
        RECT 857.700 45.600 859.800 47.700 ;
        RECT 860.700 45.600 862.800 47.700 ;
        RECT 863.700 47.400 866.400 48.600 ;
        RECT 864.600 46.500 866.400 47.400 ;
        RECT 868.200 46.500 870.900 48.600 ;
        RECT 854.700 42.600 856.500 45.600 ;
        RECT 857.700 42.600 859.500 45.600 ;
        RECT 860.700 42.600 862.500 45.600 ;
        RECT 863.700 42.000 865.500 45.600 ;
        RECT 868.200 42.600 870.000 46.500 ;
        RECT 874.200 45.600 876.300 47.700 ;
        RECT 877.200 45.600 879.300 47.700 ;
        RECT 880.200 45.600 882.300 47.700 ;
        RECT 883.200 45.600 885.300 47.700 ;
        RECT 887.400 47.400 891.600 48.600 ;
        RECT 871.200 42.000 873.000 45.600 ;
        RECT 874.200 42.600 876.000 45.600 ;
        RECT 877.200 42.600 879.000 45.600 ;
        RECT 880.200 42.600 882.000 45.600 ;
        RECT 883.200 42.600 885.000 45.600 ;
        RECT 887.400 42.600 889.200 47.400 ;
        RECT 892.500 42.000 894.300 48.600 ;
        RECT 897.900 42.600 899.700 48.600 ;
        RECT 901.500 61.050 903.000 71.400 ;
        RECT 923.400 65.400 925.200 78.000 ;
        RECT 928.500 66.900 930.300 77.400 ;
        RECT 931.500 71.400 933.300 78.000 ;
        RECT 950.100 71.400 951.900 78.000 ;
        RECT 953.100 71.400 954.900 77.400 ;
        RECT 956.100 72.000 957.900 78.000 ;
        RECT 953.400 71.100 954.900 71.400 ;
        RECT 959.100 71.400 960.900 77.400 ;
        RECT 959.100 71.100 960.000 71.400 ;
        RECT 953.400 70.200 960.000 71.100 ;
        RECT 931.200 68.100 933.000 69.900 ;
        RECT 928.500 65.400 930.900 66.900 ;
        RECT 901.500 58.950 903.900 61.050 ;
        RECT 901.500 45.600 903.000 58.950 ;
        RECT 923.100 58.050 924.900 59.850 ;
        RECT 929.700 58.050 930.900 65.400 ;
        RECT 953.100 58.050 954.900 59.850 ;
        RECT 959.100 58.050 960.000 70.200 ;
        RECT 978.600 66.900 980.400 77.400 ;
        RECT 978.000 65.400 980.400 66.900 ;
        RECT 981.600 65.400 983.400 78.000 ;
        RECT 986.100 65.400 987.900 77.400 ;
        RECT 1004.100 71.400 1005.900 78.000 ;
        RECT 1007.100 71.400 1008.900 77.400 ;
        RECT 1010.100 71.400 1011.900 78.000 ;
        RECT 1028.700 71.400 1030.500 78.000 ;
        RECT 978.000 58.050 979.200 65.400 ;
        RECT 986.700 63.900 987.900 65.400 ;
        RECT 980.100 62.700 987.900 63.900 ;
        RECT 980.100 62.100 981.900 62.700 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 928.950 55.950 931.050 58.050 ;
        RECT 931.950 55.950 934.050 58.050 ;
        RECT 949.950 55.950 952.050 58.050 ;
        RECT 952.950 55.950 955.050 58.050 ;
        RECT 955.950 55.950 958.050 58.050 ;
        RECT 958.950 55.950 961.050 58.050 ;
        RECT 977.100 55.950 979.200 58.050 ;
        RECT 926.100 54.150 927.900 55.950 ;
        RECT 929.700 51.600 930.900 55.950 ;
        RECT 932.100 54.150 933.900 55.950 ;
        RECT 950.100 54.150 951.900 55.950 ;
        RECT 956.100 54.150 957.900 55.950 ;
        RECT 959.100 52.200 960.000 55.950 ;
        RECT 929.700 50.700 933.300 51.600 ;
        RECT 923.100 47.700 930.900 49.050 ;
        RECT 901.500 42.600 903.300 45.600 ;
        RECT 904.500 42.000 906.300 45.600 ;
        RECT 923.100 42.600 924.900 47.700 ;
        RECT 926.100 42.000 927.900 46.800 ;
        RECT 929.100 42.600 930.900 47.700 ;
        RECT 932.100 48.600 933.300 50.700 ;
        RECT 932.100 42.600 933.900 48.600 ;
        RECT 950.100 42.000 951.900 51.600 ;
        RECT 956.700 51.000 960.000 52.200 ;
        RECT 956.700 42.600 958.500 51.000 ;
        RECT 977.100 48.600 978.000 55.950 ;
        RECT 980.400 51.600 981.300 62.100 ;
        RECT 982.200 58.050 984.000 59.850 ;
        RECT 1007.700 58.050 1008.900 71.400 ;
        RECT 1029.000 68.100 1030.800 69.900 ;
        RECT 1031.700 66.900 1033.500 77.400 ;
        RECT 1031.100 65.400 1033.500 66.900 ;
        RECT 1036.800 65.400 1038.600 78.000 ;
        RECT 1031.100 58.050 1032.300 65.400 ;
        RECT 1037.100 58.050 1038.900 59.850 ;
        RECT 982.500 55.950 984.600 58.050 ;
        RECT 985.800 55.950 987.900 58.050 ;
        RECT 1003.950 55.950 1006.050 58.050 ;
        RECT 1006.950 55.950 1009.050 58.050 ;
        RECT 1009.950 55.950 1012.050 58.050 ;
        RECT 1027.950 55.950 1030.050 58.050 ;
        RECT 1030.950 55.950 1033.050 58.050 ;
        RECT 1033.950 55.950 1036.050 58.050 ;
        RECT 1036.950 55.950 1039.050 58.050 ;
        RECT 985.800 54.150 987.600 55.950 ;
        RECT 1004.100 54.150 1005.900 55.950 ;
        RECT 979.200 50.700 981.300 51.600 ;
        RECT 1007.700 50.700 1008.900 55.950 ;
        RECT 1009.950 54.150 1011.750 55.950 ;
        RECT 1028.100 54.150 1029.900 55.950 ;
        RECT 1031.100 51.600 1032.300 55.950 ;
        RECT 1034.100 54.150 1035.900 55.950 ;
        RECT 979.200 49.800 984.600 50.700 ;
        RECT 977.100 42.600 978.900 48.600 ;
        RECT 980.100 42.000 981.900 48.000 ;
        RECT 983.700 45.600 984.600 49.800 ;
        RECT 1004.700 49.800 1008.900 50.700 ;
        RECT 1028.700 50.700 1032.300 51.600 ;
        RECT 983.100 42.600 984.900 45.600 ;
        RECT 986.100 42.600 987.900 45.600 ;
        RECT 1004.700 42.600 1006.500 49.800 ;
        RECT 1028.700 48.600 1029.900 50.700 ;
        RECT 986.700 42.000 987.900 42.600 ;
        RECT 1009.800 42.000 1011.600 48.600 ;
        RECT 1028.100 42.600 1029.900 48.600 ;
        RECT 1031.100 47.700 1038.900 49.050 ;
        RECT 1031.100 42.600 1032.900 47.700 ;
        RECT 1034.100 42.000 1035.900 46.800 ;
        RECT 1037.100 42.600 1038.900 47.700 ;
        RECT 17.100 32.400 18.900 38.400 ;
        RECT 20.100 32.400 21.900 39.000 ;
        RECT 23.100 35.400 24.900 38.400 ;
        RECT 17.100 25.050 18.300 32.400 ;
        RECT 23.700 31.500 24.900 35.400 ;
        RECT 19.200 30.600 24.900 31.500 ;
        RECT 41.100 32.400 42.900 38.400 ;
        RECT 44.100 32.400 45.900 39.000 ;
        RECT 47.100 35.400 48.900 38.400 ;
        RECT 19.200 29.700 21.000 30.600 ;
        RECT 17.100 22.950 19.200 25.050 ;
        RECT 17.100 15.600 18.300 22.950 ;
        RECT 20.100 18.300 21.000 29.700 ;
        RECT 41.100 25.050 42.300 32.400 ;
        RECT 47.700 31.500 48.900 35.400 ;
        RECT 43.200 30.600 48.900 31.500 ;
        RECT 65.100 35.400 66.900 38.400 ;
        RECT 65.100 31.500 66.300 35.400 ;
        RECT 68.100 32.400 69.900 39.000 ;
        RECT 71.100 32.400 72.900 38.400 ;
        RECT 65.100 30.600 70.800 31.500 ;
        RECT 43.200 29.700 45.000 30.600 ;
        RECT 22.500 22.950 24.600 25.050 ;
        RECT 22.800 21.150 24.600 22.950 ;
        RECT 41.100 22.950 43.200 25.050 ;
        RECT 19.200 17.400 21.000 18.300 ;
        RECT 19.200 16.500 24.900 17.400 ;
        RECT 17.100 3.600 18.900 15.600 ;
        RECT 20.100 3.000 21.900 13.800 ;
        RECT 23.700 9.600 24.900 16.500 ;
        RECT 23.100 3.600 24.900 9.600 ;
        RECT 41.100 15.600 42.300 22.950 ;
        RECT 44.100 18.300 45.000 29.700 ;
        RECT 69.000 29.700 70.800 30.600 ;
        RECT 46.500 22.950 48.600 25.050 ;
        RECT 46.800 21.150 48.600 22.950 ;
        RECT 65.400 22.950 67.500 25.050 ;
        RECT 65.400 21.150 67.200 22.950 ;
        RECT 43.200 17.400 45.000 18.300 ;
        RECT 69.000 18.300 69.900 29.700 ;
        RECT 71.700 25.050 72.900 32.400 ;
        RECT 89.100 33.300 90.900 38.400 ;
        RECT 92.100 34.200 93.900 39.000 ;
        RECT 95.100 33.300 96.900 38.400 ;
        RECT 89.100 31.950 96.900 33.300 ;
        RECT 98.100 32.400 99.900 38.400 ;
        RECT 117.600 34.200 119.400 38.400 ;
        RECT 116.700 32.400 119.400 34.200 ;
        RECT 120.600 32.400 122.400 39.000 ;
        RECT 98.100 30.300 99.300 32.400 ;
        RECT 95.700 29.400 99.300 30.300 ;
        RECT 92.100 25.050 93.900 26.850 ;
        RECT 95.700 25.050 96.900 29.400 ;
        RECT 98.100 25.050 99.900 26.850 ;
        RECT 116.700 25.050 117.600 32.400 ;
        RECT 118.500 30.600 120.300 31.500 ;
        RECT 125.100 30.600 126.900 38.400 ;
        RECT 118.500 29.700 126.900 30.600 ;
        RECT 143.700 31.200 145.500 38.400 ;
        RECT 148.800 32.400 150.600 39.000 ;
        RECT 167.100 32.400 168.900 38.400 ;
        RECT 170.100 32.400 171.900 39.000 ;
        RECT 173.100 35.400 174.900 38.400 ;
        RECT 143.700 30.300 147.900 31.200 ;
        RECT 70.800 22.950 72.900 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 97.950 22.950 100.050 25.050 ;
        RECT 116.100 22.950 118.200 25.050 ;
        RECT 119.400 22.950 121.500 25.050 ;
        RECT 69.000 17.400 70.800 18.300 ;
        RECT 43.200 16.500 48.900 17.400 ;
        RECT 41.100 3.600 42.900 15.600 ;
        RECT 44.100 3.000 45.900 13.800 ;
        RECT 47.700 9.600 48.900 16.500 ;
        RECT 47.100 3.600 48.900 9.600 ;
        RECT 65.100 16.500 70.800 17.400 ;
        RECT 65.100 9.600 66.300 16.500 ;
        RECT 71.700 15.600 72.900 22.950 ;
        RECT 89.100 21.150 90.900 22.950 ;
        RECT 95.700 15.600 96.900 22.950 ;
        RECT 116.700 15.600 117.600 22.950 ;
        RECT 120.000 21.150 121.800 22.950 ;
        RECT 65.100 3.600 66.900 9.600 ;
        RECT 68.100 3.000 69.900 13.800 ;
        RECT 71.100 3.600 72.900 15.600 ;
        RECT 89.400 3.000 91.200 15.600 ;
        RECT 94.500 14.100 96.900 15.600 ;
        RECT 94.500 3.600 96.300 14.100 ;
        RECT 97.200 11.100 99.000 12.900 ;
        RECT 97.500 3.000 99.300 9.600 ;
        RECT 116.100 3.600 117.900 15.600 ;
        RECT 119.100 3.000 120.900 15.000 ;
        RECT 123.000 9.600 123.900 29.700 ;
        RECT 124.950 25.050 126.750 26.850 ;
        RECT 143.100 25.050 144.900 26.850 ;
        RECT 146.700 25.050 147.900 30.300 ;
        RECT 148.950 25.050 150.750 26.850 ;
        RECT 167.100 25.050 168.300 32.400 ;
        RECT 173.700 31.500 174.900 35.400 ;
        RECT 169.200 30.600 174.900 31.500 ;
        RECT 191.100 35.400 192.900 38.400 ;
        RECT 191.100 31.500 192.300 35.400 ;
        RECT 194.100 32.400 195.900 39.000 ;
        RECT 197.100 32.400 198.900 38.400 ;
        RECT 215.100 35.400 216.900 38.400 ;
        RECT 218.100 35.400 219.900 39.000 ;
        RECT 236.100 35.400 237.900 38.400 ;
        RECT 191.100 30.600 196.800 31.500 ;
        RECT 169.200 29.700 171.000 30.600 ;
        RECT 124.800 22.950 126.900 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 167.100 22.950 169.200 25.050 ;
        RECT 146.700 9.600 147.900 22.950 ;
        RECT 167.100 15.600 168.300 22.950 ;
        RECT 170.100 18.300 171.000 29.700 ;
        RECT 195.000 29.700 196.800 30.600 ;
        RECT 172.500 22.950 174.600 25.050 ;
        RECT 172.800 21.150 174.600 22.950 ;
        RECT 191.400 22.950 193.500 25.050 ;
        RECT 191.400 21.150 193.200 22.950 ;
        RECT 169.200 17.400 171.000 18.300 ;
        RECT 195.000 18.300 195.900 29.700 ;
        RECT 197.700 25.050 198.900 32.400 ;
        RECT 215.700 25.050 216.900 35.400 ;
        RECT 236.100 31.500 237.300 35.400 ;
        RECT 239.100 32.400 240.900 39.000 ;
        RECT 242.100 32.400 243.900 38.400 ;
        RECT 245.700 35.400 247.500 39.000 ;
        RECT 248.700 35.400 250.500 38.400 ;
        RECT 236.100 30.600 241.800 31.500 ;
        RECT 240.000 29.700 241.800 30.600 ;
        RECT 196.800 22.950 198.900 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 236.400 22.950 238.500 25.050 ;
        RECT 195.000 17.400 196.800 18.300 ;
        RECT 169.200 16.500 174.900 17.400 ;
        RECT 122.100 3.600 123.900 9.600 ;
        RECT 125.100 3.000 126.900 9.600 ;
        RECT 143.100 3.000 144.900 9.600 ;
        RECT 146.100 3.600 147.900 9.600 ;
        RECT 149.100 3.000 150.900 9.600 ;
        RECT 167.100 3.600 168.900 15.600 ;
        RECT 170.100 3.000 171.900 13.800 ;
        RECT 173.700 9.600 174.900 16.500 ;
        RECT 173.100 3.600 174.900 9.600 ;
        RECT 191.100 16.500 196.800 17.400 ;
        RECT 191.100 9.600 192.300 16.500 ;
        RECT 197.700 15.600 198.900 22.950 ;
        RECT 191.100 3.600 192.900 9.600 ;
        RECT 194.100 3.000 195.900 13.800 ;
        RECT 197.100 3.600 198.900 15.600 ;
        RECT 215.700 9.600 216.900 22.950 ;
        RECT 218.100 21.150 219.900 22.950 ;
        RECT 236.400 21.150 238.200 22.950 ;
        RECT 240.000 18.300 240.900 29.700 ;
        RECT 242.700 25.050 243.900 32.400 ;
        RECT 241.800 22.950 243.900 25.050 ;
        RECT 240.000 17.400 241.800 18.300 ;
        RECT 236.100 16.500 241.800 17.400 ;
        RECT 236.100 9.600 237.300 16.500 ;
        RECT 242.700 15.600 243.900 22.950 ;
        RECT 249.000 22.050 250.500 35.400 ;
        RECT 248.100 19.950 250.500 22.050 ;
        RECT 215.100 3.600 216.900 9.600 ;
        RECT 218.100 3.000 219.900 9.600 ;
        RECT 236.100 3.600 237.900 9.600 ;
        RECT 239.100 3.000 240.900 13.800 ;
        RECT 242.100 3.600 243.900 15.600 ;
        RECT 249.000 9.600 250.500 19.950 ;
        RECT 252.300 32.400 254.100 38.400 ;
        RECT 257.700 32.400 259.500 39.000 ;
        RECT 262.800 33.600 264.600 38.400 ;
        RECT 267.000 35.400 268.800 38.400 ;
        RECT 270.000 35.400 271.800 38.400 ;
        RECT 273.000 35.400 274.800 38.400 ;
        RECT 276.000 35.400 277.800 38.400 ;
        RECT 279.000 35.400 280.800 39.000 ;
        RECT 260.400 32.400 264.600 33.600 ;
        RECT 266.700 33.300 268.800 35.400 ;
        RECT 269.700 33.300 271.800 35.400 ;
        RECT 272.700 33.300 274.800 35.400 ;
        RECT 275.700 33.300 277.800 35.400 ;
        RECT 282.000 34.500 283.800 38.400 ;
        RECT 286.500 35.400 288.300 39.000 ;
        RECT 289.500 35.400 291.300 38.400 ;
        RECT 292.500 35.400 294.300 38.400 ;
        RECT 295.500 35.400 297.300 38.400 ;
        RECT 281.100 32.400 283.800 34.500 ;
        RECT 285.600 33.600 287.400 34.500 ;
        RECT 285.600 32.400 288.300 33.600 ;
        RECT 289.200 33.300 291.300 35.400 ;
        RECT 292.200 33.300 294.300 35.400 ;
        RECT 295.200 33.300 297.300 35.400 ;
        RECT 299.700 32.400 301.500 38.400 ;
        RECT 305.100 32.400 306.900 39.000 ;
        RECT 310.500 32.400 312.300 38.400 ;
        RECT 252.300 15.600 253.200 32.400 ;
        RECT 260.400 29.100 261.900 32.400 ;
        RECT 266.100 30.600 272.700 32.400 ;
        RECT 287.400 31.800 288.300 32.400 ;
        RECT 290.400 31.800 292.200 32.400 ;
        RECT 287.400 30.600 294.600 31.800 ;
        RECT 254.100 27.300 261.900 29.100 ;
        RECT 278.100 28.500 279.900 30.300 ;
        RECT 277.800 27.900 279.900 28.500 ;
        RECT 262.800 26.400 279.900 27.900 ;
        RECT 284.100 27.900 286.200 28.050 ;
        RECT 287.400 27.900 289.200 28.800 ;
        RECT 284.100 27.000 289.200 27.900 ;
        RECT 293.700 27.600 294.600 30.600 ;
        RECT 299.700 31.500 301.200 32.400 ;
        RECT 299.700 30.300 308.100 31.500 ;
        RECT 306.300 29.700 308.100 30.300 ;
        RECT 295.500 28.800 297.600 29.700 ;
        RECT 311.100 28.800 312.300 32.400 ;
        RECT 295.500 27.600 312.300 28.800 ;
        RECT 257.700 24.900 264.300 26.400 ;
        RECT 284.100 25.950 286.200 27.000 ;
        RECT 292.800 25.800 294.600 27.600 ;
        RECT 257.700 22.050 259.200 24.900 ;
        RECT 265.500 23.700 309.900 24.900 ;
        RECT 265.500 22.200 266.400 23.700 ;
        RECT 257.100 19.950 259.200 22.050 ;
        RECT 261.300 20.400 266.400 22.200 ;
        RECT 269.100 21.900 282.600 22.800 ;
        RECT 289.800 21.900 291.600 22.500 ;
        RECT 308.100 22.050 309.900 23.700 ;
        RECT 269.100 20.700 270.000 21.900 ;
        RECT 269.100 18.900 270.900 20.700 ;
        RECT 275.100 19.200 279.000 21.000 ;
        RECT 280.500 20.700 291.600 21.900 ;
        RECT 302.100 21.750 304.200 22.050 ;
        RECT 280.500 19.800 282.600 20.700 ;
        RECT 300.300 19.950 304.200 21.750 ;
        RECT 308.100 19.950 310.200 22.050 ;
        RECT 300.300 19.200 302.100 19.950 ;
        RECT 275.100 18.900 277.200 19.200 ;
        RECT 288.600 18.300 302.100 19.200 ;
        RECT 254.100 17.700 255.900 18.300 ;
        RECT 288.600 17.700 289.800 18.300 ;
        RECT 254.100 16.500 289.800 17.700 ;
        RECT 292.500 16.500 294.600 16.800 ;
        RECT 252.300 14.700 268.800 15.600 ;
        RECT 252.300 11.400 253.200 14.700 ;
        RECT 257.100 12.600 262.800 13.800 ;
        RECT 266.700 13.500 268.800 14.700 ;
        RECT 272.100 14.400 289.800 15.600 ;
        RECT 292.500 15.300 304.500 16.500 ;
        RECT 292.500 14.700 294.600 15.300 ;
        RECT 302.700 14.700 304.500 15.300 ;
        RECT 272.100 13.500 274.200 14.400 ;
        RECT 288.600 13.800 289.800 14.400 ;
        RECT 306.000 13.800 307.800 14.100 ;
        RECT 257.100 12.000 258.900 12.600 ;
        RECT 252.300 10.500 256.200 11.400 ;
        RECT 255.000 9.600 256.200 10.500 ;
        RECT 261.600 9.600 262.800 12.600 ;
        RECT 263.700 11.700 265.500 12.300 ;
        RECT 263.700 10.500 271.800 11.700 ;
        RECT 269.700 9.600 271.800 10.500 ;
        RECT 275.100 9.600 277.800 13.500 ;
        RECT 280.500 11.100 283.800 13.200 ;
        RECT 288.600 12.600 307.800 13.800 ;
        RECT 245.700 3.000 247.500 9.600 ;
        RECT 248.700 3.600 250.500 9.600 ;
        RECT 252.000 3.000 253.800 9.600 ;
        RECT 255.000 3.600 256.800 9.600 ;
        RECT 258.000 3.000 259.800 9.600 ;
        RECT 261.000 3.600 262.800 9.600 ;
        RECT 264.000 3.000 265.800 9.600 ;
        RECT 266.700 6.600 268.800 8.700 ;
        RECT 269.700 6.600 271.800 8.700 ;
        RECT 272.700 6.600 274.800 8.700 ;
        RECT 267.000 3.600 268.800 6.600 ;
        RECT 270.000 3.600 271.800 6.600 ;
        RECT 273.000 3.600 274.800 6.600 ;
        RECT 276.000 3.600 277.800 9.600 ;
        RECT 279.000 3.000 280.800 9.600 ;
        RECT 282.000 3.600 283.800 11.100 ;
        RECT 289.200 9.600 291.300 11.700 ;
        RECT 285.900 3.000 287.700 9.600 ;
        RECT 288.900 3.600 290.700 9.600 ;
        RECT 291.600 6.600 293.700 8.700 ;
        RECT 294.600 6.600 296.700 8.700 ;
        RECT 291.900 3.600 293.700 6.600 ;
        RECT 294.900 3.600 296.700 6.600 ;
        RECT 298.500 3.000 300.300 9.600 ;
        RECT 301.500 3.600 303.300 12.600 ;
        RECT 306.000 12.300 307.800 12.600 ;
        RECT 311.100 11.400 312.300 27.600 ;
        RECT 308.700 10.500 312.300 11.400 ;
        RECT 314.700 32.400 316.500 38.400 ;
        RECT 320.100 32.400 321.900 39.000 ;
        RECT 325.500 32.400 327.300 38.400 ;
        RECT 329.700 35.400 331.500 38.400 ;
        RECT 332.700 35.400 334.500 38.400 ;
        RECT 335.700 35.400 337.500 38.400 ;
        RECT 338.700 35.400 340.500 39.000 ;
        RECT 329.700 33.300 331.800 35.400 ;
        RECT 332.700 33.300 334.800 35.400 ;
        RECT 335.700 33.300 337.800 35.400 ;
        RECT 343.200 34.500 345.000 38.400 ;
        RECT 346.200 35.400 348.000 39.000 ;
        RECT 349.200 35.400 351.000 38.400 ;
        RECT 352.200 35.400 354.000 38.400 ;
        RECT 355.200 35.400 357.000 38.400 ;
        RECT 358.200 35.400 360.000 38.400 ;
        RECT 339.600 33.600 341.400 34.500 ;
        RECT 338.700 32.400 341.400 33.600 ;
        RECT 343.200 32.400 345.900 34.500 ;
        RECT 349.200 33.300 351.300 35.400 ;
        RECT 352.200 33.300 354.300 35.400 ;
        RECT 355.200 33.300 357.300 35.400 ;
        RECT 358.200 33.300 360.300 35.400 ;
        RECT 362.400 33.600 364.200 38.400 ;
        RECT 362.400 32.400 366.600 33.600 ;
        RECT 367.500 32.400 369.300 39.000 ;
        RECT 372.900 32.400 374.700 38.400 ;
        RECT 314.700 28.800 315.900 32.400 ;
        RECT 325.800 31.500 327.300 32.400 ;
        RECT 334.800 31.800 336.600 32.400 ;
        RECT 338.700 31.800 339.600 32.400 ;
        RECT 318.900 30.300 327.300 31.500 ;
        RECT 332.400 30.600 339.600 31.800 ;
        RECT 354.300 30.600 360.900 32.400 ;
        RECT 318.900 29.700 320.700 30.300 ;
        RECT 329.400 28.800 331.500 29.700 ;
        RECT 314.700 27.600 331.500 28.800 ;
        RECT 332.400 27.600 333.300 30.600 ;
        RECT 337.800 27.900 339.600 28.800 ;
        RECT 347.100 28.500 348.900 30.300 ;
        RECT 365.100 29.100 366.600 32.400 ;
        RECT 340.800 27.900 342.900 28.050 ;
        RECT 314.700 11.400 315.900 27.600 ;
        RECT 332.400 25.800 334.200 27.600 ;
        RECT 337.800 27.000 342.900 27.900 ;
        RECT 340.800 25.950 342.900 27.000 ;
        RECT 347.100 27.900 349.200 28.500 ;
        RECT 347.100 26.400 364.200 27.900 ;
        RECT 365.100 27.300 372.900 29.100 ;
        RECT 362.700 24.900 369.300 26.400 ;
        RECT 317.100 23.700 361.500 24.900 ;
        RECT 317.100 22.050 318.900 23.700 ;
        RECT 316.800 19.950 318.900 22.050 ;
        RECT 322.800 21.750 324.900 22.050 ;
        RECT 335.400 21.900 337.200 22.500 ;
        RECT 344.400 21.900 357.900 22.800 ;
        RECT 322.800 19.950 326.700 21.750 ;
        RECT 335.400 20.700 346.500 21.900 ;
        RECT 324.900 19.200 326.700 19.950 ;
        RECT 344.400 19.800 346.500 20.700 ;
        RECT 348.000 19.200 351.900 21.000 ;
        RECT 357.000 20.700 357.900 21.900 ;
        RECT 324.900 18.300 338.400 19.200 ;
        RECT 349.800 18.900 351.900 19.200 ;
        RECT 356.100 18.900 357.900 20.700 ;
        RECT 360.600 22.200 361.500 23.700 ;
        RECT 360.600 20.400 365.700 22.200 ;
        RECT 367.800 22.050 369.300 24.900 ;
        RECT 367.800 19.950 369.900 22.050 ;
        RECT 337.200 17.700 338.400 18.300 ;
        RECT 371.100 17.700 372.900 18.300 ;
        RECT 332.400 16.500 334.500 16.800 ;
        RECT 337.200 16.500 372.900 17.700 ;
        RECT 322.500 15.300 334.500 16.500 ;
        RECT 373.800 15.600 374.700 32.400 ;
        RECT 322.500 14.700 324.300 15.300 ;
        RECT 332.400 14.700 334.500 15.300 ;
        RECT 337.200 14.400 354.900 15.600 ;
        RECT 319.200 13.800 321.000 14.100 ;
        RECT 337.200 13.800 338.400 14.400 ;
        RECT 319.200 12.600 338.400 13.800 ;
        RECT 352.800 13.500 354.900 14.400 ;
        RECT 358.200 14.700 374.700 15.600 ;
        RECT 358.200 13.500 360.300 14.700 ;
        RECT 319.200 12.300 321.000 12.600 ;
        RECT 314.700 10.500 318.300 11.400 ;
        RECT 308.700 9.600 309.600 10.500 ;
        RECT 317.400 9.600 318.300 10.500 ;
        RECT 304.500 3.000 306.300 9.600 ;
        RECT 307.500 8.700 309.600 9.600 ;
        RECT 307.500 3.600 309.300 8.700 ;
        RECT 310.500 3.000 312.300 9.600 ;
        RECT 314.700 3.000 316.500 9.600 ;
        RECT 317.400 8.700 319.500 9.600 ;
        RECT 317.700 3.600 319.500 8.700 ;
        RECT 320.700 3.000 322.500 9.600 ;
        RECT 323.700 3.600 325.500 12.600 ;
        RECT 335.700 9.600 337.800 11.700 ;
        RECT 343.200 11.100 346.500 13.200 ;
        RECT 326.700 3.000 328.500 9.600 ;
        RECT 330.300 6.600 332.400 8.700 ;
        RECT 333.300 6.600 335.400 8.700 ;
        RECT 330.300 3.600 332.100 6.600 ;
        RECT 333.300 3.600 335.100 6.600 ;
        RECT 336.300 3.600 338.100 9.600 ;
        RECT 339.300 3.000 341.100 9.600 ;
        RECT 343.200 3.600 345.000 11.100 ;
        RECT 349.200 9.600 351.900 13.500 ;
        RECT 364.200 12.600 369.900 13.800 ;
        RECT 361.500 11.700 363.300 12.300 ;
        RECT 355.200 10.500 363.300 11.700 ;
        RECT 355.200 9.600 357.300 10.500 ;
        RECT 364.200 9.600 365.400 12.600 ;
        RECT 368.100 12.000 369.900 12.600 ;
        RECT 373.800 11.400 374.700 14.700 ;
        RECT 370.800 10.500 374.700 11.400 ;
        RECT 376.500 35.400 378.300 38.400 ;
        RECT 379.500 35.400 381.300 39.000 ;
        RECT 376.500 22.050 378.000 35.400 ;
        RECT 398.100 33.300 399.900 38.400 ;
        RECT 401.100 34.200 402.900 39.000 ;
        RECT 404.100 33.300 405.900 38.400 ;
        RECT 398.100 31.950 405.900 33.300 ;
        RECT 407.100 32.400 408.900 38.400 ;
        RECT 425.100 32.400 426.900 38.400 ;
        RECT 428.100 33.300 429.900 39.000 ;
        RECT 432.600 32.400 434.400 38.400 ;
        RECT 437.100 33.300 438.900 39.000 ;
        RECT 440.100 32.400 441.900 38.400 ;
        RECT 458.100 35.400 459.900 39.000 ;
        RECT 461.100 35.400 462.900 38.400 ;
        RECT 407.100 30.300 408.300 32.400 ;
        RECT 404.700 29.400 408.300 30.300 ;
        RECT 425.700 30.600 426.900 32.400 ;
        RECT 432.900 30.900 434.100 32.400 ;
        RECT 437.100 31.500 441.900 32.400 ;
        RECT 425.700 29.700 432.000 30.600 ;
        RECT 401.100 25.050 402.900 26.850 ;
        RECT 404.700 25.050 405.900 29.400 ;
        RECT 429.900 27.600 432.000 29.700 ;
        RECT 407.100 25.050 408.900 26.850 ;
        RECT 425.400 25.050 427.200 26.850 ;
        RECT 430.200 25.800 432.000 27.600 ;
        RECT 432.900 28.800 435.900 30.900 ;
        RECT 437.100 30.300 439.200 31.500 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 425.100 24.300 427.200 25.050 ;
        RECT 425.100 22.950 432.000 24.300 ;
        RECT 376.500 19.950 378.900 22.050 ;
        RECT 398.100 21.150 399.900 22.950 ;
        RECT 370.800 9.600 372.000 10.500 ;
        RECT 376.500 9.600 378.000 19.950 ;
        RECT 404.700 15.600 405.900 22.950 ;
        RECT 430.200 22.500 432.000 22.950 ;
        RECT 432.900 23.100 434.100 28.800 ;
        RECT 435.000 25.800 437.100 27.900 ;
        RECT 435.300 24.000 437.100 25.800 ;
        RECT 461.100 25.050 462.300 35.400 ;
        RECT 479.400 32.400 481.200 39.000 ;
        RECT 484.500 31.200 486.300 38.400 ;
        RECT 503.400 32.400 505.200 39.000 ;
        RECT 508.500 31.200 510.300 38.400 ;
        RECT 527.100 35.400 528.900 39.000 ;
        RECT 530.100 35.400 531.900 38.400 ;
        RECT 482.100 30.300 486.300 31.200 ;
        RECT 506.100 30.300 510.300 31.200 ;
        RECT 479.250 25.050 481.050 26.850 ;
        RECT 482.100 25.050 483.300 30.300 ;
        RECT 485.100 25.050 486.900 26.850 ;
        RECT 503.250 25.050 505.050 26.850 ;
        RECT 506.100 25.050 507.300 30.300 ;
        RECT 509.100 25.050 510.900 26.850 ;
        RECT 530.100 25.050 531.300 35.400 ;
        RECT 548.100 33.300 549.900 38.400 ;
        RECT 551.100 34.200 552.900 39.000 ;
        RECT 554.100 33.300 555.900 38.400 ;
        RECT 548.100 31.950 555.900 33.300 ;
        RECT 557.100 32.400 558.900 38.400 ;
        RECT 557.100 30.300 558.300 32.400 ;
        RECT 575.700 31.200 577.500 38.400 ;
        RECT 580.800 32.400 582.600 39.000 ;
        RECT 599.100 35.400 600.900 39.000 ;
        RECT 602.100 35.400 603.900 38.400 ;
        RECT 605.100 35.400 606.900 39.000 ;
        RECT 575.700 30.300 579.900 31.200 ;
        RECT 554.700 29.400 558.300 30.300 ;
        RECT 551.100 25.050 552.900 26.850 ;
        RECT 554.700 25.050 555.900 29.400 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 575.100 25.050 576.900 26.850 ;
        RECT 578.700 25.050 579.900 30.300 ;
        RECT 580.950 25.050 582.750 26.850 ;
        RECT 602.700 25.050 603.600 35.400 ;
        RECT 624.000 32.400 625.800 39.000 ;
        RECT 628.500 33.600 630.300 38.400 ;
        RECT 631.500 35.400 633.300 39.000 ;
        RECT 628.500 32.400 633.600 33.600 ;
        RECT 623.100 25.050 624.900 26.850 ;
        RECT 629.250 25.050 631.050 26.850 ;
        RECT 632.700 25.050 633.600 32.400 ;
        RECT 650.100 33.300 651.900 38.400 ;
        RECT 653.100 34.200 654.900 39.000 ;
        RECT 656.100 33.300 657.900 38.400 ;
        RECT 650.100 31.950 657.900 33.300 ;
        RECT 659.100 32.400 660.900 38.400 ;
        RECT 677.400 32.400 679.200 39.000 ;
        RECT 659.100 30.300 660.300 32.400 ;
        RECT 682.500 31.200 684.300 38.400 ;
        RECT 656.700 29.400 660.300 30.300 ;
        RECT 680.100 30.300 684.300 31.200 ;
        RECT 653.100 25.050 654.900 26.850 ;
        RECT 656.700 25.050 657.900 29.400 ;
        RECT 659.100 25.050 660.900 26.850 ;
        RECT 677.250 25.050 679.050 26.850 ;
        RECT 680.100 25.050 681.300 30.300 ;
        RECT 703.500 30.000 705.300 38.400 ;
        RECT 702.000 28.800 705.300 30.000 ;
        RECT 710.100 29.400 711.900 39.000 ;
        RECT 728.700 31.200 730.500 38.400 ;
        RECT 733.800 32.400 735.600 39.000 ;
        RECT 752.100 33.300 753.900 38.400 ;
        RECT 755.100 34.200 756.900 39.000 ;
        RECT 758.100 33.300 759.900 38.400 ;
        RECT 752.100 31.950 759.900 33.300 ;
        RECT 761.100 32.400 762.900 38.400 ;
        RECT 779.100 32.400 780.900 38.400 ;
        RECT 782.100 33.300 783.900 39.000 ;
        RECT 786.300 33.000 788.100 38.400 ;
        RECT 790.800 33.300 792.600 39.000 ;
        RECT 728.700 30.300 732.900 31.200 ;
        RECT 761.100 30.300 762.300 32.400 ;
        RECT 683.100 25.050 684.900 26.850 ;
        RECT 702.000 25.050 702.900 28.800 ;
        RECT 704.100 25.050 705.900 26.850 ;
        RECT 710.100 25.050 711.900 26.850 ;
        RECT 728.100 25.050 729.900 26.850 ;
        RECT 731.700 25.050 732.900 30.300 ;
        RECT 758.700 29.400 762.300 30.300 ;
        RECT 779.100 31.500 780.600 32.400 ;
        RECT 779.100 30.000 783.600 31.500 ;
        RECT 781.500 29.400 783.600 30.000 ;
        RECT 787.200 30.900 788.100 33.000 ;
        RECT 794.100 32.400 795.900 38.400 ;
        RECT 797.700 35.400 799.500 39.000 ;
        RECT 800.700 35.400 802.500 38.400 ;
        RECT 791.400 31.500 795.900 32.400 ;
        RECT 733.950 25.050 735.750 26.850 ;
        RECT 755.100 25.050 756.900 26.850 ;
        RECT 758.700 25.050 759.900 29.400 ;
        RECT 784.500 27.900 786.300 29.700 ;
        RECT 787.200 28.800 790.200 30.900 ;
        RECT 791.400 29.100 793.500 31.500 ;
        RECT 783.900 27.000 786.000 27.900 ;
        RECT 761.100 25.050 762.900 26.850 ;
        RECT 779.400 25.800 786.000 27.000 ;
        RECT 779.400 25.200 781.200 25.800 ;
        RECT 432.900 22.200 435.300 23.100 ;
        RECT 433.800 22.050 435.300 22.200 ;
        RECT 439.800 22.950 441.900 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 779.100 22.950 781.200 25.200 ;
        RECT 429.000 19.500 432.900 21.300 ;
        RECT 430.800 19.200 432.900 19.500 ;
        RECT 433.800 19.950 435.900 22.050 ;
        RECT 439.800 21.150 441.600 22.950 ;
        RECT 458.100 21.150 459.900 22.950 ;
        RECT 433.800 18.000 434.700 19.950 ;
        RECT 427.500 15.600 429.600 17.700 ;
        RECT 433.200 16.950 434.700 18.000 ;
        RECT 433.200 15.600 434.400 16.950 ;
        RECT 346.200 3.000 348.000 9.600 ;
        RECT 349.200 3.600 351.000 9.600 ;
        RECT 352.200 6.600 354.300 8.700 ;
        RECT 355.200 6.600 357.300 8.700 ;
        RECT 358.200 6.600 360.300 8.700 ;
        RECT 352.200 3.600 354.000 6.600 ;
        RECT 355.200 3.600 357.000 6.600 ;
        RECT 358.200 3.600 360.000 6.600 ;
        RECT 361.200 3.000 363.000 9.600 ;
        RECT 364.200 3.600 366.000 9.600 ;
        RECT 367.200 3.000 369.000 9.600 ;
        RECT 370.200 3.600 372.000 9.600 ;
        RECT 373.200 3.000 375.000 9.600 ;
        RECT 376.500 3.600 378.300 9.600 ;
        RECT 379.500 3.000 381.300 9.600 ;
        RECT 398.400 3.000 400.200 15.600 ;
        RECT 403.500 14.100 405.900 15.600 ;
        RECT 425.100 14.700 429.600 15.600 ;
        RECT 403.500 3.600 405.300 14.100 ;
        RECT 406.200 11.100 408.000 12.900 ;
        RECT 406.500 3.000 408.300 9.600 ;
        RECT 425.100 3.600 426.900 14.700 ;
        RECT 428.100 3.000 429.900 13.500 ;
        RECT 432.600 3.600 434.400 15.600 ;
        RECT 437.100 15.600 439.200 16.500 ;
        RECT 437.100 14.400 441.900 15.600 ;
        RECT 437.100 3.000 438.900 13.500 ;
        RECT 440.100 3.600 441.900 14.400 ;
        RECT 461.100 9.600 462.300 22.950 ;
        RECT 482.100 9.600 483.300 22.950 ;
        RECT 506.100 9.600 507.300 22.950 ;
        RECT 527.100 21.150 528.900 22.950 ;
        RECT 530.100 9.600 531.300 22.950 ;
        RECT 548.100 21.150 549.900 22.950 ;
        RECT 554.700 15.600 555.900 22.950 ;
        RECT 458.100 3.000 459.900 9.600 ;
        RECT 461.100 3.600 462.900 9.600 ;
        RECT 479.100 3.000 480.900 9.600 ;
        RECT 482.100 3.600 483.900 9.600 ;
        RECT 485.100 3.000 486.900 9.600 ;
        RECT 503.100 3.000 504.900 9.600 ;
        RECT 506.100 3.600 507.900 9.600 ;
        RECT 509.100 3.000 510.900 9.600 ;
        RECT 527.100 3.000 528.900 9.600 ;
        RECT 530.100 3.600 531.900 9.600 ;
        RECT 548.400 3.000 550.200 15.600 ;
        RECT 553.500 14.100 555.900 15.600 ;
        RECT 553.500 3.600 555.300 14.100 ;
        RECT 556.200 11.100 558.000 12.900 ;
        RECT 578.700 9.600 579.900 22.950 ;
        RECT 599.100 21.150 600.900 22.950 ;
        RECT 602.700 15.600 603.600 22.950 ;
        RECT 604.950 21.150 606.750 22.950 ;
        RECT 626.250 21.150 628.050 22.950 ;
        RECT 632.700 15.600 633.600 22.950 ;
        RECT 650.100 21.150 651.900 22.950 ;
        RECT 656.700 15.600 657.900 22.950 ;
        RECT 600.000 14.400 603.600 15.600 ;
        RECT 556.500 3.000 558.300 9.600 ;
        RECT 575.100 3.000 576.900 9.600 ;
        RECT 578.100 3.600 579.900 9.600 ;
        RECT 581.100 3.000 582.900 9.600 ;
        RECT 600.000 3.600 601.800 14.400 ;
        RECT 605.100 3.000 606.900 15.600 ;
        RECT 623.100 14.700 630.900 15.600 ;
        RECT 623.100 3.600 624.900 14.700 ;
        RECT 626.100 3.000 627.900 13.800 ;
        RECT 629.100 3.600 630.900 14.700 ;
        RECT 632.100 3.600 633.900 15.600 ;
        RECT 650.400 3.000 652.200 15.600 ;
        RECT 655.500 14.100 657.900 15.600 ;
        RECT 655.500 3.600 657.300 14.100 ;
        RECT 658.200 11.100 660.000 12.900 ;
        RECT 680.100 9.600 681.300 22.950 ;
        RECT 702.000 10.800 702.900 22.950 ;
        RECT 707.100 21.150 708.900 22.950 ;
        RECT 703.950 15.450 706.050 16.050 ;
        RECT 727.950 15.450 730.050 16.050 ;
        RECT 703.950 14.550 730.050 15.450 ;
        RECT 703.950 13.950 706.050 14.550 ;
        RECT 727.950 13.950 730.050 14.550 ;
        RECT 702.000 9.900 708.600 10.800 ;
        RECT 702.000 9.600 702.900 9.900 ;
        RECT 658.500 3.000 660.300 9.600 ;
        RECT 677.100 3.000 678.900 9.600 ;
        RECT 680.100 3.600 681.900 9.600 ;
        RECT 683.100 3.000 684.900 9.600 ;
        RECT 701.100 3.600 702.900 9.600 ;
        RECT 707.100 9.600 708.600 9.900 ;
        RECT 731.700 9.600 732.900 22.950 ;
        RECT 752.100 21.150 753.900 22.950 ;
        RECT 758.700 15.600 759.900 22.950 ;
        RECT 783.900 22.800 786.000 24.900 ;
        RECT 783.900 21.000 785.700 22.800 ;
        RECT 787.200 22.050 788.100 28.800 ;
        RECT 789.000 24.900 791.100 27.000 ;
        RECT 789.000 23.100 790.800 24.900 ;
        RECT 793.800 22.950 795.900 25.050 ;
        RECT 787.200 20.700 790.200 22.050 ;
        RECT 793.800 21.150 795.600 22.950 ;
        RECT 801.000 22.050 802.500 35.400 ;
        RECT 788.100 19.950 790.200 20.700 ;
        RECT 800.100 19.950 802.500 22.050 ;
        RECT 785.400 17.700 787.200 19.500 ;
        RECT 781.800 16.800 787.200 17.700 ;
        RECT 781.800 15.900 783.900 16.800 ;
        RECT 704.100 3.000 705.900 9.000 ;
        RECT 707.100 3.600 708.900 9.600 ;
        RECT 710.100 3.000 711.900 9.600 ;
        RECT 728.100 3.000 729.900 9.600 ;
        RECT 731.100 3.600 732.900 9.600 ;
        RECT 734.100 3.000 735.900 9.600 ;
        RECT 752.400 3.000 754.200 15.600 ;
        RECT 757.500 14.100 759.900 15.600 ;
        RECT 779.100 14.700 783.900 15.900 ;
        RECT 788.700 15.600 789.900 19.950 ;
        RECT 786.600 14.700 789.900 15.600 ;
        RECT 790.800 15.600 792.900 16.500 ;
        RECT 757.500 3.600 759.300 14.100 ;
        RECT 760.200 11.100 762.000 12.900 ;
        RECT 760.500 3.000 762.300 9.600 ;
        RECT 779.100 3.600 780.900 14.700 ;
        RECT 782.100 3.000 783.900 13.500 ;
        RECT 786.600 3.600 788.400 14.700 ;
        RECT 790.800 14.400 795.900 15.600 ;
        RECT 790.800 3.000 792.900 13.500 ;
        RECT 794.100 3.600 795.900 14.400 ;
        RECT 801.000 9.600 802.500 19.950 ;
        RECT 804.300 32.400 806.100 38.400 ;
        RECT 809.700 32.400 811.500 39.000 ;
        RECT 814.800 33.600 816.600 38.400 ;
        RECT 819.000 35.400 820.800 38.400 ;
        RECT 822.000 35.400 823.800 38.400 ;
        RECT 825.000 35.400 826.800 38.400 ;
        RECT 828.000 35.400 829.800 38.400 ;
        RECT 831.000 35.400 832.800 39.000 ;
        RECT 812.400 32.400 816.600 33.600 ;
        RECT 818.700 33.300 820.800 35.400 ;
        RECT 821.700 33.300 823.800 35.400 ;
        RECT 824.700 33.300 826.800 35.400 ;
        RECT 827.700 33.300 829.800 35.400 ;
        RECT 834.000 34.500 835.800 38.400 ;
        RECT 838.500 35.400 840.300 39.000 ;
        RECT 841.500 35.400 843.300 38.400 ;
        RECT 844.500 35.400 846.300 38.400 ;
        RECT 847.500 35.400 849.300 38.400 ;
        RECT 833.100 32.400 835.800 34.500 ;
        RECT 837.600 33.600 839.400 34.500 ;
        RECT 837.600 32.400 840.300 33.600 ;
        RECT 841.200 33.300 843.300 35.400 ;
        RECT 844.200 33.300 846.300 35.400 ;
        RECT 847.200 33.300 849.300 35.400 ;
        RECT 851.700 32.400 853.500 38.400 ;
        RECT 857.100 32.400 858.900 39.000 ;
        RECT 862.500 32.400 864.300 38.400 ;
        RECT 804.300 15.600 805.200 32.400 ;
        RECT 812.400 29.100 813.900 32.400 ;
        RECT 818.100 30.600 824.700 32.400 ;
        RECT 839.400 31.800 840.300 32.400 ;
        RECT 842.400 31.800 844.200 32.400 ;
        RECT 839.400 30.600 846.600 31.800 ;
        RECT 806.100 27.300 813.900 29.100 ;
        RECT 830.100 28.500 831.900 30.300 ;
        RECT 829.800 27.900 831.900 28.500 ;
        RECT 814.800 26.400 831.900 27.900 ;
        RECT 836.100 27.900 838.200 28.050 ;
        RECT 839.400 27.900 841.200 28.800 ;
        RECT 836.100 27.000 841.200 27.900 ;
        RECT 845.700 27.600 846.600 30.600 ;
        RECT 851.700 31.500 853.200 32.400 ;
        RECT 851.700 30.300 860.100 31.500 ;
        RECT 858.300 29.700 860.100 30.300 ;
        RECT 847.500 28.800 849.600 29.700 ;
        RECT 863.100 28.800 864.300 32.400 ;
        RECT 881.100 35.400 882.900 38.400 ;
        RECT 881.100 31.500 882.300 35.400 ;
        RECT 884.100 32.400 885.900 39.000 ;
        RECT 887.100 32.400 888.900 38.400 ;
        RECT 881.100 30.600 886.800 31.500 ;
        RECT 847.500 27.600 864.300 28.800 ;
        RECT 809.700 24.900 816.300 26.400 ;
        RECT 836.100 25.950 838.200 27.000 ;
        RECT 844.800 25.800 846.600 27.600 ;
        RECT 809.700 22.050 811.200 24.900 ;
        RECT 817.500 23.700 861.900 24.900 ;
        RECT 817.500 22.200 818.400 23.700 ;
        RECT 809.100 19.950 811.200 22.050 ;
        RECT 813.300 20.400 818.400 22.200 ;
        RECT 821.100 21.900 834.600 22.800 ;
        RECT 841.800 21.900 843.600 22.500 ;
        RECT 860.100 22.050 861.900 23.700 ;
        RECT 821.100 20.700 822.000 21.900 ;
        RECT 821.100 18.900 822.900 20.700 ;
        RECT 827.100 19.200 831.000 21.000 ;
        RECT 832.500 20.700 843.600 21.900 ;
        RECT 854.100 21.750 856.200 22.050 ;
        RECT 832.500 19.800 834.600 20.700 ;
        RECT 852.300 19.950 856.200 21.750 ;
        RECT 860.100 19.950 862.200 22.050 ;
        RECT 852.300 19.200 854.100 19.950 ;
        RECT 827.100 18.900 829.200 19.200 ;
        RECT 840.600 18.300 854.100 19.200 ;
        RECT 806.100 17.700 807.900 18.300 ;
        RECT 840.600 17.700 841.800 18.300 ;
        RECT 806.100 16.500 841.800 17.700 ;
        RECT 844.500 16.500 846.600 16.800 ;
        RECT 804.300 14.700 820.800 15.600 ;
        RECT 804.300 11.400 805.200 14.700 ;
        RECT 809.100 12.600 814.800 13.800 ;
        RECT 818.700 13.500 820.800 14.700 ;
        RECT 824.100 14.400 841.800 15.600 ;
        RECT 844.500 15.300 856.500 16.500 ;
        RECT 844.500 14.700 846.600 15.300 ;
        RECT 854.700 14.700 856.500 15.300 ;
        RECT 824.100 13.500 826.200 14.400 ;
        RECT 840.600 13.800 841.800 14.400 ;
        RECT 858.000 13.800 859.800 14.100 ;
        RECT 809.100 12.000 810.900 12.600 ;
        RECT 804.300 10.500 808.200 11.400 ;
        RECT 807.000 9.600 808.200 10.500 ;
        RECT 813.600 9.600 814.800 12.600 ;
        RECT 815.700 11.700 817.500 12.300 ;
        RECT 815.700 10.500 823.800 11.700 ;
        RECT 821.700 9.600 823.800 10.500 ;
        RECT 827.100 9.600 829.800 13.500 ;
        RECT 832.500 11.100 835.800 13.200 ;
        RECT 840.600 12.600 859.800 13.800 ;
        RECT 797.700 3.000 799.500 9.600 ;
        RECT 800.700 3.600 802.500 9.600 ;
        RECT 804.000 3.000 805.800 9.600 ;
        RECT 807.000 3.600 808.800 9.600 ;
        RECT 810.000 3.000 811.800 9.600 ;
        RECT 813.000 3.600 814.800 9.600 ;
        RECT 816.000 3.000 817.800 9.600 ;
        RECT 818.700 6.600 820.800 8.700 ;
        RECT 821.700 6.600 823.800 8.700 ;
        RECT 824.700 6.600 826.800 8.700 ;
        RECT 819.000 3.600 820.800 6.600 ;
        RECT 822.000 3.600 823.800 6.600 ;
        RECT 825.000 3.600 826.800 6.600 ;
        RECT 828.000 3.600 829.800 9.600 ;
        RECT 831.000 3.000 832.800 9.600 ;
        RECT 834.000 3.600 835.800 11.100 ;
        RECT 841.200 9.600 843.300 11.700 ;
        RECT 837.900 3.000 839.700 9.600 ;
        RECT 840.900 3.600 842.700 9.600 ;
        RECT 843.600 6.600 845.700 8.700 ;
        RECT 846.600 6.600 848.700 8.700 ;
        RECT 843.900 3.600 845.700 6.600 ;
        RECT 846.900 3.600 848.700 6.600 ;
        RECT 850.500 3.000 852.300 9.600 ;
        RECT 853.500 3.600 855.300 12.600 ;
        RECT 858.000 12.300 859.800 12.600 ;
        RECT 863.100 11.400 864.300 27.600 ;
        RECT 885.000 29.700 886.800 30.600 ;
        RECT 881.400 22.950 883.500 25.050 ;
        RECT 881.400 21.150 883.200 22.950 ;
        RECT 885.000 18.300 885.900 29.700 ;
        RECT 887.700 25.050 888.900 32.400 ;
        RECT 886.800 22.950 888.900 25.050 ;
        RECT 885.000 17.400 886.800 18.300 ;
        RECT 860.700 10.500 864.300 11.400 ;
        RECT 881.100 16.500 886.800 17.400 ;
        RECT 860.700 9.600 861.600 10.500 ;
        RECT 881.100 9.600 882.300 16.500 ;
        RECT 887.700 15.600 888.900 22.950 ;
        RECT 856.500 3.000 858.300 9.600 ;
        RECT 859.500 8.700 861.600 9.600 ;
        RECT 859.500 3.600 861.300 8.700 ;
        RECT 862.500 3.000 864.300 9.600 ;
        RECT 881.100 3.600 882.900 9.600 ;
        RECT 884.100 3.000 885.900 13.800 ;
        RECT 887.100 3.600 888.900 15.600 ;
        RECT 890.700 32.400 892.500 38.400 ;
        RECT 896.100 32.400 897.900 39.000 ;
        RECT 901.500 32.400 903.300 38.400 ;
        RECT 905.700 35.400 907.500 38.400 ;
        RECT 908.700 35.400 910.500 38.400 ;
        RECT 911.700 35.400 913.500 38.400 ;
        RECT 914.700 35.400 916.500 39.000 ;
        RECT 905.700 33.300 907.800 35.400 ;
        RECT 908.700 33.300 910.800 35.400 ;
        RECT 911.700 33.300 913.800 35.400 ;
        RECT 919.200 34.500 921.000 38.400 ;
        RECT 922.200 35.400 924.000 39.000 ;
        RECT 925.200 35.400 927.000 38.400 ;
        RECT 928.200 35.400 930.000 38.400 ;
        RECT 931.200 35.400 933.000 38.400 ;
        RECT 934.200 35.400 936.000 38.400 ;
        RECT 915.600 33.600 917.400 34.500 ;
        RECT 914.700 32.400 917.400 33.600 ;
        RECT 919.200 32.400 921.900 34.500 ;
        RECT 925.200 33.300 927.300 35.400 ;
        RECT 928.200 33.300 930.300 35.400 ;
        RECT 931.200 33.300 933.300 35.400 ;
        RECT 934.200 33.300 936.300 35.400 ;
        RECT 938.400 33.600 940.200 38.400 ;
        RECT 938.400 32.400 942.600 33.600 ;
        RECT 943.500 32.400 945.300 39.000 ;
        RECT 948.900 32.400 950.700 38.400 ;
        RECT 890.700 28.800 891.900 32.400 ;
        RECT 901.800 31.500 903.300 32.400 ;
        RECT 910.800 31.800 912.600 32.400 ;
        RECT 914.700 31.800 915.600 32.400 ;
        RECT 894.900 30.300 903.300 31.500 ;
        RECT 908.400 30.600 915.600 31.800 ;
        RECT 930.300 30.600 936.900 32.400 ;
        RECT 894.900 29.700 896.700 30.300 ;
        RECT 905.400 28.800 907.500 29.700 ;
        RECT 890.700 27.600 907.500 28.800 ;
        RECT 908.400 27.600 909.300 30.600 ;
        RECT 913.800 27.900 915.600 28.800 ;
        RECT 923.100 28.500 924.900 30.300 ;
        RECT 941.100 29.100 942.600 32.400 ;
        RECT 916.800 27.900 918.900 28.050 ;
        RECT 890.700 11.400 891.900 27.600 ;
        RECT 908.400 25.800 910.200 27.600 ;
        RECT 913.800 27.000 918.900 27.900 ;
        RECT 916.800 25.950 918.900 27.000 ;
        RECT 923.100 27.900 925.200 28.500 ;
        RECT 923.100 26.400 940.200 27.900 ;
        RECT 941.100 27.300 948.900 29.100 ;
        RECT 938.700 24.900 945.300 26.400 ;
        RECT 893.100 23.700 937.500 24.900 ;
        RECT 893.100 22.050 894.900 23.700 ;
        RECT 892.800 19.950 894.900 22.050 ;
        RECT 898.800 21.750 900.900 22.050 ;
        RECT 911.400 21.900 913.200 22.500 ;
        RECT 920.400 21.900 933.900 22.800 ;
        RECT 898.800 19.950 902.700 21.750 ;
        RECT 911.400 20.700 922.500 21.900 ;
        RECT 900.900 19.200 902.700 19.950 ;
        RECT 920.400 19.800 922.500 20.700 ;
        RECT 924.000 19.200 927.900 21.000 ;
        RECT 933.000 20.700 933.900 21.900 ;
        RECT 900.900 18.300 914.400 19.200 ;
        RECT 925.800 18.900 927.900 19.200 ;
        RECT 932.100 18.900 933.900 20.700 ;
        RECT 936.600 22.200 937.500 23.700 ;
        RECT 936.600 20.400 941.700 22.200 ;
        RECT 943.800 22.050 945.300 24.900 ;
        RECT 943.800 19.950 945.900 22.050 ;
        RECT 913.200 17.700 914.400 18.300 ;
        RECT 947.100 17.700 948.900 18.300 ;
        RECT 908.400 16.500 910.500 16.800 ;
        RECT 913.200 16.500 948.900 17.700 ;
        RECT 898.500 15.300 910.500 16.500 ;
        RECT 949.800 15.600 950.700 32.400 ;
        RECT 898.500 14.700 900.300 15.300 ;
        RECT 908.400 14.700 910.500 15.300 ;
        RECT 913.200 14.400 930.900 15.600 ;
        RECT 895.200 13.800 897.000 14.100 ;
        RECT 913.200 13.800 914.400 14.400 ;
        RECT 895.200 12.600 914.400 13.800 ;
        RECT 928.800 13.500 930.900 14.400 ;
        RECT 934.200 14.700 950.700 15.600 ;
        RECT 934.200 13.500 936.300 14.700 ;
        RECT 895.200 12.300 897.000 12.600 ;
        RECT 890.700 10.500 894.300 11.400 ;
        RECT 893.400 9.600 894.300 10.500 ;
        RECT 890.700 3.000 892.500 9.600 ;
        RECT 893.400 8.700 895.500 9.600 ;
        RECT 893.700 3.600 895.500 8.700 ;
        RECT 896.700 3.000 898.500 9.600 ;
        RECT 899.700 3.600 901.500 12.600 ;
        RECT 911.700 9.600 913.800 11.700 ;
        RECT 919.200 11.100 922.500 13.200 ;
        RECT 902.700 3.000 904.500 9.600 ;
        RECT 906.300 6.600 908.400 8.700 ;
        RECT 909.300 6.600 911.400 8.700 ;
        RECT 906.300 3.600 908.100 6.600 ;
        RECT 909.300 3.600 911.100 6.600 ;
        RECT 912.300 3.600 914.100 9.600 ;
        RECT 915.300 3.000 917.100 9.600 ;
        RECT 919.200 3.600 921.000 11.100 ;
        RECT 925.200 9.600 927.900 13.500 ;
        RECT 940.200 12.600 945.900 13.800 ;
        RECT 937.500 11.700 939.300 12.300 ;
        RECT 931.200 10.500 939.300 11.700 ;
        RECT 931.200 9.600 933.300 10.500 ;
        RECT 940.200 9.600 941.400 12.600 ;
        RECT 944.100 12.000 945.900 12.600 ;
        RECT 949.800 11.400 950.700 14.700 ;
        RECT 946.800 10.500 950.700 11.400 ;
        RECT 952.500 35.400 954.300 38.400 ;
        RECT 955.500 35.400 957.300 39.000 ;
        RECT 952.500 22.050 954.000 35.400 ;
        RECT 974.100 32.400 975.900 38.400 ;
        RECT 974.700 30.300 975.900 32.400 ;
        RECT 977.100 33.300 978.900 38.400 ;
        RECT 980.100 34.200 981.900 39.000 ;
        RECT 983.100 33.300 984.900 38.400 ;
        RECT 977.100 31.950 984.900 33.300 ;
        RECT 1001.100 32.400 1002.900 38.400 ;
        RECT 1004.100 33.300 1005.900 39.000 ;
        RECT 1008.600 32.400 1010.400 38.400 ;
        RECT 1013.100 33.300 1014.900 39.000 ;
        RECT 1016.100 32.400 1017.900 38.400 ;
        RECT 1001.100 31.500 1005.900 32.400 ;
        RECT 1003.800 30.300 1005.900 31.500 ;
        RECT 1008.900 30.900 1010.100 32.400 ;
        RECT 974.700 29.400 978.300 30.300 ;
        RECT 974.100 25.050 975.900 26.850 ;
        RECT 977.100 25.050 978.300 29.400 ;
        RECT 1007.100 28.800 1010.100 30.900 ;
        RECT 1016.100 30.600 1017.300 32.400 ;
        RECT 980.100 25.050 981.900 26.850 ;
        RECT 1005.900 25.800 1008.000 27.900 ;
        RECT 973.950 22.950 976.050 25.050 ;
        RECT 976.950 22.950 979.050 25.050 ;
        RECT 979.950 22.950 982.050 25.050 ;
        RECT 982.950 22.950 985.050 25.050 ;
        RECT 1001.100 22.950 1003.200 25.050 ;
        RECT 1005.900 24.000 1007.700 25.800 ;
        RECT 1008.900 23.100 1010.100 28.800 ;
        RECT 1011.000 29.700 1017.300 30.600 ;
        RECT 1034.700 31.200 1036.500 38.400 ;
        RECT 1039.800 32.400 1041.600 39.000 ;
        RECT 1034.700 30.300 1038.900 31.200 ;
        RECT 1011.000 27.600 1013.100 29.700 ;
        RECT 1011.000 25.800 1012.800 27.600 ;
        RECT 1015.800 25.050 1017.600 26.850 ;
        RECT 1034.100 25.050 1035.900 26.850 ;
        RECT 1037.700 25.050 1038.900 30.300 ;
        RECT 1039.950 25.050 1041.750 26.850 ;
        RECT 1015.800 24.300 1017.900 25.050 ;
        RECT 952.500 19.950 954.900 22.050 ;
        RECT 946.800 9.600 948.000 10.500 ;
        RECT 952.500 9.600 954.000 19.950 ;
        RECT 977.100 15.600 978.300 22.950 ;
        RECT 983.100 21.150 984.900 22.950 ;
        RECT 1001.400 21.150 1003.200 22.950 ;
        RECT 1007.700 22.200 1010.100 23.100 ;
        RECT 1011.000 22.950 1017.900 24.300 ;
        RECT 1033.950 22.950 1036.050 25.050 ;
        RECT 1036.950 22.950 1039.050 25.050 ;
        RECT 1039.950 22.950 1042.050 25.050 ;
        RECT 1011.000 22.500 1012.800 22.950 ;
        RECT 1007.700 22.050 1009.200 22.200 ;
        RECT 1007.100 19.950 1009.200 22.050 ;
        RECT 1008.300 18.000 1009.200 19.950 ;
        RECT 1010.100 19.500 1014.000 21.300 ;
        RECT 1010.100 19.200 1012.200 19.500 ;
        RECT 1024.950 18.450 1027.050 19.050 ;
        RECT 1033.950 18.450 1036.050 19.050 ;
        RECT 1008.300 16.950 1009.800 18.000 ;
        RECT 1003.800 15.600 1005.900 16.500 ;
        RECT 977.100 14.100 979.500 15.600 ;
        RECT 975.000 11.100 976.800 12.900 ;
        RECT 922.200 3.000 924.000 9.600 ;
        RECT 925.200 3.600 927.000 9.600 ;
        RECT 928.200 6.600 930.300 8.700 ;
        RECT 931.200 6.600 933.300 8.700 ;
        RECT 934.200 6.600 936.300 8.700 ;
        RECT 928.200 3.600 930.000 6.600 ;
        RECT 931.200 3.600 933.000 6.600 ;
        RECT 934.200 3.600 936.000 6.600 ;
        RECT 937.200 3.000 939.000 9.600 ;
        RECT 940.200 3.600 942.000 9.600 ;
        RECT 943.200 3.000 945.000 9.600 ;
        RECT 946.200 3.600 948.000 9.600 ;
        RECT 949.200 3.000 951.000 9.600 ;
        RECT 952.500 3.600 954.300 9.600 ;
        RECT 955.500 3.000 957.300 9.600 ;
        RECT 974.700 3.000 976.500 9.600 ;
        RECT 977.700 3.600 979.500 14.100 ;
        RECT 982.800 3.000 984.600 15.600 ;
        RECT 1001.100 14.400 1005.900 15.600 ;
        RECT 1008.600 15.600 1009.800 16.950 ;
        RECT 1013.400 15.600 1015.500 17.700 ;
        RECT 1024.950 17.550 1036.050 18.450 ;
        RECT 1024.950 16.950 1027.050 17.550 ;
        RECT 1033.950 16.950 1036.050 17.550 ;
        RECT 1001.100 3.600 1002.900 14.400 ;
        RECT 1004.100 3.000 1005.900 13.500 ;
        RECT 1008.600 3.600 1010.400 15.600 ;
        RECT 1013.400 14.700 1017.900 15.600 ;
        RECT 1013.100 3.000 1014.900 13.500 ;
        RECT 1016.100 3.600 1017.900 14.700 ;
        RECT 1037.700 9.600 1038.900 22.950 ;
        RECT 1034.100 3.000 1035.900 9.600 ;
        RECT 1037.100 3.600 1038.900 9.600 ;
        RECT 1040.100 3.000 1041.900 9.600 ;
      LAYER metal2 ;
        RECT 89.700 969.300 91.800 971.400 ;
        RECT 92.700 969.300 94.800 971.400 ;
        RECT 95.700 969.300 97.800 971.400 ;
        RECT 90.300 965.700 91.500 969.300 ;
        RECT 22.950 962.100 25.050 964.200 ;
        RECT 40.950 962.100 43.050 964.200 ;
        RECT 61.950 963.450 64.050 964.200 ;
        RECT 89.400 963.600 91.500 965.700 ;
        RECT 65.400 963.450 66.600 963.600 ;
        RECT 61.950 962.400 66.600 963.450 ;
        RECT 61.950 962.100 64.050 962.400 ;
        RECT 23.400 961.350 24.600 962.100 ;
        RECT 41.400 961.350 42.600 962.100 ;
        RECT 17.100 958.950 19.200 961.050 ;
        RECT 22.500 958.950 24.600 961.050 ;
        RECT 41.400 958.950 43.500 961.050 ;
        RECT 46.800 958.950 48.900 961.050 ;
        RECT 52.950 946.950 55.050 949.050 ;
        RECT 25.950 917.100 28.050 919.200 ;
        RECT 37.950 917.100 40.050 919.200 ;
        RECT 53.400 918.600 54.450 946.950 ;
        RECT 26.400 916.350 27.600 917.100 ;
        RECT 20.100 913.950 22.200 916.050 ;
        RECT 26.100 913.950 28.200 916.050 ;
        RECT 38.400 912.900 39.450 917.100 ;
        RECT 53.400 916.350 54.600 918.600 ;
        RECT 47.400 913.950 49.500 916.050 ;
        RECT 52.800 913.950 54.900 916.050 ;
        RECT 47.400 912.900 48.600 913.650 ;
        RECT 37.950 910.800 40.050 912.900 ;
        RECT 46.950 910.800 49.050 912.900 ;
        RECT 38.400 886.200 39.450 910.800 ;
        RECT 62.400 910.050 63.450 962.100 ;
        RECT 65.400 961.350 66.600 962.400 ;
        RECT 65.400 958.950 67.500 961.050 ;
        RECT 70.800 958.950 72.900 961.050 ;
        RECT 83.400 960.450 84.600 960.600 ;
        RECT 83.400 959.400 87.450 960.450 ;
        RECT 83.400 958.350 84.600 959.400 ;
        RECT 76.800 955.950 78.900 958.050 ;
        RECT 82.800 955.950 84.900 958.050 ;
        RECT 86.400 949.050 87.450 959.400 ;
        RECT 85.950 946.950 88.050 949.050 ;
        RECT 86.400 943.050 87.450 946.950 ;
        RECT 89.400 944.700 90.900 963.600 ;
        RECT 93.300 952.800 94.500 969.300 ;
        RECT 92.400 950.700 94.500 952.800 ;
        RECT 93.300 944.700 94.500 950.700 ;
        RECT 95.700 947.700 96.900 969.300 ;
        RECT 103.800 968.400 105.900 970.500 ;
        RECT 109.200 969.300 111.300 971.400 ;
        RECT 112.200 969.300 114.300 971.400 ;
        RECT 115.200 969.300 117.300 971.400 ;
        RECT 100.800 961.950 102.900 964.050 ;
        RECT 101.400 959.400 102.600 961.650 ;
        RECT 95.700 945.600 97.800 947.700 ;
        RECT 85.950 940.950 88.050 943.050 ;
        RECT 89.400 942.600 92.400 944.700 ;
        RECT 93.300 942.600 95.400 944.700 ;
        RECT 101.400 937.050 102.450 959.400 ;
        RECT 104.400 957.900 105.300 968.400 ;
        RECT 107.100 962.400 109.200 964.500 ;
        RECT 104.400 955.800 106.500 957.900 ;
        RECT 110.100 957.000 111.300 969.300 ;
        RECT 104.400 949.200 105.300 955.800 ;
        RECT 109.800 954.900 111.900 957.000 ;
        RECT 104.400 947.100 106.500 949.200 ;
        RECT 110.100 947.700 111.300 954.900 ;
        RECT 112.800 951.600 114.300 969.300 ;
        RECT 112.800 949.500 114.900 951.600 ;
        RECT 109.800 945.600 111.900 947.700 ;
        RECT 112.800 944.700 114.300 949.500 ;
        RECT 116.100 947.700 117.300 969.300 ;
        RECT 112.200 942.600 114.300 944.700 ;
        RECT 115.200 942.600 117.300 947.700 ;
        RECT 118.200 969.300 120.300 971.400 ;
        RECT 158.700 969.300 160.800 971.400 ;
        RECT 161.700 969.300 163.800 971.400 ;
        RECT 164.700 969.300 166.800 971.400 ;
        RECT 118.200 951.600 119.700 969.300 ;
        RECT 159.300 965.700 160.500 969.300 ;
        RECT 121.950 961.950 124.050 964.050 ;
        RECT 118.200 949.500 120.300 951.600 ;
        RECT 118.200 944.700 119.700 949.500 ;
        RECT 118.200 942.600 120.300 944.700 ;
        RECT 100.950 934.950 103.050 937.050 ;
        RECT 106.950 934.950 109.050 937.050 ;
        RECT 79.950 917.100 82.050 919.200 ;
        RECT 97.950 917.100 100.050 919.200 ;
        RECT 71.100 913.950 73.200 916.050 ;
        RECT 76.500 913.950 78.600 916.050 ;
        RECT 77.400 912.450 78.600 913.650 ;
        RECT 80.400 912.450 81.450 917.100 ;
        RECT 98.400 916.350 99.600 917.100 ;
        RECT 94.950 913.950 97.050 916.050 ;
        RECT 97.950 913.950 100.050 916.050 ;
        RECT 100.950 913.950 103.050 916.050 ;
        RECT 77.400 911.400 81.450 912.450 ;
        RECT 95.400 911.400 96.600 913.650 ;
        RECT 101.400 911.400 102.600 913.650 ;
        RECT 107.400 913.050 108.450 934.950 ;
        RECT 122.400 934.050 123.450 961.950 ;
        RECT 128.400 960.450 129.600 960.600 ;
        RECT 128.400 959.400 132.450 960.450 ;
        RECT 136.950 960.000 139.050 964.050 ;
        RECT 158.400 963.600 160.500 965.700 ;
        RECT 128.400 958.350 129.600 959.400 ;
        RECT 127.800 955.950 129.900 958.050 ;
        RECT 131.400 952.050 132.450 959.400 ;
        RECT 137.400 958.350 138.600 960.000 ;
        RECT 136.800 955.950 138.900 958.050 ;
        RECT 145.800 955.950 147.900 958.050 ;
        RECT 151.800 955.950 153.900 958.050 ;
        RECT 146.400 953.400 147.600 955.650 ;
        RECT 130.950 949.950 133.050 952.050 ;
        RECT 136.950 949.950 139.050 952.050 ;
        RECT 121.950 931.950 124.050 934.050 ;
        RECT 118.950 917.100 121.050 919.200 ;
        RECT 124.950 918.000 127.050 922.050 ;
        RECT 133.950 919.950 136.050 922.050 ;
        RECT 119.400 916.350 120.600 917.100 ;
        RECT 125.400 916.350 126.600 918.000 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 121.950 913.950 124.050 916.050 ;
        RECT 124.950 913.950 127.050 916.050 ;
        RECT 127.950 913.950 130.050 916.050 ;
        RECT 61.950 907.950 64.050 910.050 ;
        RECT 73.950 907.950 76.050 910.050 ;
        RECT 41.700 891.300 43.800 893.400 ;
        RECT 44.700 891.300 46.800 893.400 ;
        RECT 47.700 891.300 49.800 893.400 ;
        RECT 42.300 887.700 43.500 891.300 ;
        RECT 22.950 884.100 25.050 886.200 ;
        RECT 37.950 884.100 40.050 886.200 ;
        RECT 41.400 885.600 43.500 887.700 ;
        RECT 23.400 883.350 24.600 884.100 ;
        RECT 17.100 880.950 19.200 883.050 ;
        RECT 22.500 880.950 24.600 883.050 ;
        RECT 17.400 879.000 18.600 880.650 ;
        RECT 16.950 874.800 19.050 879.000 ;
        RECT 28.800 877.950 30.900 880.050 ;
        RECT 34.800 877.950 36.900 880.050 ;
        RECT 29.400 876.900 30.600 877.650 ;
        RECT 28.950 874.800 31.050 876.900 ;
        RECT 29.400 859.050 30.450 874.800 ;
        RECT 7.950 856.950 10.050 859.050 ;
        RECT 28.950 856.950 31.050 859.050 ;
        RECT 8.400 805.050 9.450 856.950 ;
        RECT 29.400 843.600 30.450 856.950 ;
        RECT 29.400 841.350 30.600 843.600 ;
        RECT 28.800 838.950 30.900 841.050 ;
        RECT 34.800 838.950 36.900 841.050 ;
        RECT 17.100 835.950 19.200 838.050 ;
        RECT 22.500 835.950 24.600 838.050 ;
        RECT 23.400 833.400 24.600 835.650 ;
        RECT 23.400 826.050 24.450 833.400 ;
        RECT 22.950 823.950 25.050 826.050 ;
        RECT 38.400 823.050 39.450 884.100 ;
        RECT 41.400 866.700 42.900 885.600 ;
        RECT 45.300 874.800 46.500 891.300 ;
        RECT 44.400 872.700 46.500 874.800 ;
        RECT 45.300 866.700 46.500 872.700 ;
        RECT 47.700 869.700 48.900 891.300 ;
        RECT 55.800 890.400 57.900 892.500 ;
        RECT 61.200 891.300 63.300 893.400 ;
        RECT 64.200 891.300 66.300 893.400 ;
        RECT 67.200 891.300 69.300 893.400 ;
        RECT 52.800 883.950 54.900 886.050 ;
        RECT 53.400 881.400 54.600 883.650 ;
        RECT 47.700 867.600 49.800 869.700 ;
        RECT 53.400 868.050 54.450 881.400 ;
        RECT 56.400 879.900 57.300 890.400 ;
        RECT 59.100 884.400 61.200 886.500 ;
        RECT 56.400 877.800 58.500 879.900 ;
        RECT 62.100 879.000 63.300 891.300 ;
        RECT 56.400 871.200 57.300 877.800 ;
        RECT 61.800 876.900 63.900 879.000 ;
        RECT 56.400 869.100 58.500 871.200 ;
        RECT 62.100 869.700 63.300 876.900 ;
        RECT 64.800 873.600 66.300 891.300 ;
        RECT 64.800 871.500 66.900 873.600 ;
        RECT 41.400 864.600 44.400 866.700 ;
        RECT 45.300 864.600 47.400 866.700 ;
        RECT 52.950 865.950 55.050 868.050 ;
        RECT 61.800 867.600 63.900 869.700 ;
        RECT 64.800 866.700 66.300 871.500 ;
        RECT 68.100 869.700 69.300 891.300 ;
        RECT 64.200 864.600 66.300 866.700 ;
        RECT 67.200 864.600 69.300 869.700 ;
        RECT 70.200 891.300 72.300 893.400 ;
        RECT 70.200 873.600 71.700 891.300 ;
        RECT 70.200 871.500 72.300 873.600 ;
        RECT 70.200 866.700 71.700 871.500 ;
        RECT 70.200 864.600 72.300 866.700 ;
        RECT 41.400 852.300 44.400 854.400 ;
        RECT 45.300 852.300 47.400 854.400 ;
        RECT 64.200 852.300 66.300 854.400 ;
        RECT 41.400 833.400 42.900 852.300 ;
        RECT 45.300 846.300 46.500 852.300 ;
        RECT 44.400 844.200 46.500 846.300 ;
        RECT 41.400 831.300 43.500 833.400 ;
        RECT 42.300 827.700 43.500 831.300 ;
        RECT 45.300 827.700 46.500 844.200 ;
        RECT 47.700 849.300 49.800 851.400 ;
        RECT 47.700 827.700 48.900 849.300 ;
        RECT 56.400 847.800 58.500 849.900 ;
        RECT 61.800 849.300 63.900 851.400 ;
        RECT 52.950 841.950 55.050 844.050 ;
        RECT 53.400 837.600 54.450 841.950 ;
        RECT 56.400 841.200 57.300 847.800 ;
        RECT 62.100 842.100 63.300 849.300 ;
        RECT 64.800 847.500 66.300 852.300 ;
        RECT 67.200 849.300 69.300 854.400 ;
        RECT 64.800 845.400 66.900 847.500 ;
        RECT 56.400 839.100 58.500 841.200 ;
        RECT 61.800 840.000 63.900 842.100 ;
        RECT 53.400 835.350 54.600 837.600 ;
        RECT 52.800 832.950 54.900 835.050 ;
        RECT 56.400 828.600 57.300 839.100 ;
        RECT 59.100 832.500 61.200 834.600 ;
        RECT 41.700 825.600 43.800 827.700 ;
        RECT 44.700 825.600 46.800 827.700 ;
        RECT 47.700 825.600 49.800 827.700 ;
        RECT 55.800 826.500 57.900 828.600 ;
        RECT 62.100 827.700 63.300 840.000 ;
        RECT 64.800 827.700 66.300 845.400 ;
        RECT 68.100 827.700 69.300 849.300 ;
        RECT 61.200 825.600 63.300 827.700 ;
        RECT 64.200 825.600 66.300 827.700 ;
        RECT 67.200 825.600 69.300 827.700 ;
        RECT 70.200 852.300 72.300 854.400 ;
        RECT 70.200 847.500 71.700 852.300 ;
        RECT 70.200 845.400 72.300 847.500 ;
        RECT 70.200 827.700 71.700 845.400 ;
        RECT 70.200 825.600 72.300 827.700 ;
        RECT 74.400 825.450 75.450 907.950 ;
        RECT 79.950 895.950 82.050 898.050 ;
        RECT 80.400 882.600 81.450 895.950 ;
        RECT 80.400 882.450 81.600 882.600 ;
        RECT 80.400 881.400 84.450 882.450 ;
        RECT 80.400 880.350 81.600 881.400 ;
        RECT 79.800 877.950 81.900 880.050 ;
        RECT 79.800 838.950 81.900 841.050 ;
        RECT 80.400 837.450 81.600 838.650 ;
        RECT 83.400 837.450 84.450 881.400 ;
        RECT 88.950 881.100 91.050 883.200 ;
        RECT 89.400 880.350 90.600 881.100 ;
        RECT 88.800 877.950 90.900 880.050 ;
        RECT 88.800 838.950 90.900 841.050 ;
        RECT 89.400 837.900 90.600 838.650 ;
        RECT 80.400 836.400 84.450 837.450 ;
        RECT 88.950 835.800 91.050 837.900 ;
        RECT 76.950 825.450 79.050 826.050 ;
        RECT 74.400 824.400 79.050 825.450 ;
        RECT 76.950 823.950 79.050 824.400 ;
        RECT 37.950 820.950 40.050 823.050 ;
        RECT 58.950 820.950 61.050 823.050 ;
        RECT 17.700 813.300 19.800 815.400 ;
        RECT 20.700 813.300 22.800 815.400 ;
        RECT 23.700 813.300 25.800 815.400 ;
        RECT 18.300 809.700 19.500 813.300 ;
        RECT 17.400 807.600 19.500 809.700 ;
        RECT 7.950 802.950 10.050 805.050 ;
        RECT 4.800 799.950 6.900 802.050 ;
        RECT 10.800 799.950 12.900 802.050 ;
        RECT 5.400 798.900 6.600 799.650 ;
        RECT 4.950 796.800 7.050 798.900 ;
        RECT 17.400 788.700 18.900 807.600 ;
        RECT 21.300 796.800 22.500 813.300 ;
        RECT 20.400 794.700 22.500 796.800 ;
        RECT 21.300 788.700 22.500 794.700 ;
        RECT 23.700 791.700 24.900 813.300 ;
        RECT 31.800 812.400 33.900 814.500 ;
        RECT 37.200 813.300 39.300 815.400 ;
        RECT 40.200 813.300 42.300 815.400 ;
        RECT 43.200 813.300 45.300 815.400 ;
        RECT 28.800 805.950 30.900 808.050 ;
        RECT 29.400 803.400 30.600 805.650 ;
        RECT 29.400 796.050 30.450 803.400 ;
        RECT 32.400 801.900 33.300 812.400 ;
        RECT 35.100 806.400 37.200 808.500 ;
        RECT 32.400 799.800 34.500 801.900 ;
        RECT 38.100 801.000 39.300 813.300 ;
        RECT 28.950 793.950 31.050 796.050 ;
        RECT 32.400 793.200 33.300 799.800 ;
        RECT 37.800 798.900 39.900 801.000 ;
        RECT 23.700 789.600 25.800 791.700 ;
        RECT 32.400 791.100 34.500 793.200 ;
        RECT 38.100 791.700 39.300 798.900 ;
        RECT 40.800 795.600 42.300 813.300 ;
        RECT 40.800 793.500 42.900 795.600 ;
        RECT 37.800 789.600 39.900 791.700 ;
        RECT 40.800 788.700 42.300 793.500 ;
        RECT 44.100 791.700 45.300 813.300 ;
        RECT 17.400 786.600 20.400 788.700 ;
        RECT 21.300 786.600 23.400 788.700 ;
        RECT 40.200 786.600 42.300 788.700 ;
        RECT 43.200 786.600 45.300 791.700 ;
        RECT 46.200 813.300 48.300 815.400 ;
        RECT 46.200 795.600 47.700 813.300 ;
        RECT 55.950 803.100 58.050 805.200 ;
        RECT 56.400 802.350 57.600 803.100 ;
        RECT 55.800 799.950 57.900 802.050 ;
        RECT 46.200 793.500 48.300 795.600 ;
        RECT 46.200 788.700 47.700 793.500 ;
        RECT 59.400 793.050 60.450 820.950 ;
        RECT 70.950 811.950 73.050 814.050 ;
        RECT 65.400 804.450 66.600 804.600 ;
        RECT 65.400 803.400 69.450 804.450 ;
        RECT 65.400 802.350 66.600 803.400 ;
        RECT 64.800 799.950 66.900 802.050 ;
        RECT 58.950 790.950 61.050 793.050 ;
        RECT 64.950 790.950 67.050 793.050 ;
        RECT 46.200 786.600 48.300 788.700 ;
        RECT 52.950 766.950 55.050 769.050 ;
        RECT 25.950 761.100 28.050 763.200 ;
        RECT 43.950 761.100 46.050 763.200 ;
        RECT 53.400 762.600 54.450 766.950 ;
        RECT 17.100 757.950 19.200 760.050 ;
        RECT 22.500 757.950 24.600 760.050 ;
        RECT 23.400 756.900 24.600 757.650 ;
        RECT 22.950 754.800 25.050 756.900 ;
        RECT 26.400 753.450 27.450 761.100 ;
        RECT 44.400 760.350 45.600 761.100 ;
        RECT 53.400 760.350 54.600 762.600 ;
        RECT 44.400 757.950 46.500 760.050 ;
        RECT 49.950 757.950 52.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 59.100 757.950 61.200 760.050 ;
        RECT 23.400 752.400 27.450 753.450 ;
        RECT 50.400 755.400 51.600 757.650 ;
        RECT 59.400 755.400 60.600 757.650 ;
        RECT 23.400 729.600 24.450 752.400 ;
        RECT 50.400 751.050 51.450 755.400 ;
        RECT 52.950 751.950 55.050 754.050 ;
        RECT 34.950 748.950 37.050 751.050 ;
        RECT 49.950 748.950 52.050 751.050 ;
        RECT 23.400 727.350 24.600 729.600 ;
        RECT 17.100 724.950 19.200 727.050 ;
        RECT 22.500 724.950 24.600 727.050 ;
        RECT 10.950 712.950 13.050 715.050 ;
        RECT 4.950 700.950 7.050 703.050 ;
        RECT 5.400 532.200 6.450 700.950 ;
        RECT 11.400 646.050 12.450 712.950 ;
        RECT 28.950 700.950 31.050 703.050 ;
        RECT 29.400 687.600 30.450 700.950 ;
        RECT 35.400 691.050 36.450 748.950 ;
        RECT 40.950 728.100 43.050 730.200 ;
        RECT 41.400 727.350 42.600 728.100 ;
        RECT 41.400 724.950 43.500 727.050 ;
        RECT 46.800 724.950 48.900 727.050 ;
        RECT 47.400 722.400 48.600 724.650 ;
        RECT 47.400 703.050 48.450 722.400 ;
        RECT 46.950 700.950 49.050 703.050 ;
        RECT 41.400 696.300 44.400 698.400 ;
        RECT 45.300 696.300 47.400 698.400 ;
        RECT 34.950 688.950 37.050 691.050 ;
        RECT 29.400 685.350 30.600 687.600 ;
        RECT 28.800 682.950 30.900 685.050 ;
        RECT 34.800 682.950 36.900 685.050 ;
        RECT 17.100 679.950 19.200 682.050 ;
        RECT 22.500 679.950 24.600 682.050 ;
        RECT 23.400 678.900 24.600 679.650 ;
        RECT 22.950 676.800 25.050 678.900 ;
        RECT 31.950 676.800 34.050 678.900 ;
        RECT 41.400 677.400 42.900 696.300 ;
        RECT 45.300 690.300 46.500 696.300 ;
        RECT 44.400 688.200 46.500 690.300 ;
        RECT 16.950 650.100 19.050 652.200 ;
        RECT 22.950 650.100 25.050 652.200 ;
        RECT 28.950 650.100 31.050 652.200 ;
        RECT 17.400 649.350 18.600 650.100 ;
        RECT 23.400 649.350 24.600 650.100 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 22.950 646.950 25.050 649.050 ;
        RECT 10.950 643.950 13.050 646.050 ;
        RECT 20.400 645.900 21.600 646.650 ;
        RECT 19.950 643.800 22.050 645.900 ;
        RECT 25.950 613.950 28.050 616.050 ;
        RECT 17.100 601.950 19.200 604.050 ;
        RECT 22.500 601.950 24.600 604.050 ;
        RECT 23.400 600.450 24.600 601.650 ;
        RECT 26.400 600.450 27.450 613.950 ;
        RECT 23.400 599.400 27.450 600.450 ;
        RECT 25.950 595.950 28.050 598.050 ;
        RECT 19.950 572.100 22.050 574.200 ;
        RECT 26.400 573.600 27.450 595.950 ;
        RECT 29.400 595.050 30.450 650.100 ;
        RECT 32.400 616.050 33.450 676.800 ;
        RECT 34.950 673.950 37.050 676.050 ;
        RECT 41.400 675.300 43.500 677.400 ;
        RECT 35.400 661.050 36.450 673.950 ;
        RECT 42.300 671.700 43.500 675.300 ;
        RECT 45.300 671.700 46.500 688.200 ;
        RECT 47.700 693.300 49.800 695.400 ;
        RECT 47.700 671.700 48.900 693.300 ;
        RECT 49.950 688.950 52.050 691.050 ;
        RECT 50.400 681.450 51.450 688.950 ;
        RECT 53.400 685.050 54.450 751.950 ;
        RECT 59.400 751.050 60.450 755.400 ;
        RECT 58.950 748.950 61.050 751.050 ;
        RECT 65.400 730.200 66.450 790.950 ;
        RECT 68.400 775.050 69.450 803.400 ;
        RECT 71.400 796.050 72.450 811.950 ;
        RECT 73.950 803.100 76.050 805.200 ;
        RECT 70.950 793.950 73.050 796.050 ;
        RECT 67.950 772.950 70.050 775.050 ;
        RECT 64.950 728.100 67.050 730.200 ;
        RECT 65.400 727.350 66.600 728.100 ;
        RECT 65.400 724.950 67.500 727.050 ;
        RECT 70.800 724.950 72.900 727.050 ;
        RECT 71.400 722.400 72.600 724.650 ;
        RECT 71.400 718.050 72.450 722.400 ;
        RECT 74.400 721.050 75.450 803.100 ;
        RECT 77.400 754.050 78.450 823.950 ;
        RECT 95.400 823.050 96.450 911.400 ;
        RECT 101.400 880.050 102.450 911.400 ;
        RECT 106.950 910.950 109.050 913.050 ;
        RECT 122.400 912.900 123.600 913.650 ;
        RECT 121.950 910.800 124.050 912.900 ;
        RECT 128.400 911.400 129.600 913.650 ;
        RECT 128.400 895.050 129.450 911.400 ;
        RECT 134.400 901.050 135.450 919.950 ;
        RECT 133.950 898.950 136.050 901.050 ;
        RECT 137.400 898.050 138.450 949.950 ;
        RECT 146.400 943.050 147.450 953.400 ;
        RECT 158.400 944.700 159.900 963.600 ;
        RECT 162.300 952.800 163.500 969.300 ;
        RECT 161.400 950.700 163.500 952.800 ;
        RECT 162.300 944.700 163.500 950.700 ;
        RECT 164.700 947.700 165.900 969.300 ;
        RECT 172.800 968.400 174.900 970.500 ;
        RECT 178.200 969.300 180.300 971.400 ;
        RECT 181.200 969.300 183.300 971.400 ;
        RECT 184.200 969.300 186.300 971.400 ;
        RECT 169.800 961.950 171.900 964.050 ;
        RECT 170.400 959.400 171.600 961.650 ;
        RECT 164.700 945.600 166.800 947.700 ;
        RECT 145.950 940.950 148.050 943.050 ;
        RECT 158.400 942.600 161.400 944.700 ;
        RECT 162.300 942.600 164.400 944.700 ;
        RECT 139.950 931.950 142.050 934.050 ;
        RECT 140.400 919.200 141.450 931.950 ;
        RECT 146.400 931.050 147.450 940.950 ;
        RECT 145.950 928.950 148.050 931.050 ;
        RECT 160.950 928.950 163.050 931.050 ;
        RECT 151.950 922.950 154.050 925.050 ;
        RECT 139.950 917.100 142.050 919.200 ;
        RECT 145.950 917.100 148.050 919.200 ;
        RECT 152.400 918.600 153.450 922.950 ;
        RECT 161.400 921.600 162.450 928.950 ;
        RECT 170.400 922.050 171.450 959.400 ;
        RECT 173.400 957.900 174.300 968.400 ;
        RECT 176.100 962.400 178.200 964.500 ;
        RECT 173.400 955.800 175.500 957.900 ;
        RECT 179.100 957.000 180.300 969.300 ;
        RECT 173.400 949.200 174.300 955.800 ;
        RECT 178.800 954.900 180.900 957.000 ;
        RECT 173.400 947.100 175.500 949.200 ;
        RECT 179.100 947.700 180.300 954.900 ;
        RECT 181.800 951.600 183.300 969.300 ;
        RECT 181.800 949.500 183.900 951.600 ;
        RECT 178.800 945.600 180.900 947.700 ;
        RECT 181.800 944.700 183.300 949.500 ;
        RECT 185.100 947.700 186.300 969.300 ;
        RECT 181.200 942.600 183.300 944.700 ;
        RECT 184.200 942.600 186.300 947.700 ;
        RECT 187.200 969.300 189.300 971.400 ;
        RECT 227.700 969.300 229.800 971.400 ;
        RECT 230.700 969.300 232.800 971.400 ;
        RECT 233.700 969.300 235.800 971.400 ;
        RECT 187.200 951.600 188.700 969.300 ;
        RECT 228.300 965.700 229.500 969.300 ;
        RECT 197.400 960.450 198.600 960.600 ;
        RECT 199.950 960.450 202.050 961.200 ;
        RECT 197.400 959.400 202.050 960.450 ;
        RECT 205.950 960.000 208.050 964.050 ;
        RECT 227.400 963.600 229.500 965.700 ;
        RECT 197.400 958.350 198.600 959.400 ;
        RECT 199.950 959.100 202.050 959.400 ;
        RECT 196.800 955.950 198.900 958.050 ;
        RECT 200.400 952.050 201.450 959.100 ;
        RECT 206.400 958.350 207.600 960.000 ;
        RECT 205.800 955.950 207.900 958.050 ;
        RECT 214.800 955.950 216.900 958.050 ;
        RECT 220.800 955.950 222.900 958.050 ;
        RECT 215.400 953.400 216.600 955.650 ;
        RECT 187.200 949.500 189.300 951.600 ;
        RECT 199.950 949.950 202.050 952.050 ;
        RECT 205.950 949.950 208.050 952.050 ;
        RECT 187.200 944.700 188.700 949.500 ;
        RECT 187.200 942.600 189.300 944.700 ;
        RECT 173.400 930.300 176.400 932.400 ;
        RECT 177.300 930.300 179.400 932.400 ;
        RECT 196.200 930.300 198.300 932.400 ;
        RECT 161.400 919.350 162.600 921.600 ;
        RECT 169.950 919.950 172.050 922.050 ;
        RECT 140.400 907.050 141.450 917.100 ;
        RECT 146.400 916.350 147.600 917.100 ;
        RECT 152.400 916.350 153.600 918.600 ;
        RECT 160.800 916.950 162.900 919.050 ;
        RECT 166.800 916.950 168.900 919.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 148.950 913.950 151.050 916.050 ;
        RECT 151.950 913.950 154.050 916.050 ;
        RECT 154.950 913.950 157.050 916.050 ;
        RECT 149.400 912.900 150.600 913.650 ;
        RECT 148.950 910.800 151.050 912.900 ;
        RECT 155.400 911.400 156.600 913.650 ;
        RECT 173.400 911.400 174.900 930.300 ;
        RECT 177.300 924.300 178.500 930.300 ;
        RECT 176.400 922.200 178.500 924.300 ;
        RECT 155.400 907.050 156.450 911.400 ;
        RECT 157.950 907.950 160.050 910.050 ;
        RECT 173.400 909.300 175.500 911.400 ;
        RECT 139.950 904.950 142.050 907.050 ;
        RECT 148.950 904.950 151.050 907.050 ;
        RECT 154.950 904.950 157.050 907.050 ;
        RECT 136.950 895.950 139.050 898.050 ;
        RECT 127.950 892.950 130.050 895.050 ;
        RECT 115.950 884.100 118.050 886.200 ;
        RECT 139.950 884.100 142.050 886.200 ;
        RECT 116.400 883.350 117.600 884.100 ;
        RECT 140.400 883.350 141.600 884.100 ;
        RECT 110.100 880.950 112.200 883.050 ;
        RECT 115.500 880.950 117.600 883.050 ;
        RECT 118.800 880.950 120.900 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 142.950 880.950 145.050 883.050 ;
        RECT 100.950 877.950 103.050 880.050 ;
        RECT 110.400 879.900 111.600 880.650 ;
        RECT 109.950 877.800 112.050 879.900 ;
        RECT 119.400 878.400 120.600 880.650 ;
        RECT 100.950 865.950 103.050 868.050 ;
        RECT 94.950 820.950 97.050 823.050 ;
        RECT 88.950 811.950 91.050 814.050 ;
        RECT 79.950 808.950 82.050 811.050 ;
        RECT 80.400 801.900 81.450 808.950 ;
        RECT 89.400 807.600 90.450 811.950 ;
        RECT 96.000 807.600 100.050 808.050 ;
        RECT 89.400 805.350 90.600 807.600 ;
        RECT 95.400 805.950 100.050 807.600 ;
        RECT 95.400 805.350 96.600 805.950 ;
        RECT 85.950 802.950 88.050 805.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 86.400 801.900 87.600 802.650 ;
        RECT 92.400 801.900 93.600 802.650 ;
        RECT 79.950 799.800 82.050 801.900 ;
        RECT 85.950 799.800 88.050 801.900 ;
        RECT 91.950 799.800 94.050 801.900 ;
        RECT 91.950 766.950 94.050 769.050 ;
        RECT 82.950 761.100 85.050 763.200 ;
        RECT 92.400 762.600 93.450 766.950 ;
        RECT 83.400 760.350 84.600 761.100 ;
        RECT 92.400 760.350 93.600 762.600 ;
        RECT 101.400 762.450 102.450 865.950 ;
        RECT 119.400 844.050 120.450 878.400 ;
        RECT 121.950 877.950 124.050 880.050 ;
        RECT 137.400 878.400 138.600 880.650 ;
        RECT 143.400 878.400 144.600 880.650 ;
        RECT 112.950 840.000 115.050 844.050 ;
        RECT 118.950 841.950 121.050 844.050 ;
        RECT 113.400 838.350 114.600 840.000 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 112.950 835.950 115.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 110.400 833.400 111.600 835.650 ;
        RECT 116.400 834.900 117.600 835.650 ;
        RECT 110.400 829.050 111.450 833.400 ;
        RECT 115.950 832.800 118.050 834.900 ;
        RECT 109.950 826.950 112.050 829.050 ;
        RECT 103.950 805.950 106.050 808.050 ;
        RECT 110.400 807.450 111.450 826.950 ;
        RECT 116.400 817.050 117.450 832.800 ;
        RECT 115.950 814.950 118.050 817.050 ;
        RECT 107.400 806.400 111.450 807.450 ;
        RECT 112.950 807.000 115.050 811.050 ;
        RECT 122.400 810.450 123.450 877.950 ;
        RECT 137.400 841.200 138.450 878.400 ;
        RECT 143.400 853.050 144.450 878.400 ;
        RECT 149.400 874.050 150.450 904.950 ;
        RECT 148.950 871.950 151.050 874.050 ;
        RECT 155.400 868.050 156.450 904.950 ;
        RECT 158.400 901.050 159.450 907.950 ;
        RECT 163.950 904.950 166.050 907.050 ;
        RECT 174.300 905.700 175.500 909.300 ;
        RECT 177.300 905.700 178.500 922.200 ;
        RECT 179.700 927.300 181.800 929.400 ;
        RECT 179.700 905.700 180.900 927.300 ;
        RECT 184.950 925.950 187.050 928.050 ;
        RECT 185.400 915.600 186.450 925.950 ;
        RECT 188.400 925.800 190.500 927.900 ;
        RECT 193.800 927.300 195.900 929.400 ;
        RECT 188.400 919.200 189.300 925.800 ;
        RECT 194.100 920.100 195.300 927.300 ;
        RECT 196.800 925.500 198.300 930.300 ;
        RECT 199.200 927.300 201.300 932.400 ;
        RECT 196.800 923.400 198.900 925.500 ;
        RECT 188.400 917.100 190.500 919.200 ;
        RECT 193.800 918.000 195.900 920.100 ;
        RECT 185.400 913.350 186.600 915.600 ;
        RECT 184.800 910.950 186.900 913.050 ;
        RECT 188.400 906.600 189.300 917.100 ;
        RECT 191.100 910.500 193.200 912.600 ;
        RECT 157.800 898.950 159.900 901.050 ;
        RECT 160.950 898.950 163.050 901.050 ;
        RECT 161.400 895.050 162.450 898.950 ;
        RECT 160.950 892.950 163.050 895.050 ;
        RECT 164.400 885.600 165.450 904.950 ;
        RECT 173.700 903.600 175.800 905.700 ;
        RECT 176.700 903.600 178.800 905.700 ;
        RECT 179.700 903.600 181.800 905.700 ;
        RECT 187.800 904.500 189.900 906.600 ;
        RECT 194.100 905.700 195.300 918.000 ;
        RECT 196.800 905.700 198.300 923.400 ;
        RECT 200.100 905.700 201.300 927.300 ;
        RECT 193.200 903.600 195.300 905.700 ;
        RECT 196.200 903.600 198.300 905.700 ;
        RECT 199.200 903.600 201.300 905.700 ;
        RECT 202.200 930.300 204.300 932.400 ;
        RECT 202.200 925.500 203.700 930.300 ;
        RECT 202.200 923.400 204.300 925.500 ;
        RECT 202.200 905.700 203.700 923.400 ;
        RECT 206.400 907.050 207.450 949.950 ;
        RECT 215.400 943.050 216.450 953.400 ;
        RECT 227.400 944.700 228.900 963.600 ;
        RECT 231.300 952.800 232.500 969.300 ;
        RECT 230.400 950.700 232.500 952.800 ;
        RECT 231.300 944.700 232.500 950.700 ;
        RECT 233.700 947.700 234.900 969.300 ;
        RECT 241.800 968.400 243.900 970.500 ;
        RECT 247.200 969.300 249.300 971.400 ;
        RECT 250.200 969.300 252.300 971.400 ;
        RECT 253.200 969.300 255.300 971.400 ;
        RECT 238.800 961.950 240.900 964.050 ;
        RECT 239.400 959.400 240.600 961.650 ;
        RECT 233.700 945.600 235.800 947.700 ;
        RECT 214.950 940.950 217.050 943.050 ;
        RECT 227.400 942.600 230.400 944.700 ;
        RECT 231.300 942.600 233.400 944.700 ;
        RECT 239.400 942.450 240.450 959.400 ;
        RECT 242.400 957.900 243.300 968.400 ;
        RECT 245.100 962.400 247.200 964.500 ;
        RECT 242.400 955.800 244.500 957.900 ;
        RECT 248.100 957.000 249.300 969.300 ;
        RECT 242.400 949.200 243.300 955.800 ;
        RECT 247.800 954.900 249.900 957.000 ;
        RECT 242.400 947.100 244.500 949.200 ;
        RECT 248.100 947.700 249.300 954.900 ;
        RECT 250.800 951.600 252.300 969.300 ;
        RECT 250.800 949.500 252.900 951.600 ;
        RECT 247.800 945.600 249.900 947.700 ;
        RECT 250.800 944.700 252.300 949.500 ;
        RECT 254.100 947.700 255.300 969.300 ;
        RECT 250.200 942.600 252.300 944.700 ;
        RECT 253.200 942.600 255.300 947.700 ;
        RECT 256.200 969.300 258.300 971.400 ;
        RECT 296.700 969.300 298.800 971.400 ;
        RECT 299.700 969.300 301.800 971.400 ;
        RECT 302.700 969.300 304.800 971.400 ;
        RECT 256.200 951.600 257.700 969.300 ;
        RECT 297.300 965.700 298.500 969.300 ;
        RECT 259.950 961.950 262.050 964.050 ;
        RECT 296.400 963.600 298.500 965.700 ;
        RECT 256.200 949.500 258.300 951.600 ;
        RECT 256.200 944.700 257.700 949.500 ;
        RECT 256.200 942.600 258.300 944.700 ;
        RECT 236.400 941.400 240.450 942.450 ;
        RECT 215.400 934.050 216.450 940.950 ;
        RECT 214.950 931.950 217.050 934.050 ;
        RECT 226.950 925.950 229.050 928.050 ;
        RECT 223.950 922.950 226.050 925.050 ;
        RECT 214.950 919.950 217.050 922.050 ;
        RECT 211.800 916.950 213.900 919.050 ;
        RECT 212.400 914.400 213.600 916.650 ;
        RECT 212.400 907.050 213.450 914.400 ;
        RECT 202.200 903.600 204.300 905.700 ;
        RECT 205.950 904.950 208.050 907.050 ;
        RECT 211.950 904.950 214.050 907.050 ;
        RECT 182.700 891.300 184.800 893.400 ;
        RECT 185.700 891.300 187.800 893.400 ;
        RECT 188.700 891.300 190.800 893.400 ;
        RECT 183.300 887.700 184.500 891.300 ;
        RECT 182.400 885.600 184.500 887.700 ;
        RECT 164.400 883.350 165.600 885.600 ;
        RECT 160.950 880.950 163.050 883.050 ;
        RECT 163.950 880.950 166.050 883.050 ;
        RECT 161.400 879.900 162.600 880.650 ;
        RECT 160.950 877.800 163.050 879.900 ;
        RECT 169.800 877.950 171.900 880.050 ;
        RECT 175.800 877.950 177.900 880.050 ;
        RECT 170.400 875.400 171.600 877.650 ;
        RECT 163.950 871.950 166.050 874.050 ;
        RECT 164.400 868.050 165.450 871.950 ;
        RECT 154.950 865.950 157.050 868.050 ;
        RECT 163.950 865.950 166.050 868.050 ;
        RECT 145.950 856.950 148.050 859.050 ;
        RECT 142.950 850.950 145.050 853.050 ;
        RECT 124.950 838.950 127.050 841.050 ;
        RECT 136.950 839.100 139.050 841.200 ;
        RECT 125.400 834.900 126.450 838.950 ;
        RECT 137.400 838.350 138.600 839.100 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 134.400 834.900 135.600 835.650 ;
        RECT 124.950 832.800 127.050 834.900 ;
        RECT 133.950 832.800 136.050 834.900 ;
        RECT 139.950 832.800 142.050 834.900 ;
        RECT 127.950 826.950 130.050 829.050 ;
        RECT 133.950 826.950 136.050 829.050 ;
        RECT 130.950 823.950 133.050 826.050 ;
        RECT 127.950 814.950 130.050 817.050 ;
        RECT 119.400 809.400 123.450 810.450 ;
        RECT 119.400 808.200 120.450 809.400 ;
        RECT 104.400 801.900 105.450 805.950 ;
        RECT 103.950 799.800 106.050 801.900 ;
        RECT 104.400 772.050 105.450 799.800 ;
        RECT 103.950 769.950 106.050 772.050 ;
        RECT 101.400 761.400 105.450 762.450 ;
        RECT 83.400 757.950 85.500 760.050 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 91.950 757.950 94.050 760.050 ;
        RECT 98.100 757.950 100.200 760.050 ;
        RECT 89.400 755.400 90.600 757.650 ;
        RECT 98.400 756.900 99.600 757.650 ;
        RECT 104.400 756.900 105.450 761.400 ;
        RECT 76.950 751.950 79.050 754.050 ;
        RECT 89.400 753.450 90.450 755.400 ;
        RECT 97.950 754.800 100.050 756.900 ;
        RECT 103.950 754.800 106.050 756.900 ;
        RECT 91.950 753.450 94.050 754.050 ;
        RECT 89.400 752.400 94.050 753.450 ;
        RECT 91.950 751.950 94.050 752.400 ;
        RECT 92.400 729.600 93.450 751.950 ;
        RECT 97.950 748.950 100.050 751.050 ;
        RECT 92.400 727.350 93.600 729.600 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 91.950 724.950 94.050 727.050 ;
        RECT 94.950 724.950 97.050 727.050 ;
        RECT 89.400 722.400 90.600 724.650 ;
        RECT 95.400 723.450 96.600 724.650 ;
        RECT 95.400 723.000 99.450 723.450 ;
        RECT 95.400 722.400 100.050 723.000 ;
        RECT 73.950 718.950 76.050 721.050 ;
        RECT 70.950 715.950 73.050 718.050 ;
        RECT 89.400 715.050 90.450 722.400 ;
        RECT 91.950 718.950 94.050 721.050 ;
        RECT 97.950 718.950 100.050 722.400 ;
        RECT 88.950 712.950 91.050 715.050 ;
        RECT 64.200 696.300 66.300 698.400 ;
        RECT 56.400 691.800 58.500 693.900 ;
        RECT 61.800 693.300 63.900 695.400 ;
        RECT 56.400 685.200 57.300 691.800 ;
        RECT 62.100 686.100 63.300 693.300 ;
        RECT 64.800 691.500 66.300 696.300 ;
        RECT 67.200 693.300 69.300 698.400 ;
        RECT 64.800 689.400 66.900 691.500 ;
        RECT 52.950 682.950 55.050 685.050 ;
        RECT 56.400 683.100 58.500 685.200 ;
        RECT 61.800 684.000 63.900 686.100 ;
        RECT 53.400 681.450 54.600 681.600 ;
        RECT 50.400 680.400 54.600 681.450 ;
        RECT 53.400 679.350 54.600 680.400 ;
        RECT 52.800 676.950 54.900 679.050 ;
        RECT 56.400 672.600 57.300 683.100 ;
        RECT 59.100 676.500 61.200 678.600 ;
        RECT 41.700 669.600 43.800 671.700 ;
        RECT 44.700 669.600 46.800 671.700 ;
        RECT 47.700 669.600 49.800 671.700 ;
        RECT 55.800 670.500 57.900 672.600 ;
        RECT 62.100 671.700 63.300 684.000 ;
        RECT 64.800 671.700 66.300 689.400 ;
        RECT 68.100 671.700 69.300 693.300 ;
        RECT 61.200 669.600 63.300 671.700 ;
        RECT 64.200 669.600 66.300 671.700 ;
        RECT 67.200 669.600 69.300 671.700 ;
        RECT 70.200 696.300 72.300 698.400 ;
        RECT 70.200 691.500 71.700 696.300 ;
        RECT 70.200 689.400 72.300 691.500 ;
        RECT 70.200 671.700 71.700 689.400 ;
        RECT 73.950 688.950 76.050 691.050 ;
        RECT 70.200 669.600 72.300 671.700 ;
        RECT 34.950 658.950 37.050 661.050 ;
        RECT 46.950 658.950 49.050 661.050 ;
        RECT 40.950 650.100 43.050 652.200 ;
        RECT 47.400 651.600 48.450 658.950 ;
        RECT 74.400 652.050 75.450 688.950 ;
        RECT 79.800 682.950 81.900 685.050 ;
        RECT 88.800 682.950 90.900 685.050 ;
        RECT 80.400 680.400 81.600 682.650 ;
        RECT 89.400 680.400 90.600 682.650 ;
        RECT 80.400 679.050 81.450 680.400 ;
        RECT 79.950 676.950 82.050 679.050 ;
        RECT 41.400 649.350 42.600 650.100 ;
        RECT 47.400 649.350 48.600 651.600 ;
        RECT 73.950 649.950 76.050 652.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 71.100 646.950 73.200 649.050 ;
        RECT 44.400 645.900 45.600 646.650 ;
        RECT 37.950 643.800 40.050 645.900 ;
        RECT 43.950 643.800 46.050 645.900 ;
        RECT 50.400 644.400 51.600 646.650 ;
        RECT 71.400 645.900 72.600 646.650 ;
        RECT 80.400 646.050 81.450 676.950 ;
        RECT 89.400 673.050 90.450 680.400 ;
        RECT 92.400 679.050 93.450 718.950 ;
        RECT 94.950 715.950 97.050 718.050 ;
        RECT 91.950 676.950 94.050 679.050 ;
        RECT 88.950 670.950 91.050 673.050 ;
        RECT 95.400 652.050 96.450 715.950 ;
        RECT 98.400 678.900 99.450 718.950 ;
        RECT 104.400 709.050 105.450 754.800 ;
        RECT 107.400 754.050 108.450 806.400 ;
        RECT 113.400 805.350 114.600 807.000 ;
        RECT 118.950 806.100 121.050 808.200 ;
        RECT 119.400 805.350 120.600 806.100 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 109.950 799.950 112.050 802.050 ;
        RECT 116.400 800.400 117.600 802.650 ;
        RECT 122.400 801.900 123.600 802.650 ;
        RECT 116.400 784.050 117.450 800.400 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 128.400 801.450 129.450 814.950 ;
        RECT 131.400 805.050 132.450 823.950 ;
        RECT 140.400 817.050 141.450 832.800 ;
        RECT 139.950 814.950 142.050 817.050 ;
        RECT 139.950 806.100 142.050 808.200 ;
        RECT 146.400 808.050 147.450 856.950 ;
        RECT 148.950 841.950 151.050 844.050 ;
        RECT 149.400 835.050 150.450 841.950 ;
        RECT 157.950 839.100 160.050 841.200 ;
        RECT 164.400 840.600 165.450 865.950 ;
        RECT 170.400 859.050 171.450 875.400 ;
        RECT 182.400 866.700 183.900 885.600 ;
        RECT 186.300 874.800 187.500 891.300 ;
        RECT 185.400 872.700 187.500 874.800 ;
        RECT 186.300 866.700 187.500 872.700 ;
        RECT 188.700 869.700 189.900 891.300 ;
        RECT 196.800 890.400 198.900 892.500 ;
        RECT 202.200 891.300 204.300 893.400 ;
        RECT 205.200 891.300 207.300 893.400 ;
        RECT 208.200 891.300 210.300 893.400 ;
        RECT 193.800 883.950 195.900 886.050 ;
        RECT 194.400 881.400 195.600 883.650 ;
        RECT 188.700 867.600 190.800 869.700 ;
        RECT 182.400 864.600 185.400 866.700 ;
        RECT 186.300 864.600 188.400 866.700 ;
        RECT 169.950 856.950 172.050 859.050 ;
        RECT 175.950 853.950 178.050 856.050 ;
        RECT 158.400 838.350 159.600 839.100 ;
        RECT 164.400 838.350 165.600 840.600 ;
        RECT 172.950 839.100 175.050 841.200 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 157.950 835.950 160.050 838.050 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 166.950 835.950 169.050 838.050 ;
        RECT 148.950 832.950 151.050 835.050 ;
        RECT 155.400 834.900 156.600 835.650 ;
        RECT 154.950 832.800 157.050 834.900 ;
        RECT 161.400 833.400 162.600 835.650 ;
        RECT 167.400 834.900 168.600 835.650 ;
        RECT 155.400 814.050 156.450 832.800 ;
        RECT 157.950 819.450 160.050 823.050 ;
        RECT 161.400 819.450 162.450 833.400 ;
        RECT 166.950 832.800 169.050 834.900 ;
        RECT 173.400 823.050 174.450 839.100 ;
        RECT 176.400 834.900 177.450 853.950 ;
        RECT 187.950 839.100 190.050 841.200 ;
        RECT 194.400 841.050 195.450 881.400 ;
        RECT 197.400 879.900 198.300 890.400 ;
        RECT 200.100 884.400 202.200 886.500 ;
        RECT 197.400 877.800 199.500 879.900 ;
        RECT 203.100 879.000 204.300 891.300 ;
        RECT 197.400 871.200 198.300 877.800 ;
        RECT 202.800 876.900 204.900 879.000 ;
        RECT 197.400 869.100 199.500 871.200 ;
        RECT 203.100 869.700 204.300 876.900 ;
        RECT 205.800 873.600 207.300 891.300 ;
        RECT 205.800 871.500 207.900 873.600 ;
        RECT 196.950 865.950 199.050 868.050 ;
        RECT 202.800 867.600 204.900 869.700 ;
        RECT 205.800 866.700 207.300 871.500 ;
        RECT 209.100 869.700 210.300 891.300 ;
        RECT 188.400 838.350 189.600 839.100 ;
        RECT 193.950 838.950 196.050 841.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 175.950 832.800 178.050 834.900 ;
        RECT 185.400 833.400 186.600 835.650 ;
        RECT 191.400 834.900 192.600 835.650 ;
        RECT 185.400 829.050 186.450 833.400 ;
        RECT 190.950 832.800 193.050 834.900 ;
        RECT 197.400 832.050 198.450 865.950 ;
        RECT 205.200 864.600 207.300 866.700 ;
        RECT 208.200 864.600 210.300 869.700 ;
        RECT 211.200 891.300 213.300 893.400 ;
        RECT 211.200 873.600 212.700 891.300 ;
        RECT 215.400 874.050 216.450 919.950 ;
        RECT 220.800 916.950 222.900 919.050 ;
        RECT 221.400 915.900 222.600 916.650 ;
        RECT 220.950 913.800 223.050 915.900 ;
        RECT 220.950 904.950 223.050 907.050 ;
        RECT 221.400 895.050 222.450 904.950 ;
        RECT 220.950 892.950 223.050 895.050 ;
        RECT 221.400 882.600 222.450 892.950 ;
        RECT 221.400 880.350 222.600 882.600 ;
        RECT 220.800 877.950 222.900 880.050 ;
        RECT 211.200 871.500 213.300 873.600 ;
        RECT 214.950 871.950 217.050 874.050 ;
        RECT 211.200 866.700 212.700 871.500 ;
        RECT 211.200 864.600 213.300 866.700 ;
        RECT 224.400 862.050 225.450 922.950 ;
        RECT 227.400 913.050 228.450 925.950 ;
        RECT 226.950 910.950 229.050 913.050 ;
        RECT 236.400 898.050 237.450 941.400 ;
        RECT 260.400 931.050 261.450 961.950 ;
        RECT 265.950 959.100 268.050 961.200 ;
        RECT 275.400 960.450 276.600 960.600 ;
        RECT 275.400 959.400 279.450 960.450 ;
        RECT 266.400 958.350 267.600 959.100 ;
        RECT 275.400 958.350 276.600 959.400 ;
        RECT 265.800 955.950 267.900 958.050 ;
        RECT 274.800 955.950 276.900 958.050 ;
        RECT 278.400 943.050 279.450 959.400 ;
        RECT 283.800 955.950 285.900 958.050 ;
        RECT 289.800 955.950 291.900 958.050 ;
        RECT 284.400 953.400 285.600 955.650 ;
        RECT 277.950 940.950 280.050 943.050 ;
        RECT 268.950 937.950 271.050 940.050 ;
        RECT 259.950 928.950 262.050 931.050 ;
        RECT 244.950 918.000 247.050 922.050 ;
        RECT 250.950 918.000 253.050 922.050 ;
        RECT 256.950 919.950 259.050 922.050 ;
        RECT 259.950 919.950 262.050 922.050 ;
        RECT 245.400 916.350 246.600 918.000 ;
        RECT 251.400 916.350 252.600 918.000 ;
        RECT 241.950 913.950 244.050 916.050 ;
        RECT 244.950 913.950 247.050 916.050 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 242.400 911.400 243.600 913.650 ;
        RECT 248.400 912.900 249.600 913.650 ;
        RECT 242.400 901.050 243.450 911.400 ;
        RECT 247.950 910.800 250.050 912.900 ;
        RECT 257.400 904.050 258.450 919.950 ;
        RECT 260.400 913.050 261.450 919.950 ;
        RECT 269.400 919.200 270.450 937.950 ;
        RECT 284.400 934.050 285.450 953.400 ;
        RECT 296.400 944.700 297.900 963.600 ;
        RECT 300.300 952.800 301.500 969.300 ;
        RECT 299.400 950.700 301.500 952.800 ;
        RECT 300.300 944.700 301.500 950.700 ;
        RECT 302.700 947.700 303.900 969.300 ;
        RECT 310.800 968.400 312.900 970.500 ;
        RECT 316.200 969.300 318.300 971.400 ;
        RECT 319.200 969.300 321.300 971.400 ;
        RECT 322.200 969.300 324.300 971.400 ;
        RECT 307.800 961.950 309.900 964.050 ;
        RECT 308.400 961.050 309.600 961.650 ;
        RECT 304.950 959.400 309.600 961.050 ;
        RECT 304.950 958.950 309.000 959.400 ;
        RECT 311.400 957.900 312.300 968.400 ;
        RECT 314.100 962.400 316.200 964.500 ;
        RECT 311.400 955.800 313.500 957.900 ;
        RECT 317.100 957.000 318.300 969.300 ;
        RECT 311.400 949.200 312.300 955.800 ;
        RECT 316.800 954.900 318.900 957.000 ;
        RECT 302.700 945.600 304.800 947.700 ;
        RECT 311.400 947.100 313.500 949.200 ;
        RECT 317.100 947.700 318.300 954.900 ;
        RECT 319.800 951.600 321.300 969.300 ;
        RECT 319.800 949.500 321.900 951.600 ;
        RECT 316.800 945.600 318.900 947.700 ;
        RECT 319.800 944.700 321.300 949.500 ;
        RECT 323.100 947.700 324.300 969.300 ;
        RECT 296.400 942.600 299.400 944.700 ;
        RECT 300.300 942.600 302.400 944.700 ;
        RECT 313.950 940.950 316.050 943.050 ;
        RECT 319.200 942.600 321.300 944.700 ;
        RECT 322.200 942.600 324.300 947.700 ;
        RECT 325.200 969.300 327.300 971.400 ;
        RECT 325.200 951.600 326.700 969.300 ;
        RECT 406.950 967.950 409.050 970.050 ;
        RECT 445.950 969.450 448.050 970.050 ;
        RECT 451.950 969.450 454.050 970.050 ;
        RECT 445.950 968.400 454.050 969.450 ;
        RECT 445.950 967.950 448.050 968.400 ;
        RECT 451.950 967.950 454.050 968.400 ;
        RECT 472.950 967.950 475.050 970.050 ;
        RECT 490.950 967.950 493.050 970.050 ;
        RECT 619.950 967.950 622.050 970.050 ;
        RECT 631.950 967.950 634.050 970.050 ;
        RECT 664.950 967.950 667.050 970.050 ;
        RECT 736.950 967.950 739.050 970.050 ;
        RECT 742.950 967.950 745.050 970.050 ;
        RECT 766.950 967.950 769.050 970.050 ;
        RECT 949.950 967.950 952.050 970.050 ;
        RECT 967.950 969.450 970.050 970.050 ;
        RECT 967.950 968.400 975.450 969.450 ;
        RECT 967.950 967.950 970.050 968.400 ;
        RECT 358.950 964.950 361.050 967.050 ;
        RECT 335.400 960.450 336.600 960.600 ;
        RECT 344.400 960.450 345.600 960.600 ;
        RECT 335.400 959.400 339.450 960.450 ;
        RECT 335.400 958.350 336.600 959.400 ;
        RECT 334.800 955.950 336.900 958.050 ;
        RECT 325.200 949.500 327.300 951.600 ;
        RECT 325.200 944.700 326.700 949.500 ;
        RECT 325.200 942.600 327.300 944.700 ;
        RECT 328.950 940.950 331.050 943.050 ;
        RECT 283.950 931.950 286.050 934.050 ;
        RECT 274.950 922.950 277.050 925.050 ;
        RECT 298.950 922.950 301.050 925.050 ;
        RECT 268.950 917.100 271.050 919.200 ;
        RECT 275.400 918.600 276.450 922.950 ;
        RECT 299.400 918.600 300.450 922.950 ;
        RECT 269.400 916.350 270.600 917.100 ;
        RECT 275.400 916.350 276.600 918.600 ;
        RECT 299.400 916.350 300.600 918.600 ;
        RECT 304.950 918.000 307.050 922.050 ;
        RECT 305.400 916.350 306.600 918.000 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 301.950 913.950 304.050 916.050 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 259.950 910.950 262.050 913.050 ;
        RECT 272.400 912.900 273.600 913.650 ;
        RECT 278.400 912.900 279.600 913.650 ;
        RECT 296.400 912.900 297.600 913.650 ;
        RECT 302.400 912.900 303.600 913.650 ;
        RECT 271.950 910.800 274.050 912.900 ;
        RECT 277.950 910.800 280.050 912.900 ;
        RECT 295.950 910.800 298.050 912.900 ;
        RECT 301.950 910.800 304.050 912.900 ;
        RECT 256.950 901.950 259.050 904.050 ;
        RECT 241.950 898.950 244.050 901.050 ;
        RECT 235.950 895.950 238.050 898.050 ;
        RECT 242.400 886.200 243.450 898.950 ;
        RECT 256.950 895.950 259.050 898.050 ;
        RECT 250.950 889.950 253.050 892.050 ;
        RECT 251.400 886.200 252.450 889.950 ;
        RECT 241.950 884.100 244.050 886.200 ;
        RECT 250.950 884.100 253.050 886.200 ;
        RECT 257.400 885.600 258.450 895.950 ;
        RECT 231.000 882.600 235.050 883.050 ;
        RECT 230.400 880.950 235.050 882.600 ;
        RECT 230.400 880.350 231.600 880.950 ;
        RECT 242.400 880.050 243.450 884.100 ;
        RECT 251.400 883.350 252.600 884.100 ;
        RECT 257.400 883.350 258.600 885.600 ;
        RECT 265.950 883.950 268.050 886.050 ;
        RECT 278.400 885.600 279.450 910.800 ;
        RECT 244.950 880.950 247.050 883.050 ;
        RECT 250.950 880.950 253.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 229.800 877.950 231.900 880.050 ;
        RECT 241.950 877.950 244.050 880.050 ;
        RECT 223.950 859.950 226.050 862.050 ;
        RECT 211.950 844.950 214.050 847.050 ;
        RECT 199.950 838.950 202.050 841.050 ;
        RECT 212.400 840.600 213.450 844.950 ;
        RECT 200.400 834.900 201.450 838.950 ;
        RECT 212.400 838.350 213.600 840.600 ;
        RECT 217.950 839.100 220.050 841.200 ;
        RECT 218.400 838.350 219.600 839.100 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 199.950 832.800 202.050 834.900 ;
        RECT 209.400 833.400 210.600 835.650 ;
        RECT 215.400 834.000 216.600 835.650 ;
        RECT 196.950 829.950 199.050 832.050 ;
        RECT 184.950 826.950 187.050 829.050 ;
        RECT 199.950 823.950 202.050 826.050 ;
        RECT 172.950 820.950 175.050 823.050 ;
        RECT 193.950 820.950 196.050 823.050 ;
        RECT 157.950 819.000 162.450 819.450 ;
        RECT 158.400 818.400 162.450 819.000 ;
        RECT 154.950 811.950 157.050 814.050 ;
        RECT 155.400 808.050 156.450 811.950 ;
        RECT 140.400 805.350 141.600 806.100 ;
        RECT 145.950 805.950 148.050 808.050 ;
        RECT 154.950 805.950 157.050 808.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 142.950 802.950 145.050 805.050 ;
        RECT 137.400 801.450 138.600 802.650 ;
        RECT 128.400 800.400 138.600 801.450 ;
        RECT 143.400 800.400 144.600 802.650 ;
        RECT 115.950 781.950 118.050 784.050 ;
        RECT 122.400 781.050 123.450 799.800 ;
        RECT 133.950 796.950 136.050 799.050 ;
        RECT 121.950 778.950 124.050 781.050 ;
        RECT 130.950 769.950 133.050 772.050 ;
        RECT 109.950 763.950 112.050 766.050 ;
        RECT 106.950 751.950 109.050 754.050 ;
        RECT 110.400 750.450 111.450 763.950 ;
        RECT 112.950 761.100 115.050 763.200 ;
        RECT 121.950 761.100 124.050 763.200 ;
        RECT 107.400 749.400 111.450 750.450 ;
        RECT 107.400 721.050 108.450 749.400 ;
        RECT 113.400 739.050 114.450 761.100 ;
        RECT 122.400 760.350 123.600 761.100 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 119.400 756.000 120.600 757.650 ;
        RECT 125.400 756.900 126.600 757.650 ;
        RECT 118.950 751.950 121.050 756.000 ;
        RECT 124.950 754.800 127.050 756.900 ;
        RECT 115.950 748.950 118.050 751.050 ;
        RECT 112.950 736.950 115.050 739.050 ;
        RECT 131.400 735.450 132.450 769.950 ;
        RECT 134.400 769.050 135.450 796.950 ;
        RECT 143.400 793.050 144.450 800.400 ;
        RECT 148.800 799.950 150.900 802.050 ;
        RECT 154.800 799.950 156.900 802.050 ;
        RECT 149.400 798.900 150.600 799.650 ;
        RECT 148.950 796.800 151.050 798.900 ;
        RECT 151.950 793.950 154.050 796.050 ;
        RECT 142.950 790.950 145.050 793.050 ;
        RECT 136.950 781.950 139.050 784.050 ;
        RECT 133.950 766.950 136.050 769.050 ;
        RECT 134.400 756.900 135.450 766.950 ;
        RECT 133.950 754.800 136.050 756.900 ;
        RECT 128.400 734.400 132.450 735.450 ;
        RECT 115.950 729.000 118.050 733.050 ;
        RECT 116.400 727.350 117.600 729.000 ;
        RECT 124.950 728.100 127.050 730.200 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 115.950 724.950 118.050 727.050 ;
        RECT 113.400 723.000 114.600 724.650 ;
        RECT 106.950 718.950 109.050 721.050 ;
        RECT 112.950 718.950 115.050 723.000 ;
        RECT 103.950 706.950 106.050 709.050 ;
        RECT 112.950 683.100 115.050 685.200 ;
        RECT 113.400 682.350 114.600 683.100 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 112.950 679.950 115.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 110.400 678.900 111.600 679.650 ;
        RECT 116.400 678.900 117.600 679.650 ;
        RECT 97.950 676.800 100.050 678.900 ;
        RECT 109.950 676.800 112.050 678.900 ;
        RECT 115.950 676.800 118.050 678.900 ;
        RECT 125.400 673.050 126.450 728.100 ;
        RECT 128.400 688.050 129.450 734.400 ;
        RECT 137.400 733.050 138.450 781.950 ;
        RECT 139.950 762.450 142.050 766.050 ;
        RECT 152.400 765.450 153.450 793.950 ;
        RECT 158.400 793.050 159.450 818.400 ;
        RECT 161.700 813.300 163.800 815.400 ;
        RECT 164.700 813.300 166.800 815.400 ;
        RECT 167.700 813.300 169.800 815.400 ;
        RECT 162.300 809.700 163.500 813.300 ;
        RECT 161.400 807.600 163.500 809.700 ;
        RECT 157.950 790.950 160.050 793.050 ;
        RECT 161.400 788.700 162.900 807.600 ;
        RECT 165.300 796.800 166.500 813.300 ;
        RECT 164.400 794.700 166.500 796.800 ;
        RECT 165.300 788.700 166.500 794.700 ;
        RECT 167.700 791.700 168.900 813.300 ;
        RECT 175.800 812.400 177.900 814.500 ;
        RECT 181.200 813.300 183.300 815.400 ;
        RECT 184.200 813.300 186.300 815.400 ;
        RECT 187.200 813.300 189.300 815.400 ;
        RECT 172.800 805.950 174.900 808.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 173.400 803.400 174.600 805.650 ;
        RECT 170.400 796.050 171.450 802.950 ;
        RECT 169.950 793.950 172.050 796.050 ;
        RECT 167.700 789.600 169.800 791.700 ;
        RECT 157.950 784.950 160.050 787.050 ;
        RECT 161.400 786.600 164.400 788.700 ;
        RECT 165.300 786.600 167.400 788.700 ;
        RECT 149.400 764.400 153.450 765.450 ;
        RECT 149.400 762.600 150.450 764.400 ;
        RECT 143.400 762.450 144.600 762.600 ;
        RECT 139.950 762.000 144.600 762.450 ;
        RECT 140.400 761.400 144.600 762.000 ;
        RECT 143.400 760.350 144.600 761.400 ;
        RECT 149.400 760.350 150.600 762.600 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 146.400 755.400 147.600 757.650 ;
        RECT 152.400 756.900 153.600 757.650 ;
        RECT 158.400 756.900 159.450 784.950 ;
        RECT 173.400 781.050 174.450 803.400 ;
        RECT 176.400 801.900 177.300 812.400 ;
        RECT 179.100 806.400 181.200 808.500 ;
        RECT 176.400 799.800 178.500 801.900 ;
        RECT 182.100 801.000 183.300 813.300 ;
        RECT 176.400 793.200 177.300 799.800 ;
        RECT 181.800 798.900 183.900 801.000 ;
        RECT 176.400 791.100 178.500 793.200 ;
        RECT 182.100 791.700 183.300 798.900 ;
        RECT 184.800 795.600 186.300 813.300 ;
        RECT 184.800 793.500 186.900 795.600 ;
        RECT 181.800 789.600 183.900 791.700 ;
        RECT 184.800 788.700 186.300 793.500 ;
        RECT 188.100 791.700 189.300 813.300 ;
        RECT 184.200 786.600 186.300 788.700 ;
        RECT 187.200 786.600 189.300 791.700 ;
        RECT 190.200 813.300 192.300 815.400 ;
        RECT 190.200 795.600 191.700 813.300 ;
        RECT 190.200 793.500 192.300 795.600 ;
        RECT 190.200 788.700 191.700 793.500 ;
        RECT 190.200 786.600 192.300 788.700 ;
        RECT 194.400 787.050 195.450 820.950 ;
        RECT 200.400 804.600 201.450 823.950 ;
        RECT 209.400 814.050 210.450 833.400 ;
        RECT 214.950 831.450 217.050 834.000 ;
        RECT 214.950 830.400 219.450 831.450 ;
        RECT 214.950 829.950 217.050 830.400 ;
        RECT 208.950 811.950 211.050 814.050 ;
        RECT 214.950 805.950 217.050 808.050 ;
        RECT 200.400 804.450 201.600 804.600 ;
        RECT 209.400 804.450 210.600 804.600 ;
        RECT 200.400 803.400 204.450 804.450 ;
        RECT 200.400 802.350 201.600 803.400 ;
        RECT 199.800 799.950 201.900 802.050 ;
        RECT 193.950 784.950 196.050 787.050 ;
        RECT 160.950 778.950 163.050 781.050 ;
        RECT 172.950 778.950 175.050 781.050 ;
        RECT 184.950 778.950 187.050 781.050 ;
        RECT 161.400 763.050 162.450 778.950 ;
        RECT 163.950 772.950 166.050 775.050 ;
        RECT 160.950 760.950 163.050 763.050 ;
        RECT 146.400 751.050 147.450 755.400 ;
        RECT 151.950 754.800 154.050 756.900 ;
        RECT 157.950 754.800 160.050 756.900 ;
        RECT 148.950 751.950 151.050 754.050 ;
        RECT 145.950 748.950 148.050 751.050 ;
        RECT 133.950 728.100 136.050 733.050 ;
        RECT 136.950 730.950 139.050 733.050 ;
        RECT 139.950 728.100 142.050 730.200 ;
        RECT 145.950 728.100 148.050 730.200 ;
        RECT 134.400 727.350 135.600 728.100 ;
        RECT 140.400 727.350 141.600 728.100 ;
        RECT 133.950 724.950 136.050 727.050 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 137.400 723.900 138.600 724.650 ;
        RECT 136.950 721.800 139.050 723.900 ;
        RECT 146.400 715.050 147.450 728.100 ;
        RECT 136.950 712.950 139.050 715.050 ;
        RECT 145.950 712.950 148.050 715.050 ;
        RECT 137.400 691.050 138.450 712.950 ;
        RECT 136.950 688.950 139.050 691.050 ;
        RECT 127.950 685.950 130.050 688.050 ;
        RECT 128.400 678.900 129.450 685.950 ;
        RECT 137.400 684.600 138.450 688.950 ;
        RECT 137.400 682.350 138.600 684.600 ;
        RECT 142.950 684.000 145.050 688.050 ;
        RECT 143.400 682.350 144.600 684.000 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 127.950 676.800 130.050 678.900 ;
        RECT 134.400 678.000 135.600 679.650 ;
        RECT 140.400 678.900 141.600 679.650 ;
        RECT 133.950 673.950 136.050 678.000 ;
        RECT 139.950 676.800 142.050 678.900 ;
        RECT 124.950 670.950 127.050 673.050 ;
        RECT 140.400 663.450 141.450 676.800 ;
        RECT 149.400 667.050 150.450 751.950 ;
        RECT 151.950 742.950 154.050 745.050 ;
        RECT 152.400 711.450 153.450 742.950 ;
        RECT 161.400 732.450 162.450 760.950 ;
        RECT 164.400 757.050 165.450 772.950 ;
        RECT 172.950 761.100 175.050 763.200 ;
        RECT 173.400 760.350 174.600 761.100 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 172.950 757.950 175.050 760.050 ;
        RECT 163.950 754.950 166.050 757.050 ;
        RECT 170.400 756.900 171.600 757.650 ;
        RECT 169.950 754.800 172.050 756.900 ;
        RECT 158.400 731.400 162.450 732.450 ;
        RECT 158.400 729.600 159.450 731.400 ;
        RECT 158.400 727.350 159.600 729.600 ;
        RECT 163.950 728.100 166.050 730.200 ;
        RECT 170.400 730.050 171.450 754.800 ;
        RECT 185.400 751.050 186.450 778.950 ;
        RECT 203.400 766.050 204.450 803.400 ;
        RECT 209.400 803.400 213.450 804.450 ;
        RECT 209.400 802.350 210.600 803.400 ;
        RECT 208.800 799.950 210.900 802.050 ;
        RECT 193.950 762.000 196.050 766.050 ;
        RECT 202.950 763.950 205.050 766.050 ;
        RECT 208.950 763.950 211.050 766.050 ;
        RECT 194.400 760.350 195.600 762.000 ;
        RECT 199.950 761.100 202.050 763.200 ;
        RECT 205.950 761.100 208.050 763.200 ;
        RECT 200.400 760.350 201.600 761.100 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 199.950 757.950 202.050 760.050 ;
        RECT 191.400 755.400 192.600 757.650 ;
        RECT 197.400 755.400 198.600 757.650 ;
        RECT 206.400 757.050 207.450 761.100 ;
        RECT 184.950 748.950 187.050 751.050 ;
        RECT 191.400 745.050 192.450 755.400 ;
        RECT 197.400 751.050 198.450 755.400 ;
        RECT 205.950 754.950 208.050 757.050 ;
        RECT 196.950 748.950 199.050 751.050 ;
        RECT 209.400 745.050 210.450 763.950 ;
        RECT 212.400 763.050 213.450 803.400 ;
        RECT 215.400 766.050 216.450 805.950 ;
        RECT 218.400 781.050 219.450 830.400 ;
        RECT 224.400 787.050 225.450 859.950 ;
        RECT 245.400 856.050 246.450 880.950 ;
        RECT 247.950 877.950 250.050 880.050 ;
        RECT 254.400 878.400 255.600 880.650 ;
        RECT 260.400 879.900 261.600 880.650 ;
        RECT 266.400 879.900 267.450 883.950 ;
        RECT 278.400 883.350 279.600 885.600 ;
        RECT 283.950 884.100 286.050 886.200 ;
        RECT 284.400 883.350 285.600 884.100 ;
        RECT 277.950 880.950 280.050 883.050 ;
        RECT 280.950 880.950 283.050 883.050 ;
        RECT 283.950 880.950 286.050 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 244.950 853.950 247.050 856.050 ;
        RECT 238.950 839.100 241.050 841.200 ;
        RECT 239.400 838.350 240.600 839.100 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 236.400 834.900 237.600 835.650 ;
        RECT 245.400 834.900 246.450 853.950 ;
        RECT 235.950 832.800 238.050 834.900 ;
        RECT 244.950 832.800 247.050 834.900 ;
        RECT 229.950 829.950 232.050 832.050 ;
        RECT 230.400 817.050 231.450 829.950 ;
        RECT 232.950 826.950 235.050 829.050 ;
        RECT 233.400 823.050 234.450 826.950 ;
        RECT 232.950 820.950 235.050 823.050 ;
        RECT 235.950 817.950 238.050 820.050 ;
        RECT 229.950 814.950 232.050 817.050 ;
        RECT 229.950 806.100 232.050 808.200 ;
        RECT 236.400 807.600 237.450 817.950 ;
        RECT 230.400 805.350 231.600 806.100 ;
        RECT 236.400 805.350 237.600 807.600 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 233.400 800.400 234.600 802.650 ;
        RECT 239.400 801.000 240.600 802.650 ;
        RECT 223.950 784.950 226.050 787.050 ;
        RECT 217.950 778.950 220.050 781.050 ;
        RECT 214.950 763.950 217.050 766.050 ;
        RECT 211.950 760.950 214.050 763.050 ;
        RECT 217.950 761.100 220.050 763.200 ;
        RECT 224.400 762.600 225.450 784.950 ;
        RECT 233.400 769.050 234.450 800.400 ;
        RECT 238.950 796.950 241.050 801.000 ;
        RECT 245.400 775.050 246.450 832.800 ;
        RECT 248.400 802.050 249.450 877.950 ;
        RECT 254.400 844.050 255.450 878.400 ;
        RECT 259.950 877.800 262.050 879.900 ;
        RECT 265.950 877.800 268.050 879.900 ;
        RECT 281.400 878.400 282.600 880.650 ;
        RECT 287.400 878.400 288.600 880.650 ;
        RECT 296.400 880.050 297.450 910.800 ;
        RECT 298.950 892.950 301.050 895.050 ;
        RECT 281.400 862.050 282.450 878.400 ;
        RECT 280.950 859.950 283.050 862.050 ;
        RECT 287.400 859.050 288.450 878.400 ;
        RECT 295.950 877.950 298.050 880.050 ;
        RECT 292.950 862.950 295.050 865.050 ;
        RECT 286.950 856.950 289.050 859.050 ;
        RECT 271.950 850.950 274.050 853.050 ;
        RECT 265.950 847.950 268.050 850.050 ;
        RECT 253.950 841.950 256.050 844.050 ;
        RECT 250.950 839.100 253.050 841.200 ;
        RECT 259.950 839.100 262.050 841.200 ;
        RECT 266.400 840.600 267.450 847.950 ;
        RECT 251.400 808.200 252.450 839.100 ;
        RECT 260.400 838.350 261.600 839.100 ;
        RECT 266.400 838.350 267.600 840.600 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 265.950 835.950 268.050 838.050 ;
        RECT 257.400 833.400 258.600 835.650 ;
        RECT 263.400 834.900 264.600 835.650 ;
        RECT 272.400 834.900 273.450 850.950 ;
        RECT 286.950 844.950 289.050 847.050 ;
        RECT 277.950 841.950 280.050 844.050 ;
        RECT 274.950 839.100 277.050 841.200 ;
        RECT 257.400 829.050 258.450 833.400 ;
        RECT 262.950 832.800 265.050 834.900 ;
        RECT 271.950 832.800 274.050 834.900 ;
        RECT 275.400 831.450 276.450 839.100 ;
        RECT 278.400 835.050 279.450 841.950 ;
        RECT 286.950 839.100 289.050 841.200 ;
        RECT 293.400 840.600 294.450 862.950 ;
        RECT 287.400 838.350 288.600 839.100 ;
        RECT 293.400 838.350 294.600 840.600 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 289.950 835.950 292.050 838.050 ;
        RECT 292.950 835.950 295.050 838.050 ;
        RECT 277.950 832.950 280.050 835.050 ;
        RECT 284.400 834.900 285.600 835.650 ;
        RECT 290.400 834.900 291.600 835.650 ;
        RECT 283.950 832.800 286.050 834.900 ;
        RECT 289.950 832.800 292.050 834.900 ;
        RECT 299.400 834.450 300.450 892.950 ;
        RECT 314.400 886.200 315.450 940.950 ;
        RECT 329.400 931.050 330.450 940.950 ;
        RECT 331.950 931.950 334.050 934.050 ;
        RECT 328.950 928.950 331.050 931.050 ;
        RECT 325.950 917.100 328.050 919.200 ;
        RECT 332.400 918.600 333.450 931.950 ;
        RECT 326.400 916.350 327.600 917.100 ;
        RECT 332.400 916.350 333.600 918.600 ;
        RECT 322.950 913.950 325.050 916.050 ;
        RECT 325.950 913.950 328.050 916.050 ;
        RECT 328.950 913.950 331.050 916.050 ;
        RECT 331.950 913.950 334.050 916.050 ;
        RECT 323.400 911.400 324.600 913.650 ;
        RECT 329.400 911.400 330.600 913.650 ;
        RECT 323.400 904.050 324.450 911.400 ;
        RECT 329.400 909.450 330.450 911.400 ;
        RECT 329.400 908.400 333.450 909.450 ;
        RECT 322.950 901.950 325.050 904.050 ;
        RECT 304.950 884.100 307.050 886.200 ;
        RECT 313.800 884.100 315.900 886.200 ;
        RECT 316.950 884.100 319.050 886.200 ;
        RECT 325.950 884.100 328.050 886.200 ;
        RECT 332.400 885.600 333.450 908.400 ;
        RECT 338.400 895.050 339.450 959.400 ;
        RECT 344.400 959.400 348.450 960.450 ;
        RECT 344.400 958.350 345.600 959.400 ;
        RECT 343.800 955.950 345.900 958.050 ;
        RECT 347.400 949.050 348.450 959.400 ;
        RECT 346.950 946.950 349.050 949.050 ;
        RECT 343.950 925.950 346.050 928.050 ;
        RECT 340.950 922.950 343.050 925.050 ;
        RECT 341.400 919.200 342.450 922.950 ;
        RECT 340.950 917.100 343.050 919.200 ;
        RECT 337.950 892.950 340.050 895.050 ;
        RECT 305.400 883.350 306.600 884.100 ;
        RECT 304.950 880.950 307.050 883.050 ;
        RECT 307.950 880.950 310.050 883.050 ;
        RECT 301.950 877.950 304.050 880.050 ;
        RECT 308.400 879.900 309.600 880.650 ;
        RECT 296.400 833.400 300.450 834.450 ;
        RECT 272.400 830.400 276.450 831.450 ;
        RECT 256.950 826.950 259.050 829.050 ;
        RECT 250.950 806.100 253.050 808.200 ;
        RECT 259.950 806.100 262.050 808.200 ;
        RECT 247.950 799.950 250.050 802.050 ;
        RECT 251.400 798.450 252.450 806.100 ;
        RECT 260.400 805.350 261.600 806.100 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 253.950 799.950 256.050 802.050 ;
        RECT 257.400 801.000 258.600 802.650 ;
        RECT 248.400 797.400 252.450 798.450 ;
        RECT 244.950 772.950 247.050 775.050 ;
        RECT 232.950 766.950 235.050 769.050 ;
        RECT 218.400 760.350 219.600 761.100 ;
        RECT 224.400 760.350 225.600 762.600 ;
        RECT 232.950 761.100 235.050 763.200 ;
        RECT 248.400 762.600 249.450 797.400 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 220.950 757.950 223.050 760.050 ;
        RECT 223.950 757.950 226.050 760.050 ;
        RECT 226.950 757.950 229.050 760.050 ;
        RECT 221.400 756.900 222.600 757.650 ;
        RECT 220.950 754.800 223.050 756.900 ;
        RECT 227.400 755.400 228.600 757.650 ;
        RECT 233.400 757.050 234.450 761.100 ;
        RECT 248.400 760.350 249.600 762.600 ;
        RECT 254.400 762.450 255.450 799.950 ;
        RECT 256.950 796.950 259.050 801.000 ;
        RECT 262.950 799.800 265.050 801.900 ;
        RECT 259.950 793.950 262.050 796.050 ;
        RECT 256.950 762.450 259.050 763.200 ;
        RECT 254.400 761.400 259.050 762.450 ;
        RECT 256.950 761.100 259.050 761.400 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 247.950 757.950 250.050 760.050 ;
        RECT 250.950 757.950 253.050 760.050 ;
        RECT 190.950 742.950 193.050 745.050 ;
        RECT 208.950 742.950 211.050 745.050 ;
        RECT 223.950 742.950 226.050 745.050 ;
        RECT 220.950 739.950 223.050 742.050 ;
        RECT 181.950 736.950 184.050 739.050 ;
        RECT 164.400 727.350 165.600 728.100 ;
        RECT 169.950 727.950 172.050 730.050 ;
        RECT 157.950 724.950 160.050 727.050 ;
        RECT 160.950 724.950 163.050 727.050 ;
        RECT 163.950 724.950 166.050 727.050 ;
        RECT 166.950 724.950 169.050 727.050 ;
        RECT 161.400 722.400 162.600 724.650 ;
        RECT 167.400 722.400 168.600 724.650 ;
        RECT 152.400 710.400 156.450 711.450 ;
        RECT 151.950 683.100 154.050 685.200 ;
        RECT 152.400 670.050 153.450 683.100 ;
        RECT 155.400 679.050 156.450 710.400 ;
        RECT 161.400 709.050 162.450 722.400 ;
        RECT 163.950 718.950 166.050 721.050 ;
        RECT 160.950 706.950 163.050 709.050 ;
        RECT 164.400 688.050 165.450 718.950 ;
        RECT 167.400 706.050 168.450 722.400 ;
        RECT 172.800 721.950 174.900 724.050 ;
        RECT 178.800 721.950 180.900 724.050 ;
        RECT 173.400 720.000 174.600 721.650 ;
        RECT 172.950 715.950 175.050 720.000 ;
        RECT 175.950 718.950 178.050 721.050 ;
        RECT 166.950 703.950 169.050 706.050 ;
        RECT 163.950 685.950 166.050 688.050 ;
        RECT 160.950 683.100 163.050 685.200 ;
        RECT 166.950 684.000 169.050 688.050 ;
        RECT 161.400 682.350 162.600 683.100 ;
        RECT 167.400 682.350 168.600 684.000 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 679.950 169.050 682.050 ;
        RECT 169.950 679.950 172.050 682.050 ;
        RECT 154.950 676.950 157.050 679.050 ;
        RECT 164.400 678.900 165.600 679.650 ;
        RECT 163.950 676.800 166.050 678.900 ;
        RECT 170.400 677.400 171.600 679.650 ;
        RECT 176.400 679.050 177.450 718.950 ;
        RECT 178.950 688.950 181.050 691.050 ;
        RECT 160.950 673.950 163.050 676.050 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 157.950 667.950 160.050 670.050 ;
        RECT 148.950 664.950 151.050 667.050 ;
        RECT 140.400 662.400 144.450 663.450 ;
        RECT 110.700 657.300 112.800 659.400 ;
        RECT 113.700 657.300 115.800 659.400 ;
        RECT 116.700 657.300 118.800 659.400 ;
        RECT 111.300 653.700 112.500 657.300 ;
        RECT 85.950 649.950 88.050 652.050 ;
        RECT 94.950 649.950 97.050 652.050 ;
        RECT 110.400 651.600 112.500 653.700 ;
        RECT 34.950 637.950 37.050 640.050 ;
        RECT 31.950 613.950 34.050 616.050 ;
        RECT 31.950 607.950 34.050 610.050 ;
        RECT 32.400 598.050 33.450 607.950 ;
        RECT 35.400 601.050 36.450 637.950 ;
        RECT 38.400 607.050 39.450 643.800 ;
        RECT 50.400 640.050 51.450 644.400 ;
        RECT 70.950 643.800 73.050 645.900 ;
        RECT 79.950 643.950 82.050 646.050 ;
        RECT 49.950 637.950 52.050 640.050 ;
        RECT 64.950 637.950 67.050 640.050 ;
        RECT 40.950 609.450 43.050 610.200 ;
        RECT 65.400 610.050 66.450 637.950 ;
        RECT 80.400 631.050 81.450 643.950 ;
        RECT 86.400 640.050 87.450 649.950 ;
        RECT 89.100 646.950 91.200 649.050 ;
        RECT 97.800 643.950 99.900 646.050 ;
        RECT 103.800 643.950 105.900 646.050 ;
        RECT 98.400 642.000 99.600 643.650 ;
        RECT 85.950 637.950 88.050 640.050 ;
        RECT 97.950 637.950 100.050 642.000 ;
        RECT 110.400 632.700 111.900 651.600 ;
        RECT 114.300 640.800 115.500 657.300 ;
        RECT 113.400 638.700 115.500 640.800 ;
        RECT 114.300 632.700 115.500 638.700 ;
        RECT 116.700 635.700 117.900 657.300 ;
        RECT 124.800 656.400 126.900 658.500 ;
        RECT 130.200 657.300 132.300 659.400 ;
        RECT 133.200 657.300 135.300 659.400 ;
        RECT 136.200 657.300 138.300 659.400 ;
        RECT 121.800 649.950 123.900 652.050 ;
        RECT 122.400 648.000 123.600 649.650 ;
        RECT 121.950 643.950 124.050 648.000 ;
        RECT 125.400 645.900 126.300 656.400 ;
        RECT 128.100 650.400 130.200 652.500 ;
        RECT 125.400 643.800 127.500 645.900 ;
        RECT 131.100 645.000 132.300 657.300 ;
        RECT 125.400 637.200 126.300 643.800 ;
        RECT 130.800 642.900 132.900 645.000 ;
        RECT 116.700 633.600 118.800 635.700 ;
        RECT 125.400 635.100 127.500 637.200 ;
        RECT 131.100 635.700 132.300 642.900 ;
        RECT 133.800 639.600 135.300 657.300 ;
        RECT 133.800 637.500 135.900 639.600 ;
        RECT 130.800 633.600 132.900 635.700 ;
        RECT 133.800 632.700 135.300 637.500 ;
        RECT 137.100 635.700 138.300 657.300 ;
        RECT 79.950 628.950 82.050 631.050 ;
        RECT 110.400 630.600 113.400 632.700 ;
        RECT 114.300 630.600 116.400 632.700 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 133.200 630.600 135.300 632.700 ;
        RECT 136.200 630.600 138.300 635.700 ;
        RECT 139.200 657.300 141.300 659.400 ;
        RECT 139.200 639.600 140.700 657.300 ;
        RECT 139.200 637.500 141.300 639.600 ;
        RECT 139.200 632.700 140.700 637.500 ;
        RECT 139.200 630.600 141.300 632.700 ;
        RECT 68.400 618.300 71.400 620.400 ;
        RECT 72.300 618.300 74.400 620.400 ;
        RECT 91.200 618.300 93.300 620.400 ;
        RECT 40.950 608.400 48.450 609.450 ;
        RECT 40.950 608.100 43.050 608.400 ;
        RECT 37.800 604.950 39.900 607.050 ;
        RECT 40.950 604.950 43.050 607.050 ;
        RECT 47.400 606.600 48.450 608.400 ;
        RECT 64.950 607.950 67.050 610.050 ;
        RECT 41.400 604.350 42.600 604.950 ;
        RECT 47.400 604.350 48.600 606.600 ;
        RECT 55.800 604.950 57.900 607.050 ;
        RECT 61.800 604.950 63.900 607.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 46.950 601.950 49.050 604.050 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 62.400 603.450 63.600 604.650 ;
        RECT 65.400 603.450 66.450 607.950 ;
        RECT 62.400 602.400 66.450 603.450 ;
        RECT 34.950 598.950 37.050 601.050 ;
        RECT 44.400 600.900 45.600 601.650 ;
        RECT 43.950 598.800 46.050 600.900 ;
        RECT 50.400 599.400 51.600 601.650 ;
        RECT 31.950 595.950 34.050 598.050 ;
        RECT 28.950 592.950 31.050 595.050 ;
        RECT 50.400 577.050 51.450 599.400 ;
        RECT 52.950 592.950 55.050 595.050 ;
        RECT 49.950 574.950 52.050 577.050 ;
        RECT 20.400 571.350 21.600 572.100 ;
        RECT 26.400 571.350 27.600 573.600 ;
        RECT 37.950 572.100 40.050 574.200 ;
        RECT 46.950 572.100 49.050 574.200 ;
        RECT 53.400 573.600 54.450 592.950 ;
        RECT 59.400 583.050 60.450 601.950 ;
        RECT 68.400 599.400 69.900 618.300 ;
        RECT 72.300 612.300 73.500 618.300 ;
        RECT 71.400 610.200 73.500 612.300 ;
        RECT 64.950 595.950 67.050 598.050 ;
        RECT 68.400 597.300 70.500 599.400 ;
        RECT 58.950 580.950 61.050 583.050 ;
        RECT 58.950 574.950 61.050 577.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 17.400 566.400 18.600 568.650 ;
        RECT 23.400 567.900 24.600 568.650 ;
        RECT 17.400 547.050 18.450 566.400 ;
        RECT 22.950 565.800 25.050 567.900 ;
        RECT 28.950 565.800 31.050 567.900 ;
        RECT 16.950 544.950 19.050 547.050 ;
        RECT 17.400 540.300 20.400 542.400 ;
        RECT 21.300 540.300 23.400 542.400 ;
        RECT 4.950 530.100 7.050 532.200 ;
        RECT 5.400 529.350 6.600 530.100 ;
        RECT 13.950 529.950 16.050 532.050 ;
        RECT 4.800 526.950 6.900 529.050 ;
        RECT 10.800 526.950 12.900 529.050 ;
        RECT 14.400 496.050 15.450 529.950 ;
        RECT 17.400 521.400 18.900 540.300 ;
        RECT 21.300 534.300 22.500 540.300 ;
        RECT 20.400 532.200 22.500 534.300 ;
        RECT 17.400 519.300 19.500 521.400 ;
        RECT 18.300 515.700 19.500 519.300 ;
        RECT 21.300 515.700 22.500 532.200 ;
        RECT 23.700 537.300 25.800 539.400 ;
        RECT 23.700 515.700 24.900 537.300 ;
        RECT 25.950 532.950 28.050 535.050 ;
        RECT 26.400 525.450 27.450 532.950 ;
        RECT 29.400 529.050 30.450 565.800 ;
        RECT 38.400 565.050 39.450 572.100 ;
        RECT 47.400 571.350 48.600 572.100 ;
        RECT 53.400 571.350 54.600 573.600 ;
        RECT 43.950 568.950 46.050 571.050 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 44.400 567.900 45.600 568.650 ;
        RECT 50.400 567.900 51.600 568.650 ;
        RECT 43.950 565.800 46.050 567.900 ;
        RECT 49.950 565.800 52.050 567.900 ;
        RECT 37.950 562.950 40.050 565.050 ;
        RECT 49.950 562.650 52.050 564.750 ;
        RECT 40.200 540.300 42.300 542.400 ;
        RECT 32.400 535.800 34.500 537.900 ;
        RECT 37.800 537.300 39.900 539.400 ;
        RECT 32.400 529.200 33.300 535.800 ;
        RECT 38.100 530.100 39.300 537.300 ;
        RECT 40.800 535.500 42.300 540.300 ;
        RECT 43.200 537.300 45.300 542.400 ;
        RECT 40.800 533.400 42.900 535.500 ;
        RECT 28.950 526.950 31.050 529.050 ;
        RECT 32.400 527.100 34.500 529.200 ;
        RECT 37.800 528.000 39.900 530.100 ;
        RECT 29.400 525.450 30.600 525.600 ;
        RECT 26.400 524.400 30.600 525.450 ;
        RECT 29.400 523.350 30.600 524.400 ;
        RECT 28.800 520.950 30.900 523.050 ;
        RECT 32.400 516.600 33.300 527.100 ;
        RECT 35.100 520.500 37.200 522.600 ;
        RECT 17.700 513.600 19.800 515.700 ;
        RECT 20.700 513.600 22.800 515.700 ;
        RECT 23.700 513.600 25.800 515.700 ;
        RECT 31.800 514.500 33.900 516.600 ;
        RECT 38.100 515.700 39.300 528.000 ;
        RECT 40.800 515.700 42.300 533.400 ;
        RECT 44.100 515.700 45.300 537.300 ;
        RECT 37.200 513.600 39.300 515.700 ;
        RECT 40.200 513.600 42.300 515.700 ;
        RECT 43.200 513.600 45.300 515.700 ;
        RECT 46.200 540.300 48.300 542.400 ;
        RECT 46.200 535.500 47.700 540.300 ;
        RECT 46.200 533.400 48.300 535.500 ;
        RECT 46.200 515.700 47.700 533.400 ;
        RECT 46.200 513.600 48.300 515.700 ;
        RECT 4.950 493.950 7.050 496.050 ;
        RECT 13.950 493.950 16.050 496.050 ;
        RECT 16.950 494.100 19.050 496.200 ;
        RECT 25.950 494.100 28.050 496.200 ;
        RECT 40.950 494.100 43.050 496.200 ;
        RECT 5.400 454.200 6.450 493.950 ;
        RECT 17.400 493.350 18.600 494.100 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 20.400 489.000 21.600 490.650 ;
        RECT 19.950 484.950 22.050 489.000 ;
        RECT 26.400 481.050 27.450 494.100 ;
        RECT 41.400 493.350 42.600 494.100 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 38.400 488.400 39.600 490.650 ;
        RECT 25.950 478.950 28.050 481.050 ;
        RECT 38.400 469.050 39.450 488.400 ;
        RECT 50.400 487.050 51.450 562.650 ;
        RECT 55.800 526.950 57.900 529.050 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 56.400 524.400 57.600 526.650 ;
        RECT 49.950 484.950 52.050 487.050 ;
        RECT 53.400 483.450 54.450 523.950 ;
        RECT 56.400 502.050 57.450 524.400 ;
        RECT 59.400 517.050 60.450 574.950 ;
        RECT 65.400 547.050 66.450 595.950 ;
        RECT 69.300 593.700 70.500 597.300 ;
        RECT 72.300 593.700 73.500 610.200 ;
        RECT 74.700 615.300 76.800 617.400 ;
        RECT 74.700 593.700 75.900 615.300 ;
        RECT 83.400 613.800 85.500 615.900 ;
        RECT 88.800 615.300 90.900 617.400 ;
        RECT 83.400 607.200 84.300 613.800 ;
        RECT 89.100 608.100 90.300 615.300 ;
        RECT 91.800 613.500 93.300 618.300 ;
        RECT 94.200 615.300 96.300 620.400 ;
        RECT 91.800 611.400 93.900 613.500 ;
        RECT 83.400 605.100 85.500 607.200 ;
        RECT 88.800 606.000 90.900 608.100 ;
        RECT 79.950 602.100 82.050 604.200 ;
        RECT 80.400 601.350 81.600 602.100 ;
        RECT 79.800 598.950 81.900 601.050 ;
        RECT 83.400 594.600 84.300 605.100 ;
        RECT 86.100 598.500 88.200 600.600 ;
        RECT 68.700 591.600 70.800 593.700 ;
        RECT 71.700 591.600 73.800 593.700 ;
        RECT 74.700 591.600 76.800 593.700 ;
        RECT 82.800 592.500 84.900 594.600 ;
        RECT 89.100 593.700 90.300 606.000 ;
        RECT 91.800 593.700 93.300 611.400 ;
        RECT 95.100 593.700 96.300 615.300 ;
        RECT 88.200 591.600 90.300 593.700 ;
        RECT 91.200 591.600 93.300 593.700 ;
        RECT 94.200 591.600 96.300 593.700 ;
        RECT 97.200 618.300 99.300 620.400 ;
        RECT 124.950 619.950 127.050 622.050 ;
        RECT 97.200 613.500 98.700 618.300 ;
        RECT 118.950 616.950 121.050 619.050 ;
        RECT 97.200 611.400 99.300 613.500 ;
        RECT 97.200 593.700 98.700 611.400 ;
        RECT 109.950 607.950 112.050 610.050 ;
        RECT 106.800 604.950 108.900 607.050 ;
        RECT 100.950 602.100 103.050 604.200 ;
        RECT 107.400 603.900 108.600 604.650 ;
        RECT 97.200 591.600 99.300 593.700 ;
        RECT 101.400 589.050 102.450 602.100 ;
        RECT 106.950 601.800 109.050 603.900 ;
        RECT 70.950 586.950 73.050 589.050 ;
        RECT 79.950 586.950 82.050 589.050 ;
        RECT 100.950 586.950 103.050 589.050 ;
        RECT 71.400 573.600 72.450 586.950 ;
        RECT 71.400 571.350 72.600 573.600 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 74.400 566.400 75.600 568.650 ;
        RECT 64.950 544.950 67.050 547.050 ;
        RECT 70.950 544.950 73.050 547.050 ;
        RECT 64.800 526.950 66.900 529.050 ;
        RECT 65.400 524.400 66.600 526.650 ;
        RECT 65.400 517.050 66.450 524.400 ;
        RECT 58.950 514.950 61.050 517.050 ;
        RECT 64.950 514.950 67.050 517.050 ;
        RECT 71.400 514.050 72.450 544.950 ;
        RECT 74.400 541.050 75.450 566.400 ;
        RECT 76.950 544.950 79.050 547.050 ;
        RECT 73.950 538.950 76.050 541.050 ;
        RECT 70.950 511.950 73.050 514.050 ;
        RECT 61.950 505.950 64.050 508.050 ;
        RECT 55.950 499.950 58.050 502.050 ;
        RECT 62.400 495.600 63.450 505.950 ;
        RECT 70.950 499.950 73.050 502.050 ;
        RECT 62.400 493.350 63.600 495.600 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 64.950 490.950 67.050 493.050 ;
        RECT 59.400 489.000 60.600 490.650 ;
        RECT 58.950 484.950 61.050 489.000 ;
        RECT 65.400 488.400 66.600 490.650 ;
        RECT 50.400 482.400 54.450 483.450 ;
        RECT 28.950 466.950 31.050 469.050 ;
        RECT 37.950 466.950 40.050 469.050 ;
        RECT 17.400 462.300 20.400 464.400 ;
        RECT 21.300 462.300 23.400 464.400 ;
        RECT 4.950 452.100 7.050 454.200 ;
        RECT 5.400 451.350 6.600 452.100 ;
        RECT 13.950 451.950 16.050 454.050 ;
        RECT 4.800 448.950 6.900 451.050 ;
        RECT 10.800 448.950 12.900 451.050 ;
        RECT 10.950 442.950 13.050 445.050 ;
        RECT 11.400 406.050 12.450 442.950 ;
        RECT 14.400 424.050 15.450 451.950 ;
        RECT 17.400 443.400 18.900 462.300 ;
        RECT 21.300 456.300 22.500 462.300 ;
        RECT 20.400 454.200 22.500 456.300 ;
        RECT 17.400 441.300 19.500 443.400 ;
        RECT 18.300 437.700 19.500 441.300 ;
        RECT 21.300 437.700 22.500 454.200 ;
        RECT 23.700 459.300 25.800 461.400 ;
        RECT 23.700 437.700 24.900 459.300 ;
        RECT 29.400 447.600 30.450 466.950 ;
        RECT 40.200 462.300 42.300 464.400 ;
        RECT 32.400 457.800 34.500 459.900 ;
        RECT 37.800 459.300 39.900 461.400 ;
        RECT 32.400 451.200 33.300 457.800 ;
        RECT 38.100 452.100 39.300 459.300 ;
        RECT 40.800 457.500 42.300 462.300 ;
        RECT 43.200 459.300 45.300 464.400 ;
        RECT 40.800 455.400 42.900 457.500 ;
        RECT 32.400 449.100 34.500 451.200 ;
        RECT 37.800 450.000 39.900 452.100 ;
        RECT 29.400 445.350 30.600 447.600 ;
        RECT 28.800 442.950 30.900 445.050 ;
        RECT 32.400 438.600 33.300 449.100 ;
        RECT 35.100 442.500 37.200 444.600 ;
        RECT 17.700 435.600 19.800 437.700 ;
        RECT 20.700 435.600 22.800 437.700 ;
        RECT 23.700 435.600 25.800 437.700 ;
        RECT 31.800 436.500 33.900 438.600 ;
        RECT 38.100 437.700 39.300 450.000 ;
        RECT 40.800 437.700 42.300 455.400 ;
        RECT 44.100 437.700 45.300 459.300 ;
        RECT 37.200 435.600 39.300 437.700 ;
        RECT 40.200 435.600 42.300 437.700 ;
        RECT 43.200 435.600 45.300 437.700 ;
        RECT 46.200 462.300 48.300 464.400 ;
        RECT 46.200 457.500 47.700 462.300 ;
        RECT 46.200 455.400 48.300 457.500 ;
        RECT 46.200 437.700 47.700 455.400 ;
        RECT 50.400 445.050 51.450 482.400 ;
        RECT 65.400 469.050 66.450 488.400 ;
        RECT 64.950 466.950 67.050 469.050 ;
        RECT 58.950 457.950 61.050 460.050 ;
        RECT 55.800 448.950 57.900 451.050 ;
        RECT 56.400 446.400 57.600 448.650 ;
        RECT 49.950 442.950 52.050 445.050 ;
        RECT 56.400 439.050 57.450 446.400 ;
        RECT 46.200 435.600 48.300 437.700 ;
        RECT 55.950 436.950 58.050 439.050 ;
        RECT 13.950 421.950 16.050 424.050 ;
        RECT 28.950 421.950 31.050 424.050 ;
        RECT 16.950 416.100 19.050 418.200 ;
        RECT 22.950 416.100 25.050 418.200 ;
        RECT 17.400 415.350 18.600 416.100 ;
        RECT 23.400 415.350 24.600 416.100 ;
        RECT 16.950 412.950 19.050 415.050 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 22.950 412.950 25.050 415.050 ;
        RECT 20.400 410.400 21.600 412.650 ;
        RECT 16.950 406.950 19.050 409.050 ;
        RECT 10.950 403.950 13.050 406.050 ;
        RECT 17.400 400.050 18.450 406.950 ;
        RECT 20.400 406.050 21.450 410.400 ;
        RECT 29.400 406.050 30.450 421.950 ;
        RECT 31.950 416.100 34.050 418.200 ;
        RECT 40.950 416.100 43.050 418.200 ;
        RECT 46.950 416.100 49.050 418.200 ;
        RECT 19.950 403.950 22.050 406.050 ;
        RECT 28.950 403.950 31.050 406.050 ;
        RECT 16.950 397.950 19.050 400.050 ;
        RECT 25.950 397.950 28.050 400.050 ;
        RECT 16.950 376.950 19.050 379.050 ;
        RECT 17.400 372.600 18.450 376.950 ;
        RECT 17.400 370.350 18.600 372.600 ;
        RECT 16.950 367.950 19.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 20.400 365.400 21.600 367.650 ;
        RECT 20.400 361.050 21.450 365.400 ;
        RECT 26.400 361.050 27.450 397.950 ;
        RECT 19.950 358.950 22.050 361.050 ;
        RECT 25.950 358.950 28.050 361.050 ;
        RECT 29.400 352.050 30.450 403.950 ;
        RECT 32.400 397.050 33.450 416.100 ;
        RECT 41.400 415.350 42.600 416.100 ;
        RECT 47.400 415.350 48.600 416.100 ;
        RECT 59.400 415.050 60.450 457.950 ;
        RECT 71.400 457.050 72.450 499.950 ;
        RECT 70.950 454.950 73.050 457.050 ;
        RECT 64.800 448.950 66.900 451.050 ;
        RECT 65.400 447.450 66.600 448.650 ;
        RECT 62.400 446.400 66.600 447.450 ;
        RECT 62.400 427.050 63.450 446.400 ;
        RECT 64.950 442.950 67.050 445.050 ;
        RECT 61.950 424.950 64.050 427.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 37.950 409.950 40.050 412.050 ;
        RECT 44.400 410.400 45.600 412.650 ;
        RECT 50.400 411.900 51.600 412.650 ;
        RECT 31.950 394.950 34.050 397.050 ;
        RECT 38.400 379.050 39.450 409.950 ;
        RECT 40.950 406.950 43.050 409.050 ;
        RECT 37.950 376.950 40.050 379.050 ;
        RECT 41.400 372.600 42.450 406.950 ;
        RECT 44.400 394.050 45.450 410.400 ;
        RECT 49.950 409.800 52.050 411.900 ;
        RECT 55.800 409.950 57.900 412.050 ;
        RECT 61.800 409.950 63.900 412.050 ;
        RECT 56.400 408.000 57.600 409.650 ;
        RECT 65.400 409.050 66.450 442.950 ;
        RECT 71.400 439.050 72.450 454.950 ;
        RECT 77.400 445.050 78.450 544.950 ;
        RECT 80.400 523.050 81.450 586.950 ;
        RECT 91.950 580.950 94.050 583.050 ;
        RECT 92.400 573.600 93.450 580.950 ;
        RECT 92.400 571.350 93.600 573.600 ;
        RECT 97.950 572.100 100.050 574.200 ;
        RECT 106.950 572.100 109.050 574.200 ;
        RECT 98.400 571.350 99.600 572.100 ;
        RECT 91.950 568.950 94.050 571.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 95.400 566.400 96.600 568.650 ;
        RECT 101.400 567.000 102.600 568.650 ;
        RECT 95.400 565.050 96.450 566.400 ;
        RECT 94.950 562.950 97.050 565.050 ;
        RECT 100.950 562.950 103.050 567.000 ;
        RECT 88.950 538.950 91.050 541.050 ;
        RECT 89.400 532.050 90.450 538.950 ;
        RECT 88.950 529.950 91.050 532.050 ;
        RECT 89.400 528.600 90.450 529.950 ;
        RECT 95.400 529.200 96.450 562.950 ;
        RECT 107.400 562.050 108.450 572.100 ;
        RECT 110.400 564.900 111.450 607.950 ;
        RECT 115.800 604.950 117.900 607.050 ;
        RECT 116.400 602.400 117.600 604.650 ;
        RECT 116.400 598.050 117.450 602.400 ;
        RECT 115.950 595.950 118.050 598.050 ;
        RECT 119.400 592.050 120.450 616.950 ;
        RECT 121.950 610.950 124.050 613.050 ;
        RECT 112.950 589.950 115.050 592.050 ;
        RECT 118.950 589.950 121.050 592.050 ;
        RECT 109.950 562.800 112.050 564.900 ;
        RECT 106.950 559.950 109.050 562.050 ;
        RECT 113.400 541.050 114.450 589.950 ;
        RECT 122.400 588.450 123.450 610.950 ;
        RECT 119.400 587.400 123.450 588.450 ;
        RECT 119.400 574.200 120.450 587.400 ;
        RECT 118.950 572.100 121.050 574.200 ;
        RECT 125.400 573.600 126.450 619.950 ;
        RECT 128.400 603.900 129.450 628.950 ;
        RECT 130.950 625.950 133.050 628.050 ;
        RECT 127.950 601.800 130.050 603.900 ;
        RECT 128.400 589.050 129.450 601.800 ;
        RECT 127.950 586.950 130.050 589.050 ;
        RECT 119.400 571.350 120.600 572.100 ;
        RECT 125.400 571.350 126.600 573.600 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 121.950 568.950 124.050 571.050 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 115.950 565.950 118.050 568.050 ;
        RECT 122.400 566.400 123.600 568.650 ;
        RECT 116.400 556.050 117.450 565.950 ;
        RECT 122.400 565.050 123.450 566.400 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 118.950 563.400 123.450 565.050 ;
        RECT 118.950 562.950 123.000 563.400 ;
        RECT 128.400 562.050 129.450 565.950 ;
        RECT 127.950 559.950 130.050 562.050 ;
        RECT 115.950 553.950 118.050 556.050 ;
        RECT 103.950 538.950 106.050 541.050 ;
        RECT 112.950 538.950 115.050 541.050 ;
        RECT 124.950 538.950 127.050 541.050 ;
        RECT 100.950 535.950 103.050 538.050 ;
        RECT 89.400 526.350 90.600 528.600 ;
        RECT 94.950 527.100 97.050 529.200 ;
        RECT 95.400 526.350 96.600 527.100 ;
        RECT 85.950 523.950 88.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 79.950 520.950 82.050 523.050 ;
        RECT 86.400 522.900 87.600 523.650 ;
        RECT 85.950 520.800 88.050 522.900 ;
        RECT 92.400 521.400 93.600 523.650 ;
        RECT 101.400 523.050 102.450 535.950 ;
        RECT 92.400 519.450 93.450 521.400 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 89.400 518.400 93.450 519.450 ;
        RECT 89.400 496.200 90.450 518.400 ;
        RECT 97.950 505.950 100.050 508.050 ;
        RECT 82.950 494.100 85.050 496.200 ;
        RECT 88.950 494.100 91.050 496.200 ;
        RECT 83.400 493.350 84.600 494.100 ;
        RECT 89.400 493.350 90.600 494.100 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 88.950 490.950 91.050 493.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 86.400 489.900 87.600 490.650 ;
        RECT 85.950 487.800 88.050 489.900 ;
        RECT 92.400 489.000 93.600 490.650 ;
        RECT 98.400 489.900 99.450 505.950 ;
        RECT 91.950 484.950 94.050 489.000 ;
        RECT 97.950 487.800 100.050 489.900 ;
        RECT 104.400 487.050 105.450 538.950 ;
        RECT 112.950 529.950 115.050 535.050 ;
        RECT 115.950 527.100 118.050 529.200 ;
        RECT 116.400 526.350 117.600 527.100 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 113.400 522.000 114.600 523.650 ;
        RECT 112.950 517.950 115.050 522.000 ;
        RECT 113.400 514.050 114.450 517.950 ;
        RECT 125.400 517.050 126.450 538.950 ;
        RECT 131.400 535.050 132.450 625.950 ;
        RECT 143.400 619.050 144.450 662.400 ;
        RECT 148.950 647.100 151.050 649.200 ;
        RECT 149.400 646.350 150.600 647.100 ;
        RECT 148.800 643.950 150.900 646.050 ;
        RECT 152.400 622.050 153.450 667.950 ;
        RECT 158.400 649.200 159.450 667.950 ;
        RECT 157.950 647.100 160.050 649.200 ;
        RECT 158.400 646.350 159.600 647.100 ;
        RECT 157.800 643.950 159.900 646.050 ;
        RECT 161.400 634.050 162.450 673.950 ;
        RECT 160.950 631.950 163.050 634.050 ;
        RECT 164.400 630.450 165.450 676.800 ;
        RECT 170.400 673.050 171.450 677.400 ;
        RECT 175.950 676.950 178.050 679.050 ;
        RECT 179.400 673.050 180.450 688.950 ;
        RECT 182.400 679.050 183.450 736.950 ;
        RECT 185.700 735.300 187.800 737.400 ;
        RECT 188.700 735.300 190.800 737.400 ;
        RECT 191.700 735.300 193.800 737.400 ;
        RECT 186.300 731.700 187.500 735.300 ;
        RECT 185.400 729.600 187.500 731.700 ;
        RECT 185.400 710.700 186.900 729.600 ;
        RECT 189.300 718.800 190.500 735.300 ;
        RECT 188.400 716.700 190.500 718.800 ;
        RECT 189.300 710.700 190.500 716.700 ;
        RECT 191.700 713.700 192.900 735.300 ;
        RECT 199.800 734.400 201.900 736.500 ;
        RECT 205.200 735.300 207.300 737.400 ;
        RECT 208.200 735.300 210.300 737.400 ;
        RECT 211.200 735.300 213.300 737.400 ;
        RECT 196.800 727.950 198.900 730.050 ;
        RECT 197.400 726.900 198.600 727.650 ;
        RECT 196.950 724.800 199.050 726.900 ;
        RECT 200.400 723.900 201.300 734.400 ;
        RECT 203.100 728.400 205.200 730.500 ;
        RECT 200.400 721.800 202.500 723.900 ;
        RECT 206.100 723.000 207.300 735.300 ;
        RECT 200.400 715.200 201.300 721.800 ;
        RECT 205.800 720.900 207.900 723.000 ;
        RECT 191.700 711.600 193.800 713.700 ;
        RECT 200.400 713.100 202.500 715.200 ;
        RECT 206.100 713.700 207.300 720.900 ;
        RECT 208.800 717.600 210.300 735.300 ;
        RECT 208.800 715.500 210.900 717.600 ;
        RECT 205.800 711.600 207.900 713.700 ;
        RECT 208.800 710.700 210.300 715.500 ;
        RECT 212.100 713.700 213.300 735.300 ;
        RECT 185.400 708.600 188.400 710.700 ;
        RECT 189.300 708.600 191.400 710.700 ;
        RECT 208.200 708.600 210.300 710.700 ;
        RECT 211.200 708.600 213.300 713.700 ;
        RECT 214.200 735.300 216.300 737.400 ;
        RECT 214.200 717.600 215.700 735.300 ;
        RECT 217.950 733.950 220.050 736.050 ;
        RECT 218.400 726.900 219.450 733.950 ;
        RECT 221.400 730.200 222.450 739.950 ;
        RECT 220.950 728.100 223.050 730.200 ;
        RECT 217.950 724.800 220.050 726.900 ;
        RECT 224.400 726.600 225.450 742.950 ;
        RECT 227.400 742.050 228.450 755.400 ;
        RECT 232.950 754.950 235.050 757.050 ;
        RECT 245.400 756.900 246.600 757.650 ;
        RECT 244.950 754.800 247.050 756.900 ;
        RECT 251.400 755.400 252.600 757.650 ;
        RECT 232.950 745.950 235.050 748.050 ;
        RECT 226.950 739.950 229.050 742.050 ;
        RECT 224.400 724.350 225.600 726.600 ;
        RECT 223.800 721.950 225.900 724.050 ;
        RECT 214.200 715.500 216.300 717.600 ;
        RECT 214.200 710.700 215.700 715.500 ;
        RECT 214.200 708.600 216.300 710.700 ;
        RECT 227.400 709.050 228.450 739.950 ;
        RECT 233.400 726.600 234.450 745.950 ;
        RECT 245.400 735.450 246.450 754.800 ;
        RECT 251.400 748.050 252.450 755.400 ;
        RECT 250.950 745.950 253.050 748.050 ;
        RECT 245.400 734.400 249.450 735.450 ;
        RECT 241.950 730.950 244.050 733.050 ;
        RECT 233.400 724.350 234.600 726.600 ;
        RECT 232.800 721.950 234.900 724.050 ;
        RECT 226.950 706.950 229.050 709.050 ;
        RECT 211.950 703.950 214.050 706.050 ;
        RECT 193.950 688.950 196.050 691.050 ;
        RECT 187.950 684.000 190.050 688.050 ;
        RECT 194.400 684.600 195.450 688.950 ;
        RECT 212.400 684.600 213.450 703.950 ;
        RECT 188.400 682.350 189.600 684.000 ;
        RECT 194.400 682.350 195.600 684.600 ;
        RECT 212.400 682.350 213.600 684.600 ;
        RECT 220.950 682.950 223.050 685.050 ;
        RECT 232.950 683.100 235.050 685.200 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 190.950 679.950 193.050 682.050 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 181.950 676.950 184.050 679.050 ;
        RECT 191.400 677.400 192.600 679.650 ;
        RECT 169.950 672.450 172.050 673.050 ;
        RECT 161.400 629.400 165.450 630.450 ;
        RECT 167.400 671.400 172.050 672.450 ;
        RECT 151.950 619.950 154.050 622.050 ;
        RECT 136.950 616.950 139.050 619.050 ;
        RECT 142.950 616.950 145.050 619.050 ;
        RECT 137.400 606.600 138.450 616.950 ;
        RECT 142.950 610.950 145.050 613.050 ;
        RECT 143.400 606.600 144.450 610.950 ;
        RECT 161.400 610.050 162.450 629.400 ;
        RECT 167.400 613.050 168.450 671.400 ;
        RECT 169.950 670.950 172.050 671.400 ;
        RECT 178.950 670.950 181.050 673.050 ;
        RECT 172.950 664.950 175.050 667.050 ;
        RECT 173.400 652.200 174.450 664.950 ;
        RECT 191.400 658.050 192.450 677.400 ;
        RECT 196.950 676.950 199.050 679.050 ;
        RECT 215.400 677.400 216.600 679.650 ;
        RECT 178.950 655.950 181.050 658.050 ;
        RECT 190.950 655.950 193.050 658.050 ;
        RECT 172.950 650.100 175.050 652.200 ;
        RECT 179.400 651.600 180.450 655.950 ;
        RECT 173.400 625.050 174.450 650.100 ;
        RECT 179.400 649.350 180.600 651.600 ;
        RECT 184.950 650.100 187.050 652.200 ;
        RECT 185.400 649.350 186.600 650.100 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 182.400 645.900 183.600 646.650 ;
        RECT 181.950 643.800 184.050 645.900 ;
        RECT 197.400 645.450 198.450 676.950 ;
        RECT 202.950 650.100 205.050 652.200 ;
        RECT 211.950 650.100 214.050 652.200 ;
        RECT 203.400 649.350 204.600 650.100 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 197.400 644.400 201.450 645.450 ;
        RECT 206.400 645.000 207.600 646.650 ;
        RECT 181.950 631.950 184.050 634.050 ;
        RECT 172.950 622.950 175.050 625.050 ;
        RECT 166.950 610.950 169.050 613.050 ;
        RECT 178.950 610.950 181.050 613.050 ;
        RECT 154.950 607.950 157.050 610.050 ;
        RECT 160.950 607.950 163.050 610.050 ;
        RECT 137.400 604.350 138.600 606.600 ;
        RECT 143.400 604.350 144.600 606.600 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 140.400 600.900 141.600 601.650 ;
        RECT 139.950 598.800 142.050 600.900 ;
        RECT 146.400 599.400 147.600 601.650 ;
        RECT 155.400 601.050 156.450 607.950 ;
        RECT 157.950 605.100 160.050 607.200 ;
        RECT 163.950 605.100 166.050 607.200 ;
        RECT 169.950 606.000 172.050 610.050 ;
        RECT 146.400 583.050 147.450 599.400 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 158.400 583.050 159.450 605.100 ;
        RECT 164.400 604.350 165.600 605.100 ;
        RECT 170.400 604.350 171.600 606.000 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 167.400 599.400 168.600 601.650 ;
        RECT 173.400 599.400 174.600 601.650 ;
        RECT 160.950 589.950 163.050 592.050 ;
        RECT 145.950 580.950 148.050 583.050 ;
        RECT 157.950 580.950 160.050 583.050 ;
        RECT 133.950 574.950 136.050 577.050 ;
        RECT 136.950 574.950 139.050 577.050 ;
        RECT 134.400 541.050 135.450 574.950 ;
        RECT 137.400 559.050 138.450 574.950 ;
        RECT 142.950 573.000 145.050 577.050 ;
        RECT 148.950 573.000 151.050 577.050 ;
        RECT 161.400 574.200 162.450 589.950 ;
        RECT 167.400 586.050 168.450 599.400 ;
        RECT 173.400 592.050 174.450 599.400 ;
        RECT 172.950 589.950 175.050 592.050 ;
        RECT 179.400 586.050 180.450 610.950 ;
        RECT 182.400 595.050 183.450 631.950 ;
        RECT 193.950 606.000 196.050 610.050 ;
        RECT 194.400 604.350 195.600 606.000 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 191.400 600.000 192.600 601.650 ;
        RECT 190.950 595.950 193.050 600.000 ;
        RECT 200.400 598.050 201.450 644.400 ;
        RECT 205.950 640.950 208.050 645.000 ;
        RECT 212.400 637.050 213.450 650.100 ;
        RECT 215.400 649.200 216.450 677.400 ;
        RECT 221.400 652.050 222.450 682.950 ;
        RECT 233.400 682.350 234.600 683.100 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 236.400 677.400 237.600 679.650 ;
        RECT 236.400 673.050 237.450 677.400 ;
        RECT 235.950 670.950 238.050 673.050 ;
        RECT 223.950 655.950 226.050 658.050 ;
        RECT 238.950 655.950 241.050 658.050 ;
        RECT 220.950 649.950 223.050 652.050 ;
        RECT 224.400 651.600 225.450 655.950 ;
        RECT 224.400 649.350 225.600 651.600 ;
        RECT 229.950 650.100 232.050 652.200 ;
        RECT 230.400 649.350 231.600 650.100 ;
        RECT 214.950 647.100 217.050 649.200 ;
        RECT 211.950 634.950 214.050 637.050 ;
        RECT 215.400 631.050 216.450 647.100 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 226.950 646.950 229.050 649.050 ;
        RECT 229.950 646.950 232.050 649.050 ;
        RECT 232.950 646.950 235.050 649.050 ;
        RECT 227.400 645.900 228.600 646.650 ;
        RECT 226.950 643.800 229.050 645.900 ;
        RECT 233.400 644.400 234.600 646.650 ;
        RECT 225.000 642.750 228.000 643.050 ;
        RECT 223.950 640.950 229.050 642.750 ;
        RECT 223.950 640.650 226.050 640.950 ;
        RECT 226.950 640.650 229.050 640.950 ;
        RECT 233.400 634.050 234.450 644.400 ;
        RECT 235.950 643.950 238.050 646.050 ;
        RECT 236.400 637.050 237.450 643.950 ;
        RECT 235.950 634.950 238.050 637.050 ;
        RECT 232.950 631.950 235.050 634.050 ;
        RECT 214.950 628.950 217.050 631.050 ;
        RECT 239.400 619.050 240.450 655.950 ;
        RECT 238.950 616.950 241.050 619.050 ;
        RECT 202.950 613.950 205.050 616.050 ;
        RECT 203.400 601.050 204.450 613.950 ;
        RECT 242.400 613.050 243.450 730.950 ;
        RECT 248.400 715.050 249.450 734.400 ;
        RECT 257.400 730.200 258.450 761.100 ;
        RECT 260.400 733.050 261.450 793.950 ;
        RECT 263.400 757.050 264.450 799.800 ;
        RECT 272.400 769.050 273.450 830.400 ;
        RECT 280.950 817.950 283.050 820.050 ;
        RECT 281.400 807.600 282.450 817.950 ;
        RECT 281.400 805.350 282.600 807.600 ;
        RECT 292.950 806.100 295.050 808.200 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 278.400 801.900 279.600 802.650 ;
        RECT 277.950 799.800 280.050 801.900 ;
        RECT 284.400 801.450 285.600 802.650 ;
        RECT 284.400 800.400 288.450 801.450 ;
        RECT 287.400 790.050 288.450 800.400 ;
        RECT 286.950 787.950 289.050 790.050 ;
        RECT 271.950 766.950 274.050 769.050 ;
        RECT 277.950 766.950 280.050 769.050 ;
        RECT 271.950 761.100 274.050 763.200 ;
        RECT 278.400 762.600 279.450 766.950 ;
        RECT 272.400 760.350 273.600 761.100 ;
        RECT 278.400 760.350 279.600 762.600 ;
        RECT 268.950 757.950 271.050 760.050 ;
        RECT 271.950 757.950 274.050 760.050 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 262.950 754.950 265.050 757.050 ;
        RECT 269.400 755.400 270.600 757.650 ;
        RECT 275.400 755.400 276.600 757.650 ;
        RECT 262.950 733.950 265.050 736.050 ;
        RECT 259.950 730.950 262.050 733.050 ;
        RECT 256.950 728.100 259.050 730.200 ;
        RECT 263.400 729.600 264.450 733.950 ;
        RECT 257.400 727.350 258.600 728.100 ;
        RECT 263.400 727.350 264.600 729.600 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 262.950 724.950 265.050 727.050 ;
        RECT 254.400 723.000 255.600 724.650 ;
        RECT 260.400 723.900 261.600 724.650 ;
        RECT 269.400 723.900 270.450 755.400 ;
        RECT 275.400 753.450 276.450 755.400 ;
        RECT 272.400 752.400 276.450 753.450 ;
        RECT 253.950 718.950 256.050 723.000 ;
        RECT 259.950 721.800 262.050 723.900 ;
        RECT 268.950 721.800 271.050 723.900 ;
        RECT 272.400 721.050 273.450 752.400 ;
        RECT 287.400 748.050 288.450 787.950 ;
        RECT 286.950 745.950 289.050 748.050 ;
        RECT 287.400 733.050 288.450 745.950 ;
        RECT 293.400 739.050 294.450 806.100 ;
        RECT 296.400 801.450 297.450 833.400 ;
        RECT 302.400 808.200 303.450 877.950 ;
        RECT 307.950 877.800 310.050 879.900 ;
        RECT 314.400 859.050 315.450 884.100 ;
        RECT 317.400 880.050 318.450 884.100 ;
        RECT 326.400 883.350 327.600 884.100 ;
        RECT 332.400 883.350 333.600 885.600 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 325.950 880.950 328.050 883.050 ;
        RECT 328.950 880.950 331.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 316.950 877.950 319.050 880.050 ;
        RECT 313.950 856.950 316.050 859.050 ;
        RECT 317.400 853.050 318.450 877.950 ;
        RECT 320.400 874.050 321.450 880.950 ;
        RECT 329.400 878.400 330.600 880.650 ;
        RECT 335.400 878.400 336.600 880.650 ;
        RECT 319.950 871.950 322.050 874.050 ;
        RECT 325.950 871.950 328.050 874.050 ;
        RECT 322.950 856.950 325.050 859.050 ;
        RECT 316.950 850.950 319.050 853.050 ;
        RECT 317.400 849.450 318.450 850.950 ;
        RECT 317.400 848.400 321.450 849.450 ;
        RECT 307.950 844.950 310.050 847.050 ;
        RECT 310.950 846.450 313.050 847.050 ;
        RECT 316.950 846.450 319.050 847.050 ;
        RECT 310.950 845.400 319.050 846.450 ;
        RECT 310.950 844.950 313.050 845.400 ;
        RECT 316.950 844.950 319.050 845.400 ;
        RECT 308.400 841.050 309.450 844.950 ;
        RECT 307.800 838.950 309.900 841.050 ;
        RECT 310.950 839.100 313.050 841.200 ;
        RECT 316.950 840.000 319.050 843.900 ;
        RECT 320.400 841.200 321.450 848.400 ;
        RECT 311.400 838.350 312.600 839.100 ;
        RECT 317.400 838.350 318.600 840.000 ;
        RECT 319.950 839.100 322.050 841.200 ;
        RECT 310.950 835.950 313.050 838.050 ;
        RECT 313.950 835.950 316.050 838.050 ;
        RECT 316.950 835.950 319.050 838.050 ;
        RECT 314.400 834.900 315.600 835.650 ;
        RECT 313.950 832.800 316.050 834.900 ;
        RECT 319.950 832.950 322.050 835.050 ;
        RECT 307.950 826.950 310.050 829.050 ;
        RECT 301.950 806.100 304.050 808.200 ;
        RECT 308.400 807.600 309.450 826.950 ;
        RECT 316.950 823.950 319.050 826.050 ;
        RECT 302.400 805.350 303.600 806.100 ;
        RECT 308.400 805.350 309.600 807.600 ;
        RECT 301.950 802.950 304.050 805.050 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 296.400 800.400 300.450 801.450 ;
        RECT 295.950 778.950 298.050 781.050 ;
        RECT 292.950 736.950 295.050 739.050 ;
        RECT 274.950 727.950 277.050 730.050 ;
        RECT 280.950 729.000 283.050 733.050 ;
        RECT 286.950 730.950 289.050 733.050 ;
        RECT 271.950 718.950 274.050 721.050 ;
        RECT 247.950 712.950 250.050 715.050 ;
        RECT 256.800 688.500 258.900 690.600 ;
        RECT 254.100 679.950 256.200 682.050 ;
        RECT 257.100 681.300 258.300 688.500 ;
        RECT 260.400 685.350 261.600 687.600 ;
        RECT 266.400 687.300 268.500 689.400 ;
        RECT 260.100 682.950 262.200 685.050 ;
        RECT 263.100 683.700 265.200 685.800 ;
        RECT 263.100 681.300 264.000 683.700 ;
        RECT 257.100 680.100 264.000 681.300 ;
        RECT 254.400 678.900 255.600 679.650 ;
        RECT 253.950 676.800 256.050 678.900 ;
        RECT 257.100 674.700 258.000 680.100 ;
        RECT 258.900 678.300 261.000 679.200 ;
        RECT 266.700 678.300 267.600 687.300 ;
        RECT 275.400 685.200 276.450 727.950 ;
        RECT 281.400 727.350 282.600 729.000 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 284.400 723.000 285.600 724.650 ;
        RECT 283.950 718.950 286.050 723.000 ;
        RECT 268.950 683.100 271.050 685.200 ;
        RECT 274.950 683.100 277.050 685.200 ;
        RECT 289.950 683.100 292.050 685.200 ;
        RECT 296.400 684.450 297.450 778.950 ;
        RECT 299.400 762.600 300.450 800.400 ;
        RECT 305.400 800.400 306.600 802.650 ;
        RECT 311.400 801.000 312.600 802.650 ;
        RECT 305.400 787.050 306.450 800.400 ;
        RECT 310.950 793.950 313.050 801.000 ;
        RECT 317.400 799.050 318.450 823.950 ;
        RECT 320.400 820.050 321.450 832.950 ;
        RECT 319.950 817.950 322.050 820.050 ;
        RECT 323.400 802.050 324.450 856.950 ;
        RECT 326.400 829.050 327.450 871.950 ;
        RECT 329.400 844.050 330.450 878.400 ;
        RECT 335.400 856.050 336.450 878.400 ;
        RECT 334.950 853.950 337.050 856.050 ;
        RECT 335.400 850.050 336.450 853.950 ;
        RECT 334.950 847.950 337.050 850.050 ;
        RECT 341.400 847.050 342.450 917.100 ;
        RECT 344.400 913.050 345.450 925.950 ;
        RECT 347.400 922.050 348.450 946.950 ;
        RECT 346.950 919.950 349.050 922.050 ;
        RECT 352.950 917.100 355.050 919.200 ;
        RECT 353.400 916.350 354.600 917.100 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 343.950 910.950 346.050 913.050 ;
        RECT 350.400 912.900 351.600 913.650 ;
        RECT 349.950 910.800 352.050 912.900 ;
        RECT 359.400 888.450 360.450 964.950 ;
        RECT 367.950 962.100 370.050 964.200 ;
        RECT 373.950 963.000 376.050 967.050 ;
        RECT 368.400 961.350 369.600 962.100 ;
        RECT 374.400 961.350 375.600 963.000 ;
        RECT 379.950 961.950 382.050 964.050 ;
        RECT 391.950 962.100 394.050 964.200 ;
        RECT 397.950 962.100 400.050 964.200 ;
        RECT 364.950 958.950 367.050 961.050 ;
        RECT 367.950 958.950 370.050 961.050 ;
        RECT 370.950 958.950 373.050 961.050 ;
        RECT 373.950 958.950 376.050 961.050 ;
        RECT 365.400 957.450 366.600 958.650 ;
        RECT 362.400 956.400 366.600 957.450 ;
        RECT 371.400 957.000 372.600 958.650 ;
        RECT 362.400 928.050 363.450 956.400 ;
        RECT 370.950 952.950 373.050 957.000 ;
        RECT 380.400 955.050 381.450 961.950 ;
        RECT 392.400 961.350 393.600 962.100 ;
        RECT 398.400 961.350 399.600 962.100 ;
        RECT 391.950 958.950 394.050 961.050 ;
        RECT 394.950 958.950 397.050 961.050 ;
        RECT 397.950 958.950 400.050 961.050 ;
        RECT 400.950 958.950 403.050 961.050 ;
        RECT 395.400 957.900 396.600 958.650 ;
        RECT 394.950 955.800 397.050 957.900 ;
        RECT 401.400 956.400 402.600 958.650 ;
        RECT 407.400 957.900 408.450 967.950 ;
        RECT 421.950 962.100 424.050 964.200 ;
        RECT 422.400 961.350 423.600 962.100 ;
        RECT 430.950 961.950 433.050 964.050 ;
        RECT 442.950 962.100 445.050 964.200 ;
        RECT 448.950 962.100 451.050 967.050 ;
        RECT 473.400 963.600 474.450 967.950 ;
        RECT 418.950 958.950 421.050 961.050 ;
        RECT 421.950 958.950 424.050 961.050 ;
        RECT 424.950 958.950 427.050 961.050 ;
        RECT 379.950 952.950 382.050 955.050 ;
        RECT 364.950 937.950 367.050 940.050 ;
        RECT 365.400 931.050 366.450 937.950 ;
        RECT 364.950 928.950 367.050 931.050 ;
        RECT 361.950 925.950 364.050 928.050 ;
        RECT 365.400 912.900 366.450 928.950 ;
        RECT 401.400 925.050 402.450 956.400 ;
        RECT 406.950 955.800 409.050 957.900 ;
        RECT 419.400 957.450 420.600 958.650 ;
        RECT 425.400 957.900 426.600 958.650 ;
        RECT 416.400 956.400 420.600 957.450 ;
        RECT 416.400 952.050 417.450 956.400 ;
        RECT 424.950 955.800 427.050 957.900 ;
        RECT 415.950 949.950 418.050 952.050 ;
        RECT 379.950 922.950 382.050 925.050 ;
        RECT 400.950 922.950 403.050 925.050 ;
        RECT 406.950 922.950 409.050 925.050 ;
        RECT 373.950 918.000 376.050 922.050 ;
        RECT 380.400 918.600 381.450 922.950 ;
        RECT 388.950 919.950 391.050 922.050 ;
        RECT 374.400 916.350 375.600 918.000 ;
        RECT 380.400 916.350 381.600 918.600 ;
        RECT 385.950 916.950 388.050 919.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 373.950 913.950 376.050 916.050 ;
        RECT 376.950 913.950 379.050 916.050 ;
        RECT 379.950 913.950 382.050 916.050 ;
        RECT 364.950 910.800 367.050 912.900 ;
        RECT 371.400 911.400 372.600 913.650 ;
        RECT 377.400 912.900 378.600 913.650 ;
        RECT 386.400 912.900 387.450 916.950 ;
        RECT 371.400 907.050 372.450 911.400 ;
        RECT 376.950 910.800 379.050 912.900 ;
        RECT 385.950 910.800 388.050 912.900 ;
        RECT 367.950 905.400 372.450 907.050 ;
        RECT 367.950 904.950 372.000 905.400 ;
        RECT 389.400 904.050 390.450 919.950 ;
        RECT 407.400 918.600 408.450 922.950 ;
        RECT 416.400 918.600 417.450 949.950 ;
        RECT 425.400 949.050 426.450 955.800 ;
        RECT 424.950 946.950 427.050 949.050 ;
        RECT 421.950 937.950 424.050 940.050 ;
        RECT 418.950 922.950 421.050 925.050 ;
        RECT 407.400 916.350 408.600 918.600 ;
        RECT 416.400 916.350 417.600 918.600 ;
        RECT 400.800 913.950 402.900 916.050 ;
        RECT 406.950 913.950 409.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 415.500 913.950 417.600 916.050 ;
        RECT 401.400 912.900 402.600 913.650 ;
        RECT 410.400 912.900 411.600 913.650 ;
        RECT 400.950 910.800 403.050 912.900 ;
        RECT 397.950 907.950 400.050 910.050 ;
        RECT 388.950 901.950 391.050 904.050 ;
        RECT 394.950 898.950 397.050 901.050 ;
        RECT 385.950 889.950 388.050 892.050 ;
        RECT 361.950 888.450 364.050 889.050 ;
        RECT 359.400 887.400 364.050 888.450 ;
        RECT 355.950 884.100 358.050 886.200 ;
        RECT 361.950 885.000 364.050 887.400 ;
        RECT 356.400 883.350 357.600 884.100 ;
        RECT 362.400 883.350 363.600 885.000 ;
        RECT 367.950 883.950 370.050 886.050 ;
        RECT 379.950 884.100 382.050 886.200 ;
        RECT 386.400 885.600 387.450 889.950 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 361.950 880.950 364.050 883.050 ;
        RECT 353.400 878.400 354.600 880.650 ;
        RECT 359.400 879.900 360.600 880.650 ;
        RECT 368.400 879.900 369.450 883.950 ;
        RECT 380.400 883.350 381.600 884.100 ;
        RECT 386.400 883.350 387.600 885.600 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 382.950 880.950 385.050 883.050 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 353.400 874.050 354.450 878.400 ;
        RECT 358.950 877.800 361.050 879.900 ;
        RECT 367.950 877.800 370.050 879.900 ;
        RECT 383.400 878.400 384.600 880.650 ;
        RECT 389.400 879.900 390.600 880.650 ;
        RECT 352.950 871.950 355.050 874.050 ;
        RECT 376.950 871.950 379.050 874.050 ;
        RECT 355.950 868.950 358.050 871.050 ;
        RECT 343.950 865.950 346.050 868.050 ;
        RECT 344.400 859.050 345.450 865.950 ;
        RECT 356.400 865.050 357.450 868.950 ;
        RECT 355.950 862.950 358.050 865.050 ;
        RECT 343.950 856.950 346.050 859.050 ;
        RECT 336.000 846.900 339.000 847.050 ;
        RECT 334.950 846.450 339.000 846.900 ;
        RECT 334.950 844.950 339.450 846.450 ;
        RECT 340.950 844.950 343.050 847.050 ;
        RECT 334.950 844.800 337.050 844.950 ;
        RECT 328.950 841.950 331.050 844.050 ;
        RECT 338.400 843.450 339.450 844.950 ;
        RECT 338.400 842.400 342.450 843.450 ;
        RECT 329.400 835.050 330.450 841.950 ;
        RECT 341.400 841.200 342.450 842.400 ;
        RECT 334.950 839.100 337.050 841.200 ;
        RECT 340.950 839.100 343.050 841.200 ;
        RECT 335.400 838.350 336.600 839.100 ;
        RECT 341.400 838.350 342.600 839.100 ;
        RECT 334.950 835.950 337.050 838.050 ;
        RECT 337.950 835.950 340.050 838.050 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 352.950 835.950 355.050 838.050 ;
        RECT 328.950 832.950 331.050 835.050 ;
        RECT 338.400 833.400 339.600 835.650 ;
        RECT 344.400 834.900 345.600 835.650 ;
        RECT 328.950 829.800 331.050 831.900 ;
        RECT 325.950 826.950 328.050 829.050 ;
        RECT 329.400 823.050 330.450 829.800 ;
        RECT 328.950 820.950 331.050 823.050 ;
        RECT 329.400 807.600 330.450 820.950 ;
        RECT 329.400 805.350 330.600 807.600 ;
        RECT 335.400 807.450 336.600 807.600 ;
        RECT 338.400 807.450 339.450 833.400 ;
        RECT 343.950 832.800 346.050 834.900 ;
        RECT 353.400 823.050 354.450 835.950 ;
        RECT 352.950 820.950 355.050 823.050 ;
        RECT 356.400 820.050 357.450 862.950 ;
        RECT 373.950 859.950 376.050 862.050 ;
        RECT 364.950 839.100 367.050 841.200 ;
        RECT 365.400 838.350 366.600 839.100 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 362.400 834.000 363.600 835.650 ;
        RECT 361.950 829.950 364.050 834.000 ;
        RECT 368.400 833.400 369.600 835.650 ;
        RECT 374.400 834.900 375.450 859.950 ;
        RECT 362.400 826.050 363.450 829.950 ;
        RECT 361.950 823.950 364.050 826.050 ;
        RECT 368.400 823.050 369.450 833.400 ;
        RECT 373.950 832.800 376.050 834.900 ;
        RECT 377.400 832.050 378.450 871.950 ;
        RECT 383.400 844.050 384.450 878.400 ;
        RECT 388.950 877.800 391.050 879.900 ;
        RECT 395.400 874.050 396.450 898.950 ;
        RECT 394.950 871.950 397.050 874.050 ;
        RECT 398.400 871.050 399.450 907.950 ;
        RECT 401.400 886.200 402.450 910.800 ;
        RECT 409.950 907.950 412.050 912.900 ;
        RECT 412.950 889.950 415.050 892.050 ;
        RECT 400.950 884.100 403.050 886.200 ;
        RECT 406.950 884.100 409.050 886.200 ;
        RECT 413.400 885.600 414.450 889.950 ;
        RECT 397.950 868.950 400.050 871.050 ;
        RECT 394.950 865.950 397.050 868.050 ;
        RECT 385.950 859.950 388.050 862.050 ;
        RECT 382.950 841.950 385.050 844.050 ;
        RECT 386.400 840.600 387.450 859.950 ;
        RECT 395.400 859.050 396.450 865.950 ;
        RECT 394.950 856.950 397.050 859.050 ;
        RECT 386.400 838.350 387.600 840.600 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 389.400 834.900 390.600 835.650 ;
        RECT 395.400 834.900 396.450 856.950 ;
        RECT 401.400 856.050 402.450 884.100 ;
        RECT 407.400 883.350 408.600 884.100 ;
        RECT 413.400 883.350 414.600 885.600 ;
        RECT 419.400 885.450 420.450 922.950 ;
        RECT 422.400 901.050 423.450 937.950 ;
        RECT 421.950 898.950 424.050 901.050 ;
        RECT 419.400 884.400 423.450 885.450 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 410.400 878.400 411.600 880.650 ;
        RECT 416.400 879.900 417.600 880.650 ;
        RECT 422.400 879.900 423.450 884.400 ;
        RECT 410.400 871.050 411.450 878.400 ;
        RECT 415.950 877.800 418.050 879.900 ;
        RECT 421.950 877.800 424.050 879.900 ;
        RECT 425.400 874.050 426.450 946.950 ;
        RECT 431.400 919.050 432.450 961.950 ;
        RECT 443.400 961.350 444.600 962.100 ;
        RECT 449.400 961.350 450.600 962.100 ;
        RECT 473.400 961.350 474.600 963.600 ;
        RECT 478.950 962.100 481.050 964.200 ;
        RECT 484.950 962.100 487.050 964.200 ;
        RECT 479.400 961.350 480.600 962.100 ;
        RECT 442.950 958.950 445.050 961.050 ;
        RECT 445.950 958.950 448.050 961.050 ;
        RECT 448.950 958.950 451.050 961.050 ;
        RECT 451.950 958.950 454.050 961.050 ;
        RECT 469.950 958.950 472.050 961.050 ;
        RECT 472.950 958.950 475.050 961.050 ;
        RECT 475.950 958.950 478.050 961.050 ;
        RECT 478.950 958.950 481.050 961.050 ;
        RECT 446.400 956.400 447.600 958.650 ;
        RECT 452.400 956.400 453.600 958.650 ;
        RECT 470.400 956.400 471.600 958.650 ;
        RECT 476.400 956.400 477.600 958.650 ;
        RECT 485.400 958.050 486.450 962.100 ;
        RECT 446.400 952.050 447.450 956.400 ;
        RECT 445.950 949.950 448.050 952.050 ;
        RECT 448.950 946.950 451.050 949.050 ;
        RECT 430.950 916.950 433.050 919.050 ;
        RECT 439.950 917.100 442.050 919.200 ;
        RECT 440.400 916.350 441.600 917.100 ;
        RECT 436.950 913.950 439.050 916.050 ;
        RECT 439.950 913.950 442.050 916.050 ;
        RECT 437.400 912.900 438.600 913.650 ;
        RECT 436.950 910.800 439.050 912.900 ;
        RECT 449.400 907.050 450.450 946.950 ;
        RECT 439.950 904.950 442.050 907.050 ;
        RECT 448.950 904.950 451.050 907.050 ;
        RECT 433.950 901.950 436.050 904.050 ;
        RECT 434.400 885.600 435.450 901.950 ;
        RECT 440.400 885.600 441.450 904.950 ;
        RECT 452.400 904.050 453.450 956.400 ;
        RECT 470.400 949.050 471.450 956.400 ;
        RECT 476.400 954.450 477.450 956.400 ;
        RECT 484.950 955.950 487.050 958.050 ;
        RECT 476.400 953.400 480.450 954.450 ;
        RECT 472.950 949.950 475.050 952.050 ;
        RECT 469.950 946.950 472.050 949.050 ;
        RECT 466.950 928.950 469.050 931.050 ;
        RECT 460.950 917.100 463.050 922.050 ;
        RECT 467.400 919.200 468.450 928.950 ;
        RECT 466.950 917.100 469.050 919.200 ;
        RECT 461.400 916.350 462.600 917.100 ;
        RECT 467.400 916.350 468.600 917.100 ;
        RECT 457.950 913.950 460.050 916.050 ;
        RECT 460.950 913.950 463.050 916.050 ;
        RECT 463.950 913.950 466.050 916.050 ;
        RECT 466.950 913.950 469.050 916.050 ;
        RECT 458.400 911.400 459.600 913.650 ;
        RECT 464.400 912.900 465.600 913.650 ;
        RECT 451.950 901.950 454.050 904.050 ;
        RECT 434.400 883.350 435.600 885.600 ;
        RECT 440.400 883.350 441.600 885.600 ;
        RECT 442.950 883.950 448.050 886.050 ;
        RECT 430.950 880.950 433.050 883.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 439.950 880.950 442.050 883.050 ;
        RECT 431.400 878.400 432.600 880.650 ;
        RECT 437.400 879.900 438.600 880.650 ;
        RECT 446.400 879.900 447.450 883.950 ;
        RECT 424.950 871.950 427.050 874.050 ;
        RECT 409.950 868.950 412.050 871.050 ;
        RECT 431.400 862.050 432.450 878.400 ;
        RECT 436.950 877.800 439.050 879.900 ;
        RECT 445.950 877.800 448.050 879.900 ;
        RECT 452.400 868.050 453.450 901.950 ;
        RECT 458.400 888.450 459.450 911.400 ;
        RECT 463.950 910.800 466.050 912.900 ;
        RECT 460.950 901.950 463.050 904.050 ;
        RECT 455.400 888.000 459.450 888.450 ;
        RECT 454.950 887.400 459.450 888.000 ;
        RECT 454.950 883.950 457.050 887.400 ;
        RECT 461.400 885.600 462.450 901.950 ;
        RECT 466.950 895.950 469.050 898.050 ;
        RECT 461.400 883.350 462.600 885.600 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 460.950 880.950 463.050 883.050 ;
        RECT 458.400 879.900 459.600 880.650 ;
        RECT 457.950 877.800 460.050 879.900 ;
        RECT 451.950 865.950 454.050 868.050 ;
        RECT 430.950 859.950 433.050 862.050 ;
        RECT 436.950 859.950 439.050 862.050 ;
        RECT 400.950 853.950 403.050 856.050 ;
        RECT 400.950 847.950 403.050 850.050 ;
        RECT 397.950 844.950 400.050 847.050 ;
        RECT 388.950 832.800 391.050 834.900 ;
        RECT 394.950 832.800 397.050 834.900 ;
        RECT 376.950 829.950 379.050 832.050 ;
        RECT 394.950 823.950 397.050 826.050 ;
        RECT 367.950 820.950 370.050 823.050 ;
        RECT 355.950 817.950 358.050 820.050 ;
        RECT 361.950 817.950 364.050 820.050 ;
        RECT 346.950 811.950 349.050 814.050 ;
        RECT 335.400 806.400 339.450 807.450 ;
        RECT 335.400 805.350 336.600 806.400 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 322.950 799.950 325.050 802.050 ;
        RECT 332.400 800.400 333.600 802.650 ;
        RECT 316.950 796.950 319.050 799.050 ;
        RECT 304.950 784.950 307.050 787.050 ;
        RECT 332.400 769.050 333.450 800.400 ;
        RECT 334.950 775.950 337.050 778.050 ;
        RECT 331.950 766.950 334.050 769.050 ;
        RECT 299.400 760.350 300.600 762.600 ;
        RECT 299.100 757.950 301.200 760.050 ;
        RECT 317.100 757.950 319.200 760.050 ;
        RECT 316.950 730.950 319.050 733.050 ;
        RECT 304.950 728.100 307.050 730.200 ;
        RECT 305.400 727.350 306.600 728.100 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 302.400 722.400 303.600 724.650 ;
        RECT 308.400 722.400 309.600 724.650 ;
        RECT 302.400 718.050 303.450 722.400 ;
        RECT 301.950 715.950 304.050 718.050 ;
        RECT 308.400 700.050 309.450 722.400 ;
        RECT 317.400 700.050 318.450 730.950 ;
        RECT 319.950 727.950 322.050 730.050 ;
        RECT 325.950 729.000 328.050 733.050 ;
        RECT 307.950 697.950 310.050 700.050 ;
        RECT 316.950 697.950 319.050 700.050 ;
        RECT 296.400 683.400 300.450 684.450 ;
        RECT 269.400 682.350 270.600 683.100 ;
        RECT 268.800 679.950 270.900 682.050 ;
        RECT 275.400 678.900 276.450 683.100 ;
        RECT 290.400 682.350 291.600 683.100 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 287.400 678.900 288.600 679.650 ;
        RECT 258.900 677.100 267.600 678.300 ;
        RECT 256.800 672.600 258.900 674.700 ;
        RECT 260.100 674.100 262.200 676.200 ;
        RECT 264.000 675.300 266.100 677.100 ;
        RECT 271.800 676.800 273.900 678.900 ;
        RECT 274.950 676.800 277.050 678.900 ;
        RECT 286.950 676.800 289.050 678.900 ;
        RECT 293.400 677.400 294.600 679.650 ;
        RECT 260.400 673.050 261.600 673.800 ;
        RECT 272.400 673.050 273.450 676.800 ;
        RECT 293.400 673.050 294.450 677.400 ;
        RECT 259.950 670.950 262.050 673.050 ;
        RECT 265.950 670.950 268.050 673.050 ;
        RECT 271.950 670.950 274.050 673.050 ;
        RECT 292.950 670.950 295.050 673.050 ;
        RECT 244.950 652.950 247.050 655.050 ;
        RECT 241.950 610.950 244.050 613.050 ;
        RECT 245.400 610.050 246.450 652.950 ;
        RECT 250.950 650.100 253.050 652.200 ;
        RECT 256.950 650.100 259.050 652.200 ;
        RECT 251.400 649.350 252.600 650.100 ;
        RECT 257.400 649.350 258.600 650.100 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 256.950 646.950 259.050 649.050 ;
        RECT 259.950 646.950 262.050 649.050 ;
        RECT 254.400 645.000 255.600 646.650 ;
        RECT 260.400 645.900 261.600 646.650 ;
        RECT 266.400 645.900 267.450 670.950 ;
        RECT 292.950 655.950 295.050 658.050 ;
        RECT 284.400 654.000 291.450 654.450 ;
        RECT 284.400 653.400 292.050 654.000 ;
        RECT 268.950 649.950 271.050 652.050 ;
        RECT 277.950 650.100 280.050 652.200 ;
        RECT 284.400 651.600 285.450 653.400 ;
        RECT 253.950 640.950 256.050 645.000 ;
        RECT 259.950 643.800 262.050 645.900 ;
        RECT 265.950 643.800 268.050 645.900 ;
        RECT 253.950 628.950 256.050 631.050 ;
        RECT 250.950 616.950 253.050 619.050 ;
        RECT 214.950 606.000 217.050 610.050 ;
        RECT 229.950 607.950 232.050 610.050 ;
        RECT 238.950 609.450 243.000 610.050 ;
        RECT 238.950 607.950 243.450 609.450 ;
        RECT 244.950 607.950 247.050 610.050 ;
        RECT 215.400 604.350 216.600 606.000 ;
        RECT 220.950 605.100 223.050 607.200 ;
        RECT 226.950 605.100 229.050 607.200 ;
        RECT 221.400 604.350 222.600 605.100 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 202.950 598.950 205.050 601.050 ;
        RECT 212.400 600.900 213.600 601.650 ;
        RECT 211.950 598.800 214.050 600.900 ;
        RECT 218.400 600.000 219.600 601.650 ;
        RECT 199.950 595.950 202.050 598.050 ;
        RECT 217.950 595.950 220.050 600.000 ;
        RECT 181.950 592.950 184.050 595.050 ;
        RECT 166.950 585.450 169.050 586.050 ;
        RECT 164.400 584.400 169.050 585.450 ;
        RECT 143.400 571.350 144.600 573.000 ;
        RECT 149.400 571.350 150.600 573.000 ;
        RECT 160.950 572.100 163.050 574.200 ;
        RECT 142.950 568.950 145.050 571.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 146.400 567.900 147.600 568.650 ;
        RECT 145.950 565.800 148.050 567.900 ;
        RECT 154.800 565.950 156.900 568.050 ;
        RECT 160.800 565.950 162.900 568.050 ;
        RECT 155.400 564.900 156.600 565.650 ;
        RECT 154.950 562.800 157.050 564.900 ;
        RECT 136.950 556.950 139.050 559.050 ;
        RECT 133.950 538.950 136.050 541.050 ;
        RECT 164.400 538.050 165.450 584.400 ;
        RECT 166.950 583.950 169.050 584.400 ;
        RECT 178.950 583.950 181.050 586.050 ;
        RECT 167.700 579.300 169.800 581.400 ;
        RECT 170.700 579.300 172.800 581.400 ;
        RECT 173.700 579.300 175.800 581.400 ;
        RECT 168.300 575.700 169.500 579.300 ;
        RECT 167.400 573.600 169.500 575.700 ;
        RECT 167.400 554.700 168.900 573.600 ;
        RECT 171.300 562.800 172.500 579.300 ;
        RECT 170.400 560.700 172.500 562.800 ;
        RECT 171.300 554.700 172.500 560.700 ;
        RECT 173.700 557.700 174.900 579.300 ;
        RECT 181.800 578.400 183.900 580.500 ;
        RECT 187.200 579.300 189.300 581.400 ;
        RECT 190.200 579.300 192.300 581.400 ;
        RECT 193.200 579.300 195.300 581.400 ;
        RECT 178.800 571.950 180.900 574.050 ;
        RECT 179.400 570.900 180.600 571.650 ;
        RECT 178.950 568.800 181.050 570.900 ;
        RECT 182.400 567.900 183.300 578.400 ;
        RECT 185.100 572.400 187.200 574.500 ;
        RECT 182.400 565.800 184.500 567.900 ;
        RECT 188.100 567.000 189.300 579.300 ;
        RECT 182.400 559.200 183.300 565.800 ;
        RECT 187.800 564.900 189.900 567.000 ;
        RECT 173.700 555.600 175.800 557.700 ;
        RECT 182.400 557.100 184.500 559.200 ;
        RECT 188.100 557.700 189.300 564.900 ;
        RECT 190.800 561.600 192.300 579.300 ;
        RECT 190.800 559.500 192.900 561.600 ;
        RECT 187.800 555.600 189.900 557.700 ;
        RECT 190.800 554.700 192.300 559.500 ;
        RECT 194.100 557.700 195.300 579.300 ;
        RECT 167.400 552.600 170.400 554.700 ;
        RECT 171.300 552.600 173.400 554.700 ;
        RECT 190.200 552.600 192.300 554.700 ;
        RECT 193.200 552.600 195.300 557.700 ;
        RECT 196.200 579.300 198.300 581.400 ;
        RECT 196.200 561.600 197.700 579.300 ;
        RECT 200.400 571.050 201.450 595.950 ;
        RECT 220.950 592.950 223.050 595.050 ;
        RECT 205.950 586.950 208.050 589.050 ;
        RECT 199.950 568.950 202.050 571.050 ;
        RECT 206.400 570.600 207.450 586.950 ;
        RECT 208.950 571.950 211.050 574.050 ;
        RECT 206.400 568.350 207.600 570.600 ;
        RECT 205.800 565.950 207.900 568.050 ;
        RECT 196.200 559.500 198.300 561.600 ;
        RECT 196.200 554.700 197.700 559.500 ;
        RECT 196.200 552.600 198.300 554.700 ;
        RECT 202.950 550.950 205.050 553.050 ;
        RECT 193.950 541.950 196.050 547.050 ;
        RECT 203.400 544.050 204.450 550.950 ;
        RECT 202.950 541.950 205.050 544.050 ;
        RECT 209.400 541.050 210.450 571.950 ;
        RECT 215.400 570.450 216.600 570.600 ;
        RECT 215.400 569.400 219.450 570.450 ;
        RECT 215.400 568.350 216.600 569.400 ;
        RECT 214.800 565.950 216.900 568.050 ;
        RECT 218.400 559.050 219.450 569.400 ;
        RECT 221.400 562.050 222.450 592.950 ;
        RECT 223.950 580.950 226.050 583.050 ;
        RECT 220.950 559.950 223.050 562.050 ;
        RECT 217.950 556.950 220.050 559.050 ;
        RECT 193.950 538.800 196.050 540.900 ;
        RECT 208.950 538.950 211.050 541.050 ;
        RECT 163.950 535.950 166.050 538.050 ;
        RECT 172.950 535.950 175.050 538.050 ;
        RECT 130.950 532.950 133.050 535.050 ;
        RECT 136.950 532.950 139.050 535.050 ;
        RECT 137.400 528.600 138.450 532.950 ;
        RECT 137.400 526.350 138.600 528.600 ;
        RECT 142.950 527.100 145.050 529.200 ;
        RECT 148.950 527.100 151.050 529.200 ;
        RECT 163.950 527.100 166.050 529.200 ;
        RECT 143.400 526.350 144.600 527.100 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 134.400 522.900 135.600 523.650 ;
        RECT 133.950 520.800 136.050 522.900 ;
        RECT 140.400 521.400 141.600 523.650 ;
        RECT 124.950 514.950 127.050 517.050 ;
        RECT 140.400 514.050 141.450 521.400 ;
        RECT 112.950 511.950 115.050 514.050 ;
        RECT 139.950 511.950 142.050 514.050 ;
        RECT 149.400 511.050 150.450 527.100 ;
        RECT 164.400 526.350 165.600 527.100 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 161.400 521.400 162.600 523.650 ;
        RECT 151.950 517.950 154.050 520.050 ;
        RECT 148.950 508.950 151.050 511.050 ;
        RECT 109.950 494.100 112.050 496.200 ;
        RECT 115.950 494.100 118.050 496.200 ;
        RECT 124.950 494.100 127.050 496.200 ;
        RECT 139.950 494.100 142.050 496.200 ;
        RECT 110.400 493.350 111.600 494.100 ;
        RECT 116.400 493.350 117.600 494.100 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 115.950 490.950 118.050 493.050 ;
        RECT 118.950 490.950 121.050 493.050 ;
        RECT 113.400 489.000 114.600 490.650 ;
        RECT 103.950 484.950 106.050 487.050 ;
        RECT 112.950 484.950 115.050 489.000 ;
        RECT 119.400 488.400 120.600 490.650 ;
        RECT 125.400 490.050 126.450 494.100 ;
        RECT 140.400 493.350 141.600 494.100 ;
        RECT 148.950 493.950 151.050 496.050 ;
        RECT 136.950 490.950 139.050 493.050 ;
        RECT 139.950 490.950 142.050 493.050 ;
        RECT 142.950 490.950 145.050 493.050 ;
        RECT 115.950 484.950 118.050 487.050 ;
        RECT 116.400 460.050 117.450 484.950 ;
        RECT 119.400 483.450 120.450 488.400 ;
        RECT 124.950 487.950 127.050 490.050 ;
        RECT 137.400 489.900 138.600 490.650 ;
        RECT 143.400 489.900 144.600 490.650 ;
        RECT 136.950 487.800 139.050 489.900 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 119.400 483.000 123.450 483.450 ;
        RECT 118.950 482.400 123.450 483.000 ;
        RECT 118.950 478.950 121.050 482.400 ;
        RECT 115.950 457.950 118.050 460.050 ;
        RECT 88.950 449.100 91.050 451.200 ;
        RECT 89.400 448.350 90.600 449.100 ;
        RECT 100.950 448.950 103.050 451.050 ;
        RECT 109.950 449.100 112.050 451.200 ;
        RECT 116.400 450.600 117.450 457.950 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 76.950 442.950 79.050 445.050 ;
        RECT 86.400 444.900 87.600 445.650 ;
        RECT 85.950 442.800 88.050 444.900 ;
        RECT 70.950 436.950 73.050 439.050 ;
        RECT 68.700 423.300 70.800 425.400 ;
        RECT 71.700 423.300 73.800 425.400 ;
        RECT 74.700 423.300 76.800 425.400 ;
        RECT 69.300 419.700 70.500 423.300 ;
        RECT 68.400 417.600 70.500 419.700 ;
        RECT 55.950 403.950 58.050 408.000 ;
        RECT 58.950 406.950 61.050 409.050 ;
        RECT 64.950 406.950 67.050 409.050 ;
        RECT 43.950 391.950 46.050 394.050 ;
        RECT 44.400 376.050 45.450 391.950 ;
        RECT 46.950 376.950 49.050 379.050 ;
        RECT 43.950 373.950 46.050 376.050 ;
        RECT 47.400 372.600 48.450 376.950 ;
        RECT 52.950 373.950 55.050 376.050 ;
        RECT 41.400 370.350 42.600 372.600 ;
        RECT 47.400 370.350 48.600 372.600 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 38.400 365.400 39.600 367.650 ;
        RECT 44.400 366.900 45.600 367.650 ;
        RECT 53.400 366.900 54.450 373.950 ;
        RECT 38.400 352.050 39.450 365.400 ;
        RECT 43.950 364.800 46.050 366.900 ;
        RECT 52.950 364.800 55.050 366.900 ;
        RECT 7.950 349.950 10.050 352.050 ;
        RECT 28.950 349.950 31.050 352.050 ;
        RECT 37.950 349.950 40.050 352.050 ;
        RECT 8.400 337.050 9.450 349.950 ;
        RECT 17.700 345.300 19.800 347.400 ;
        RECT 20.700 345.300 22.800 347.400 ;
        RECT 23.700 345.300 25.800 347.400 ;
        RECT 18.300 341.700 19.500 345.300 ;
        RECT 17.400 339.600 19.500 341.700 ;
        RECT 7.950 334.950 10.050 337.050 ;
        RECT 4.800 331.950 6.900 334.050 ;
        RECT 10.800 331.950 12.900 334.050 ;
        RECT 5.400 330.900 6.600 331.650 ;
        RECT 4.950 328.800 7.050 330.900 ;
        RECT 17.400 320.700 18.900 339.600 ;
        RECT 21.300 328.800 22.500 345.300 ;
        RECT 20.400 326.700 22.500 328.800 ;
        RECT 21.300 320.700 22.500 326.700 ;
        RECT 23.700 323.700 24.900 345.300 ;
        RECT 31.800 344.400 33.900 346.500 ;
        RECT 37.200 345.300 39.300 347.400 ;
        RECT 40.200 345.300 42.300 347.400 ;
        RECT 43.200 345.300 45.300 347.400 ;
        RECT 28.800 337.950 30.900 340.050 ;
        RECT 29.400 336.000 30.600 337.650 ;
        RECT 28.950 331.950 31.050 336.000 ;
        RECT 32.400 333.900 33.300 344.400 ;
        RECT 35.100 338.400 37.200 340.500 ;
        RECT 32.400 331.800 34.500 333.900 ;
        RECT 38.100 333.000 39.300 345.300 ;
        RECT 32.400 325.200 33.300 331.800 ;
        RECT 37.800 330.900 39.900 333.000 ;
        RECT 23.700 321.600 25.800 323.700 ;
        RECT 32.400 323.100 34.500 325.200 ;
        RECT 38.100 323.700 39.300 330.900 ;
        RECT 40.800 327.600 42.300 345.300 ;
        RECT 40.800 325.500 42.900 327.600 ;
        RECT 37.800 321.600 39.900 323.700 ;
        RECT 40.800 320.700 42.300 325.500 ;
        RECT 44.100 323.700 45.300 345.300 ;
        RECT 17.400 318.600 20.400 320.700 ;
        RECT 21.300 318.600 23.400 320.700 ;
        RECT 40.200 318.600 42.300 320.700 ;
        RECT 43.200 318.600 45.300 323.700 ;
        RECT 46.200 345.300 48.300 347.400 ;
        RECT 46.200 327.600 47.700 345.300 ;
        RECT 55.950 340.950 58.050 343.050 ;
        RECT 56.400 336.600 57.450 340.950 ;
        RECT 56.400 334.350 57.600 336.600 ;
        RECT 55.800 331.950 57.900 334.050 ;
        RECT 46.200 325.500 48.300 327.600 ;
        RECT 46.200 320.700 47.700 325.500 ;
        RECT 46.200 318.600 48.300 320.700 ;
        RECT 16.950 293.100 19.050 295.200 ;
        RECT 22.950 293.100 25.050 295.200 ;
        RECT 37.950 293.100 40.050 295.200 ;
        RECT 43.950 293.100 46.050 295.200 ;
        RECT 49.950 293.100 52.050 295.200 ;
        RECT 17.400 292.350 18.600 293.100 ;
        RECT 23.400 292.350 24.600 293.100 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 22.950 289.950 25.050 292.050 ;
        RECT 25.950 289.950 28.050 292.050 ;
        RECT 13.950 286.950 16.050 289.050 ;
        RECT 20.400 288.000 21.600 289.650 ;
        RECT 26.400 288.900 27.600 289.650 ;
        RECT 38.400 289.050 39.450 293.100 ;
        RECT 44.400 292.350 45.600 293.100 ;
        RECT 50.400 292.350 51.600 293.100 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 49.950 289.950 52.050 292.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 10.950 283.950 13.050 286.050 ;
        RECT 11.400 211.050 12.450 283.950 ;
        RECT 14.400 268.050 15.450 286.950 ;
        RECT 19.950 283.950 22.050 288.000 ;
        RECT 25.950 286.800 28.050 288.900 ;
        RECT 37.950 286.950 40.050 289.050 ;
        RECT 47.400 287.400 48.600 289.650 ;
        RECT 53.400 288.900 54.600 289.650 ;
        RECT 59.400 289.050 60.450 406.950 ;
        RECT 68.400 398.700 69.900 417.600 ;
        RECT 72.300 406.800 73.500 423.300 ;
        RECT 71.400 404.700 73.500 406.800 ;
        RECT 72.300 398.700 73.500 404.700 ;
        RECT 74.700 401.700 75.900 423.300 ;
        RECT 82.800 422.400 84.900 424.500 ;
        RECT 88.200 423.300 90.300 425.400 ;
        RECT 91.200 423.300 93.300 425.400 ;
        RECT 94.200 423.300 96.300 425.400 ;
        RECT 79.800 415.950 81.900 418.050 ;
        RECT 80.400 414.900 81.600 415.650 ;
        RECT 79.950 412.800 82.050 414.900 ;
        RECT 83.400 411.900 84.300 422.400 ;
        RECT 86.100 416.400 88.200 418.500 ;
        RECT 83.400 409.800 85.500 411.900 ;
        RECT 89.100 411.000 90.300 423.300 ;
        RECT 83.400 403.200 84.300 409.800 ;
        RECT 88.800 408.900 90.900 411.000 ;
        RECT 74.700 399.600 76.800 401.700 ;
        RECT 83.400 401.100 85.500 403.200 ;
        RECT 89.100 401.700 90.300 408.900 ;
        RECT 91.800 405.600 93.300 423.300 ;
        RECT 91.800 403.500 93.900 405.600 ;
        RECT 88.800 399.600 90.900 401.700 ;
        RECT 91.800 398.700 93.300 403.500 ;
        RECT 95.100 401.700 96.300 423.300 ;
        RECT 68.400 396.600 71.400 398.700 ;
        RECT 72.300 396.600 74.400 398.700 ;
        RECT 91.200 396.600 93.300 398.700 ;
        RECT 94.200 396.600 96.300 401.700 ;
        RECT 97.200 423.300 99.300 425.400 ;
        RECT 101.400 423.450 102.450 448.950 ;
        RECT 110.400 448.350 111.600 449.100 ;
        RECT 116.400 448.350 117.600 450.600 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 107.400 444.900 108.600 445.650 ;
        RECT 106.950 442.800 109.050 444.900 ;
        RECT 113.400 443.400 114.600 445.650 ;
        RECT 106.950 436.950 109.050 439.050 ;
        RECT 97.200 405.600 98.700 423.300 ;
        RECT 101.400 422.400 105.450 423.450 ;
        RECT 104.400 414.900 105.450 422.400 ;
        RECT 103.950 412.800 106.050 414.900 ;
        RECT 107.400 414.600 108.450 436.950 ;
        RECT 113.400 436.050 114.450 443.400 ;
        RECT 118.950 442.800 121.050 444.900 ;
        RECT 112.950 433.950 115.050 436.050 ;
        RECT 107.400 414.450 108.600 414.600 ;
        RECT 107.400 413.400 111.450 414.450 ;
        RECT 115.950 414.000 118.050 418.050 ;
        RECT 107.400 412.350 108.600 413.400 ;
        RECT 106.800 409.950 108.900 412.050 ;
        RECT 97.200 403.500 99.300 405.600 ;
        RECT 97.200 398.700 98.700 403.500 ;
        RECT 97.200 396.600 99.300 398.700 ;
        RECT 67.950 388.950 70.050 391.050 ;
        RECT 110.400 390.450 111.450 413.400 ;
        RECT 116.400 412.350 117.600 414.000 ;
        RECT 115.800 409.950 117.900 412.050 ;
        RECT 107.400 389.400 111.450 390.450 ;
        RECT 68.400 372.600 69.450 388.950 ;
        RECT 103.950 385.950 106.050 388.050 ;
        RECT 93.000 375.450 97.050 376.050 ;
        RECT 92.400 373.950 97.050 375.450 ;
        RECT 68.400 370.350 69.600 372.600 ;
        RECT 79.950 370.950 82.050 373.050 ;
        RECT 92.400 372.600 93.450 373.950 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 67.950 367.950 70.050 370.050 ;
        RECT 70.950 367.950 73.050 370.050 ;
        RECT 65.400 365.400 66.600 367.650 ;
        RECT 71.400 365.400 72.600 367.650 ;
        RECT 65.400 361.050 66.450 365.400 ;
        RECT 64.950 358.950 67.050 361.050 ;
        RECT 65.400 336.600 66.450 358.950 ;
        RECT 71.400 352.050 72.450 365.400 ;
        RECT 73.950 364.950 76.050 367.050 ;
        RECT 70.950 349.950 73.050 352.050 ;
        RECT 65.400 334.350 66.600 336.600 ;
        RECT 64.800 331.950 66.900 334.050 ;
        RECT 71.400 319.050 72.450 349.950 ;
        RECT 70.950 316.950 73.050 319.050 ;
        RECT 61.950 313.950 64.050 316.050 ;
        RECT 22.950 283.950 25.050 286.050 ;
        RECT 13.950 265.950 16.050 268.050 ;
        RECT 23.400 267.450 24.450 283.950 ;
        RECT 38.400 280.050 39.450 286.950 ;
        RECT 43.950 283.950 46.050 286.050 ;
        RECT 37.950 277.950 40.050 280.050 ;
        RECT 19.800 264.300 21.900 266.400 ;
        RECT 23.400 265.200 24.600 267.450 ;
        RECT 16.950 260.100 19.050 262.200 ;
        RECT 17.400 259.350 18.600 260.100 ;
        RECT 17.100 256.950 19.200 259.050 ;
        RECT 20.100 258.900 21.000 264.300 ;
        RECT 23.100 262.800 25.200 264.900 ;
        RECT 27.000 261.900 29.100 263.700 ;
        RECT 21.900 260.700 30.600 261.900 ;
        RECT 21.900 259.800 24.000 260.700 ;
        RECT 20.100 257.700 27.000 258.900 ;
        RECT 20.100 250.500 21.300 257.700 ;
        RECT 23.100 253.950 25.200 256.050 ;
        RECT 26.100 255.300 27.000 257.700 ;
        RECT 23.400 251.400 24.600 253.650 ;
        RECT 26.100 253.200 28.200 255.300 ;
        RECT 29.700 251.700 30.600 260.700 ;
        RECT 31.800 256.950 33.900 259.050 ;
        RECT 32.400 255.900 33.600 256.650 ;
        RECT 31.950 253.800 34.050 255.900 ;
        RECT 40.950 253.800 43.050 255.900 ;
        RECT 19.800 248.400 21.900 250.500 ;
        RECT 29.400 249.600 31.500 251.700 ;
        RECT 41.400 241.050 42.450 253.800 ;
        RECT 44.400 247.050 45.450 283.950 ;
        RECT 47.400 271.050 48.450 287.400 ;
        RECT 52.950 286.800 55.050 288.900 ;
        RECT 58.950 286.950 61.050 289.050 ;
        RECT 46.950 268.950 49.050 271.050 ;
        RECT 58.950 268.950 61.050 271.050 ;
        RECT 52.950 260.100 55.050 262.200 ;
        RECT 53.400 259.350 54.600 260.100 ;
        RECT 49.950 256.950 52.050 259.050 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 50.400 254.400 51.600 256.650 ;
        RECT 43.950 244.950 46.050 247.050 ;
        RECT 40.950 238.950 43.050 241.050 ;
        RECT 28.950 232.950 31.050 235.050 ;
        RECT 22.950 226.950 25.050 229.050 ;
        RECT 16.950 215.100 19.050 217.200 ;
        RECT 23.400 216.600 24.450 226.950 ;
        RECT 17.400 214.350 18.600 215.100 ;
        RECT 23.400 214.350 24.600 216.600 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 19.950 211.950 22.050 214.050 ;
        RECT 22.950 211.950 25.050 214.050 ;
        RECT 10.950 208.950 13.050 211.050 ;
        RECT 20.400 210.900 21.600 211.650 ;
        RECT 19.950 208.800 22.050 210.900 ;
        RECT 19.950 190.950 22.050 193.050 ;
        RECT 20.400 183.600 21.450 190.950 ;
        RECT 20.400 181.350 21.600 183.600 ;
        RECT 25.950 181.950 28.050 184.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 17.400 177.000 18.600 178.650 ;
        RECT 16.950 172.950 19.050 177.000 ;
        RECT 26.400 142.050 27.450 181.950 ;
        RECT 29.400 175.050 30.450 232.950 ;
        RECT 34.950 220.950 37.050 223.050 ;
        RECT 31.950 215.100 34.050 217.200 ;
        RECT 32.400 193.050 33.450 215.100 ;
        RECT 31.950 190.950 34.050 193.050 ;
        RECT 28.950 172.950 31.050 175.050 ;
        RECT 29.400 145.050 30.450 172.950 ;
        RECT 28.950 142.950 31.050 145.050 ;
        RECT 25.950 139.950 28.050 142.050 ;
        RECT 19.950 137.100 22.050 139.200 ;
        RECT 26.400 138.600 27.450 139.950 ;
        RECT 32.400 139.200 33.450 190.950 ;
        RECT 35.400 184.050 36.450 220.950 ;
        RECT 41.400 216.600 42.450 238.950 ;
        RECT 50.400 223.050 51.450 254.400 ;
        RECT 52.950 244.950 55.050 247.050 ;
        RECT 49.950 220.950 52.050 223.050 ;
        RECT 41.400 214.350 42.600 216.600 ;
        RECT 47.400 216.450 48.600 216.600 ;
        RECT 50.400 216.450 51.450 220.950 ;
        RECT 47.400 215.400 51.450 216.450 ;
        RECT 47.400 214.350 48.600 215.400 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 46.950 211.950 49.050 214.050 ;
        RECT 44.400 209.400 45.600 211.650 ;
        RECT 44.400 190.050 45.450 209.400 ;
        RECT 53.400 208.050 54.450 244.950 ;
        RECT 59.400 211.050 60.450 268.950 ;
        RECT 62.400 262.200 63.450 313.950 ;
        RECT 74.400 307.050 75.450 364.950 ;
        RECT 80.400 361.050 81.450 370.950 ;
        RECT 92.400 370.350 93.600 372.600 ;
        RECT 88.950 367.950 91.050 370.050 ;
        RECT 91.950 367.950 94.050 370.050 ;
        RECT 94.950 367.950 97.050 370.050 ;
        RECT 89.400 366.900 90.600 367.650 ;
        RECT 88.950 364.800 91.050 366.900 ;
        RECT 95.400 365.400 96.600 367.650 ;
        RECT 104.400 367.050 105.450 385.950 ;
        RECT 79.950 360.450 82.050 361.050 ;
        RECT 79.950 359.400 84.450 360.450 ;
        RECT 79.950 358.950 82.050 359.400 ;
        RECT 64.950 304.950 67.050 307.050 ;
        RECT 73.950 304.950 76.050 307.050 ;
        RECT 61.950 260.100 64.050 262.200 ;
        RECT 65.400 255.900 66.450 304.950 ;
        RECT 76.950 298.950 79.050 301.050 ;
        RECT 70.950 293.100 73.050 295.200 ;
        RECT 77.400 294.600 78.450 298.950 ;
        RECT 71.400 292.350 72.600 293.100 ;
        RECT 77.400 292.350 78.600 294.600 ;
        RECT 70.950 289.950 73.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 74.400 288.900 75.600 289.650 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 73.950 265.950 76.050 268.050 ;
        RECT 74.400 261.600 75.450 265.950 ;
        RECT 74.400 259.350 75.600 261.600 ;
        RECT 70.950 256.950 73.050 259.050 ;
        RECT 73.950 256.950 76.050 259.050 ;
        RECT 76.950 256.950 79.050 259.050 ;
        RECT 71.400 255.900 72.600 256.650 ;
        RECT 64.950 253.800 67.050 255.900 ;
        RECT 70.950 253.800 73.050 255.900 ;
        RECT 77.400 254.400 78.600 256.650 ;
        RECT 65.400 235.050 66.450 253.800 ;
        RECT 64.950 232.950 67.050 235.050 ;
        RECT 77.400 232.050 78.450 254.400 ;
        RECT 76.950 229.950 79.050 232.050 ;
        RECT 64.950 226.950 67.050 229.050 ;
        RECT 65.400 216.600 66.450 226.950 ;
        RECT 77.400 226.050 78.450 229.950 ;
        RECT 70.950 223.950 73.050 226.050 ;
        RECT 76.950 223.950 79.050 226.050 ;
        RECT 65.400 214.350 66.600 216.600 ;
        RECT 71.400 216.450 72.450 223.950 ;
        RECT 76.950 217.950 79.050 220.050 ;
        RECT 71.400 215.400 75.450 216.450 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 58.950 208.950 61.050 211.050 ;
        RECT 68.400 209.400 69.600 211.650 ;
        RECT 46.950 205.950 49.050 208.050 ;
        RECT 52.950 205.950 55.050 208.050 ;
        RECT 37.950 187.950 40.050 190.050 ;
        RECT 43.950 187.950 46.050 190.050 ;
        RECT 34.950 181.950 37.050 184.050 ;
        RECT 38.400 183.600 39.450 187.950 ;
        RECT 47.400 186.450 48.450 205.950 ;
        RECT 68.400 196.050 69.450 209.400 ;
        RECT 74.400 196.050 75.450 215.400 ;
        RECT 67.950 193.950 70.050 196.050 ;
        RECT 73.950 193.950 76.050 196.050 ;
        RECT 58.950 190.950 61.050 193.050 ;
        RECT 44.400 185.400 48.450 186.450 ;
        RECT 44.400 183.600 45.450 185.400 ;
        RECT 38.400 181.350 39.600 183.600 ;
        RECT 44.400 181.350 45.600 183.600 ;
        RECT 52.950 181.950 55.050 184.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 41.400 176.400 42.600 178.650 ;
        RECT 47.400 177.900 48.600 178.650 ;
        RECT 53.400 177.900 54.450 181.950 ;
        RECT 59.400 177.900 60.450 190.950 ;
        RECT 67.950 182.100 70.050 184.200 ;
        RECT 68.400 181.350 69.600 182.100 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 70.950 178.950 73.050 181.050 ;
        RECT 65.400 177.900 66.600 178.650 ;
        RECT 71.400 177.900 72.600 178.650 ;
        RECT 41.400 172.050 42.450 176.400 ;
        RECT 46.950 175.800 49.050 177.900 ;
        RECT 52.950 175.800 55.050 177.900 ;
        RECT 58.950 175.800 61.050 177.900 ;
        RECT 64.950 175.800 67.050 177.900 ;
        RECT 70.950 175.800 73.050 177.900 ;
        RECT 40.950 169.950 43.050 172.050 ;
        RECT 77.400 157.050 78.450 217.950 ;
        RECT 83.400 216.450 84.450 359.400 ;
        RECT 88.800 334.950 90.900 337.050 ;
        RECT 95.400 328.050 96.450 365.400 ;
        RECT 103.950 364.950 106.050 367.050 ;
        RECT 107.400 342.450 108.450 389.400 ;
        RECT 119.400 382.050 120.450 442.800 ;
        RECT 122.400 427.050 123.450 482.400 ;
        RECT 137.400 450.600 138.450 487.800 ;
        RECT 142.950 484.950 145.050 489.900 ;
        RECT 149.400 469.050 150.450 493.950 ;
        RECT 148.950 466.950 151.050 469.050 ;
        RECT 137.400 448.350 138.600 450.600 ;
        RECT 145.950 449.100 148.050 451.200 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 134.400 444.900 135.600 445.650 ;
        RECT 133.950 439.950 136.050 444.900 ;
        RECT 140.400 443.400 141.600 445.650 ;
        RECT 121.950 424.950 124.050 427.050 ;
        RECT 130.950 424.950 133.050 427.050 ;
        RECT 127.950 416.100 130.050 418.200 ;
        RECT 128.400 397.050 129.450 416.100 ;
        RECT 127.950 394.950 130.050 397.050 ;
        RECT 118.950 379.950 121.050 382.050 ;
        RECT 112.950 371.100 115.050 373.200 ;
        RECT 118.950 372.000 121.050 376.050 ;
        RECT 113.400 370.350 114.600 371.100 ;
        RECT 119.400 370.350 120.600 372.000 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 116.400 366.000 117.600 367.650 ;
        RECT 122.400 366.900 123.600 367.650 ;
        RECT 115.950 363.450 118.050 366.000 ;
        RECT 121.950 364.800 124.050 366.900 ;
        RECT 113.400 362.400 118.050 363.450 ;
        RECT 109.950 342.450 112.050 343.050 ;
        RECT 107.400 341.400 112.050 342.450 ;
        RECT 109.950 340.950 112.050 341.400 ;
        RECT 106.800 334.950 108.900 337.050 ;
        RECT 107.400 333.450 108.600 334.650 ;
        RECT 110.400 333.450 111.450 340.950 ;
        RECT 107.400 332.400 111.450 333.450 ;
        RECT 94.950 325.950 97.050 328.050 ;
        RECT 106.950 322.950 109.050 325.050 ;
        RECT 85.950 316.950 88.050 319.050 ;
        RECT 86.400 220.200 87.450 316.950 ;
        RECT 100.950 298.950 103.050 301.050 ;
        RECT 88.950 293.100 91.050 295.200 ;
        RECT 94.950 293.100 97.050 295.200 ;
        RECT 101.400 294.600 102.450 298.950 ;
        RECT 107.400 294.600 108.450 322.950 ;
        RECT 113.400 316.050 114.450 362.400 ;
        RECT 115.950 361.950 118.050 362.400 ;
        RECT 115.950 352.950 118.050 355.050 ;
        RECT 112.950 313.950 115.050 316.050 ;
        RECT 89.400 280.050 90.450 293.100 ;
        RECT 95.400 292.350 96.600 293.100 ;
        RECT 101.400 292.350 102.600 294.600 ;
        RECT 107.400 292.350 108.600 294.600 ;
        RECT 112.950 293.100 115.050 295.200 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 98.400 287.400 99.600 289.650 ;
        RECT 104.400 288.900 105.600 289.650 ;
        RECT 98.400 280.050 99.450 287.400 ;
        RECT 103.950 286.800 106.050 288.900 ;
        RECT 103.950 280.950 106.050 283.050 ;
        RECT 88.950 277.950 91.050 280.050 ;
        RECT 97.950 277.950 100.050 280.050 ;
        RECT 97.950 260.100 100.050 262.200 ;
        RECT 104.400 261.600 105.450 280.950 ;
        RECT 98.400 259.350 99.600 260.100 ;
        RECT 104.400 259.350 105.600 261.600 ;
        RECT 109.950 260.100 112.050 262.200 ;
        RECT 94.950 256.950 97.050 259.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 95.400 254.400 96.600 256.650 ;
        RECT 101.400 254.400 102.600 256.650 ;
        RECT 95.400 229.050 96.450 254.400 ;
        RECT 101.400 244.050 102.450 254.400 ;
        RECT 106.950 253.950 109.050 256.050 ;
        RECT 100.950 241.950 103.050 244.050 ;
        RECT 94.950 226.950 97.050 229.050 ;
        RECT 91.950 220.950 94.050 223.050 ;
        RECT 85.950 218.100 88.050 220.200 ;
        RECT 80.400 215.400 84.450 216.450 ;
        RECT 80.400 187.050 81.450 215.400 ;
        RECT 85.950 214.950 88.050 217.050 ;
        RECT 92.400 216.600 93.450 220.950 ;
        RECT 86.400 214.350 87.600 214.950 ;
        RECT 92.400 214.350 93.600 216.600 ;
        RECT 103.950 215.100 106.050 217.200 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 89.400 210.900 90.600 211.650 ;
        RECT 88.950 208.800 91.050 210.900 ;
        RECT 95.400 209.400 96.600 211.650 ;
        RECT 82.950 193.950 85.050 196.050 ;
        RECT 79.950 184.950 82.050 187.050 ;
        RECT 76.950 154.950 79.050 157.050 ;
        RECT 76.950 142.950 79.050 145.050 ;
        RECT 20.400 136.350 21.600 137.100 ;
        RECT 26.400 136.350 27.600 138.600 ;
        RECT 31.950 138.450 34.050 139.200 ;
        RECT 31.950 137.400 36.450 138.450 ;
        RECT 31.950 137.100 34.050 137.400 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 28.950 133.950 31.050 136.050 ;
        RECT 17.400 131.400 18.600 133.650 ;
        RECT 23.400 131.400 24.600 133.650 ;
        RECT 29.400 132.900 30.600 133.650 ;
        RECT 13.950 112.950 16.050 115.050 ;
        RECT 14.400 105.450 15.450 112.950 ;
        RECT 17.400 109.050 18.450 131.400 ;
        RECT 23.400 121.050 24.450 131.400 ;
        RECT 28.950 130.800 31.050 132.900 ;
        RECT 22.950 118.950 25.050 121.050 ;
        RECT 16.950 106.950 19.050 109.050 ;
        RECT 17.400 105.450 18.600 105.600 ;
        RECT 14.400 104.400 18.600 105.450 ;
        RECT 17.400 103.350 18.600 104.400 ;
        RECT 22.950 104.100 25.050 109.050 ;
        RECT 23.400 103.350 24.600 104.100 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 20.400 99.900 21.600 100.650 ;
        RECT 19.950 97.800 22.050 99.900 ;
        RECT 29.400 94.050 30.450 130.800 ;
        RECT 35.400 115.050 36.450 137.400 ;
        RECT 40.950 137.100 43.050 139.200 ;
        RECT 46.950 138.000 49.050 142.050 ;
        RECT 41.400 133.050 42.450 137.100 ;
        RECT 47.400 136.350 48.600 138.000 ;
        RECT 52.950 137.100 55.050 139.200 ;
        RECT 64.950 137.100 67.050 139.200 ;
        RECT 70.950 137.100 73.050 139.200 ;
        RECT 77.400 138.600 78.450 142.950 ;
        RECT 80.400 142.050 81.450 184.950 ;
        RECT 83.400 178.050 84.450 193.950 ;
        RECT 95.400 193.050 96.450 209.400 ;
        RECT 104.400 199.050 105.450 215.100 ;
        RECT 103.950 196.950 106.050 199.050 ;
        RECT 88.950 190.950 91.050 193.050 ;
        RECT 94.950 190.950 97.050 193.050 ;
        RECT 89.400 183.600 90.450 190.950 ;
        RECT 89.400 181.350 90.600 183.600 ;
        RECT 94.950 182.100 97.050 184.200 ;
        RECT 100.950 182.100 103.050 184.200 ;
        RECT 95.400 181.350 96.600 182.100 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 82.950 175.950 85.050 178.050 ;
        RECT 92.400 176.400 93.600 178.650 ;
        RECT 101.400 177.900 102.450 182.100 ;
        RECT 92.400 172.050 93.450 176.400 ;
        RECT 100.950 175.800 103.050 177.900 ;
        RECT 91.950 169.950 94.050 172.050 ;
        RECT 91.950 166.800 94.050 168.900 ;
        RECT 79.950 139.950 82.050 142.050 ;
        RECT 85.950 139.950 88.050 142.050 ;
        RECT 53.400 136.350 54.600 137.100 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 40.950 130.950 43.050 133.050 ;
        RECT 50.400 132.900 51.600 133.650 ;
        RECT 65.400 133.050 66.450 137.100 ;
        RECT 71.400 136.350 72.600 137.100 ;
        RECT 77.400 136.350 78.600 138.600 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 49.950 130.800 52.050 132.900 ;
        RECT 64.950 130.950 67.050 133.050 ;
        RECT 74.400 131.400 75.600 133.650 ;
        RECT 80.400 131.400 81.600 133.650 ;
        RECT 34.950 112.950 37.050 115.050 ;
        RECT 31.950 104.100 34.050 106.200 ;
        RECT 28.950 91.950 31.050 94.050 ;
        RECT 16.950 79.950 19.050 82.050 ;
        RECT 17.400 60.600 18.450 79.950 ;
        RECT 32.400 73.050 33.450 104.100 ;
        RECT 35.400 82.050 36.450 112.950 ;
        RECT 43.950 104.100 46.050 106.200 ;
        RECT 50.400 105.600 51.450 130.800 ;
        RECT 67.950 118.950 70.050 121.050 ;
        RECT 68.400 105.600 69.450 118.950 ;
        RECT 74.400 105.600 75.450 131.400 ;
        RECT 80.400 121.050 81.450 131.400 ;
        RECT 79.950 118.950 82.050 121.050 ;
        RECT 44.400 103.350 45.600 104.100 ;
        RECT 50.400 103.350 51.600 105.600 ;
        RECT 68.400 103.350 69.600 105.600 ;
        RECT 74.400 103.350 75.600 105.600 ;
        RECT 82.950 103.950 85.050 106.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 41.400 98.400 42.600 100.650 ;
        RECT 47.400 99.900 48.600 100.650 ;
        RECT 71.400 99.900 72.600 100.650 ;
        RECT 41.400 93.450 42.450 98.400 ;
        RECT 46.950 97.800 49.050 99.900 ;
        RECT 70.950 97.800 73.050 99.900 ;
        RECT 83.400 97.050 84.450 103.950 ;
        RECT 82.950 94.950 85.050 97.050 ;
        RECT 38.400 92.400 42.450 93.450 ;
        RECT 34.950 79.950 37.050 82.050 ;
        RECT 22.950 70.950 25.050 73.050 ;
        RECT 31.950 70.950 34.050 73.050 ;
        RECT 23.400 60.600 24.450 70.950 ;
        RECT 17.400 58.350 18.600 60.600 ;
        RECT 23.400 58.350 24.600 60.600 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 20.400 54.900 21.600 55.650 ;
        RECT 38.400 55.050 39.450 92.400 ;
        RECT 40.950 73.950 43.050 76.050 ;
        RECT 67.950 73.950 70.050 76.050 ;
        RECT 41.400 60.600 42.450 73.950 ;
        RECT 68.400 60.600 69.450 73.950 ;
        RECT 82.950 61.950 85.050 64.050 ;
        RECT 41.400 58.350 42.600 60.600 ;
        RECT 50.400 60.450 51.600 60.600 ;
        RECT 50.400 59.400 54.450 60.450 ;
        RECT 50.400 58.350 51.600 59.400 ;
        RECT 41.100 55.950 43.200 58.050 ;
        RECT 44.400 55.950 46.500 58.050 ;
        RECT 49.800 55.950 51.900 58.050 ;
        RECT 19.950 52.800 22.050 54.900 ;
        RECT 37.950 52.950 40.050 55.050 ;
        RECT 44.400 54.000 45.600 55.650 ;
        RECT 43.950 49.950 46.050 54.000 ;
        RECT 22.950 31.950 25.050 34.050 ;
        RECT 46.950 31.950 49.050 34.050 ;
        RECT 23.400 27.600 24.450 31.950 ;
        RECT 47.400 27.600 48.450 31.950 ;
        RECT 23.400 25.350 24.600 27.600 ;
        RECT 47.400 25.350 48.600 27.600 ;
        RECT 17.100 22.950 19.200 25.050 ;
        RECT 22.500 22.950 24.600 25.050 ;
        RECT 41.100 22.950 43.200 25.050 ;
        RECT 46.500 22.950 48.600 25.050 ;
        RECT 53.400 21.900 54.450 59.400 ;
        RECT 68.400 58.350 69.600 60.600 ;
        RECT 73.950 59.100 76.050 61.200 ;
        RECT 74.400 58.350 75.600 59.100 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 70.950 55.950 73.050 58.050 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 71.400 54.000 72.600 55.650 ;
        RECT 77.400 54.900 78.600 55.650 ;
        RECT 83.400 55.050 84.450 61.950 ;
        RECT 70.950 49.950 73.050 54.000 ;
        RECT 76.950 52.800 79.050 54.900 ;
        RECT 82.950 52.950 85.050 55.050 ;
        RECT 86.400 52.050 87.450 139.950 ;
        RECT 92.400 127.050 93.450 166.800 ;
        RECT 101.400 148.050 102.450 175.800 ;
        RECT 107.400 169.050 108.450 253.950 ;
        RECT 110.400 241.050 111.450 260.100 ;
        RECT 113.400 256.050 114.450 293.100 ;
        RECT 116.400 283.050 117.450 352.950 ;
        RECT 128.400 352.050 129.450 394.950 ;
        RECT 131.400 364.050 132.450 424.950 ;
        RECT 140.400 424.050 141.450 443.400 ;
        RECT 146.400 424.050 147.450 449.100 ;
        RECT 149.400 436.050 150.450 466.950 ;
        RECT 152.400 444.450 153.450 517.950 ;
        RECT 161.400 517.050 162.450 521.400 ;
        RECT 160.950 514.950 163.050 517.050 ;
        RECT 161.400 498.450 162.450 514.950 ;
        RECT 173.400 499.050 174.450 535.950 ;
        RECT 175.950 526.950 178.050 529.050 ;
        RECT 178.950 528.600 183.000 529.050 ;
        RECT 178.950 526.950 183.600 528.600 ;
        RECT 187.950 527.100 190.050 529.200 ;
        RECT 176.400 499.050 177.450 526.950 ;
        RECT 182.400 526.350 183.600 526.950 ;
        RECT 188.400 526.350 189.600 527.100 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 178.950 520.950 181.050 523.050 ;
        RECT 185.400 521.400 186.600 523.650 ;
        RECT 179.400 502.050 180.450 520.950 ;
        RECT 185.400 511.050 186.450 521.400 ;
        RECT 184.950 508.950 187.050 511.050 ;
        RECT 194.400 502.050 195.450 538.800 ;
        RECT 208.950 535.800 211.050 537.900 ;
        RECT 199.950 527.100 202.050 529.200 ;
        RECT 209.400 528.600 210.450 535.800 ;
        RECT 200.400 520.050 201.450 527.100 ;
        RECT 209.400 526.350 210.600 528.600 ;
        RECT 214.950 527.100 217.050 529.200 ;
        RECT 218.400 529.050 219.450 556.950 ;
        RECT 220.950 553.950 223.050 556.050 ;
        RECT 215.400 526.350 216.600 527.100 ;
        RECT 217.950 526.950 220.050 529.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 211.950 523.950 214.050 526.050 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 206.400 522.900 207.600 523.650 ;
        RECT 205.950 520.800 208.050 522.900 ;
        RECT 212.400 521.400 213.600 523.650 ;
        RECT 199.950 517.950 202.050 520.050 ;
        RECT 196.950 502.950 199.050 505.050 ;
        RECT 202.950 502.950 205.050 505.050 ;
        RECT 178.950 499.950 181.050 502.050 ;
        RECT 187.950 499.950 190.050 502.050 ;
        RECT 193.950 499.950 196.050 502.050 ;
        RECT 158.400 497.400 162.450 498.450 ;
        RECT 158.400 481.050 159.450 497.400 ;
        RECT 166.950 495.000 169.050 499.050 ;
        RECT 172.950 496.950 175.050 499.050 ;
        RECT 175.950 496.950 178.050 499.050 ;
        RECT 177.000 495.600 181.050 496.050 ;
        RECT 167.400 493.350 168.600 495.000 ;
        RECT 176.400 493.950 181.050 495.600 ;
        RECT 184.950 493.950 187.050 496.050 ;
        RECT 176.400 493.350 177.600 493.950 ;
        RECT 161.400 490.950 163.500 493.050 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 176.100 490.950 178.200 493.050 ;
        RECT 161.400 489.900 162.600 490.650 ;
        RECT 160.950 487.800 163.050 489.900 ;
        RECT 170.400 489.000 171.600 490.650 ;
        RECT 169.950 484.950 172.050 489.000 ;
        RECT 185.400 487.050 186.450 493.950 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 157.950 478.950 160.050 481.050 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 172.950 457.950 175.050 460.050 ;
        RECT 157.950 449.100 160.050 451.200 ;
        RECT 163.950 449.100 166.050 451.200 ;
        RECT 158.400 448.350 159.600 449.100 ;
        RECT 164.400 448.350 165.600 449.100 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 161.400 444.900 162.600 445.650 ;
        RECT 152.400 443.400 156.450 444.450 ;
        RECT 151.950 436.950 154.050 439.050 ;
        RECT 148.950 433.950 151.050 436.050 ;
        RECT 139.950 421.950 142.050 424.050 ;
        RECT 145.950 421.950 148.050 424.050 ;
        RECT 136.950 416.100 139.050 418.200 ;
        RECT 137.400 415.350 138.600 416.100 ;
        RECT 136.950 412.950 139.050 415.050 ;
        RECT 139.950 412.950 142.050 415.050 ;
        RECT 140.400 411.900 141.600 412.650 ;
        RECT 146.400 412.050 147.450 421.950 ;
        RECT 148.950 416.100 151.050 418.200 ;
        RECT 139.950 409.800 142.050 411.900 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 149.400 388.050 150.450 416.100 ;
        RECT 148.950 385.950 151.050 388.050 ;
        RECT 142.950 382.950 145.050 385.050 ;
        RECT 143.400 372.600 144.450 382.950 ;
        RECT 143.400 370.350 144.600 372.600 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 140.400 365.400 141.600 367.650 ;
        RECT 146.400 366.900 147.600 367.650 ;
        RECT 130.950 361.950 133.050 364.050 ;
        RECT 140.400 361.050 141.450 365.400 ;
        RECT 145.950 364.800 148.050 366.900 ;
        RECT 152.400 364.050 153.450 436.950 ;
        RECT 155.400 417.450 156.450 443.400 ;
        RECT 160.950 442.800 163.050 444.900 ;
        RECT 167.400 444.000 168.600 445.650 ;
        RECT 166.950 439.950 169.050 444.000 ;
        RECT 169.950 442.950 172.050 445.050 ;
        RECT 163.950 424.950 166.050 427.050 ;
        RECT 157.950 417.450 160.050 418.200 ;
        RECT 155.400 416.400 160.050 417.450 ;
        RECT 157.950 416.100 160.050 416.400 ;
        RECT 164.400 417.600 165.450 424.950 ;
        RECT 158.400 415.350 159.600 416.100 ;
        RECT 164.400 415.350 165.600 417.600 ;
        RECT 157.950 412.950 160.050 415.050 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 161.400 411.900 162.600 412.650 ;
        RECT 160.950 409.800 163.050 411.900 ;
        RECT 170.400 394.050 171.450 442.950 ;
        RECT 169.950 391.950 172.050 394.050 ;
        RECT 173.400 375.450 174.450 457.950 ;
        RECT 176.400 451.200 177.450 478.950 ;
        RECT 188.400 454.050 189.450 499.950 ;
        RECT 197.400 499.200 198.450 502.950 ;
        RECT 196.950 497.100 199.050 499.200 ;
        RECT 193.950 493.950 199.050 496.050 ;
        RECT 203.400 495.600 204.450 502.950 ;
        RECT 206.400 496.050 207.450 520.800 ;
        RECT 212.400 514.050 213.450 521.400 ;
        RECT 211.950 511.950 214.050 514.050 ;
        RECT 221.400 511.050 222.450 553.950 ;
        RECT 224.400 523.050 225.450 580.950 ;
        RECT 227.400 559.050 228.450 605.100 ;
        RECT 226.950 556.950 229.050 559.050 ;
        RECT 230.400 529.050 231.450 607.950 ;
        RECT 232.950 604.950 235.050 607.050 ;
        RECT 242.400 606.600 243.450 607.950 ;
        RECT 233.400 600.900 234.450 604.950 ;
        RECT 242.400 604.350 243.600 606.600 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 239.400 600.900 240.600 601.650 ;
        RECT 245.400 600.900 246.600 601.650 ;
        RECT 232.950 598.800 235.050 600.900 ;
        RECT 238.950 598.800 241.050 600.900 ;
        RECT 244.950 598.800 247.050 600.900 ;
        RECT 233.400 592.050 234.450 598.800 ;
        RECT 235.950 595.950 238.050 598.050 ;
        RECT 232.950 589.950 235.050 592.050 ;
        RECT 236.400 574.200 237.450 595.950 ;
        RECT 244.950 580.950 247.050 583.050 ;
        RECT 245.400 576.450 246.450 580.950 ;
        RECT 242.400 575.400 246.450 576.450 ;
        RECT 235.950 572.100 238.050 574.200 ;
        RECT 242.400 573.600 243.450 575.400 ;
        RECT 236.400 571.350 237.600 572.100 ;
        RECT 242.400 571.350 243.600 573.600 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 244.950 568.950 247.050 571.050 ;
        RECT 232.950 565.950 235.050 568.050 ;
        RECT 239.400 567.000 240.600 568.650 ;
        RECT 226.950 526.950 229.050 529.050 ;
        RECT 229.950 526.950 232.050 529.050 ;
        RECT 233.400 528.600 234.450 565.950 ;
        RECT 238.950 562.950 241.050 567.000 ;
        RECT 245.400 566.400 246.600 568.650 ;
        RECT 251.400 567.900 252.450 616.950 ;
        RECT 245.400 553.050 246.450 566.400 ;
        RECT 250.950 565.800 253.050 567.900 ;
        RECT 244.950 550.950 247.050 553.050 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 220.950 508.950 223.050 511.050 ;
        RECT 227.400 504.450 228.450 526.950 ;
        RECT 233.400 526.350 234.600 528.600 ;
        RECT 238.950 528.000 241.050 532.050 ;
        RECT 239.400 526.350 240.600 528.000 ;
        RECT 250.950 526.950 253.050 529.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 236.400 521.400 237.600 523.650 ;
        RECT 242.400 521.400 243.600 523.650 ;
        RECT 232.950 508.950 235.050 511.050 ;
        RECT 229.950 504.450 232.050 505.050 ;
        RECT 227.400 503.400 232.050 504.450 ;
        RECT 229.950 502.950 232.050 503.400 ;
        RECT 197.400 493.350 198.600 493.950 ;
        RECT 203.400 493.350 204.600 495.600 ;
        RECT 205.950 493.950 208.050 496.050 ;
        RECT 220.950 494.100 223.050 496.200 ;
        RECT 221.400 493.350 222.600 494.100 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 191.400 475.050 192.450 490.950 ;
        RECT 200.400 488.400 201.600 490.650 ;
        RECT 224.400 488.400 225.600 490.650 ;
        RECT 200.400 475.050 201.450 488.400 ;
        RECT 224.400 487.050 225.450 488.400 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 223.950 484.950 226.050 487.050 ;
        RECT 190.950 472.950 193.050 475.050 ;
        RECT 199.950 472.950 202.050 475.050 ;
        RECT 211.950 472.950 214.050 475.050 ;
        RECT 187.950 451.950 190.050 454.050 ;
        RECT 175.950 449.100 178.050 451.200 ;
        RECT 184.950 449.100 187.050 451.200 ;
        RECT 191.400 450.600 192.450 472.950 ;
        RECT 199.950 466.950 202.050 469.050 ;
        RECT 196.950 451.950 199.050 454.050 ;
        RECT 176.400 424.050 177.450 449.100 ;
        RECT 185.400 448.350 186.600 449.100 ;
        RECT 191.400 448.350 192.600 450.600 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 190.950 445.950 193.050 448.050 ;
        RECT 188.400 444.900 189.600 445.650 ;
        RECT 187.950 442.800 190.050 444.900 ;
        RECT 184.950 430.950 187.050 433.050 ;
        RECT 175.950 421.950 178.050 424.050 ;
        RECT 176.400 411.450 177.450 421.950 ;
        RECT 185.400 417.600 186.450 430.950 ;
        RECT 185.400 415.350 186.600 417.600 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 176.400 410.400 180.450 411.450 ;
        RECT 170.400 374.400 174.450 375.450 ;
        RECT 157.950 371.100 160.050 373.200 ;
        RECT 163.950 371.100 166.050 373.200 ;
        RECT 170.400 372.600 171.450 374.400 ;
        RECT 158.400 366.450 159.450 371.100 ;
        RECT 164.400 370.350 165.600 371.100 ;
        RECT 170.400 370.350 171.600 372.600 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 158.400 365.400 162.450 366.450 ;
        RECT 142.950 361.950 145.050 364.050 ;
        RECT 151.950 361.950 154.050 364.050 ;
        RECT 139.950 358.950 142.050 361.050 ;
        RECT 127.950 349.950 130.050 352.050 ;
        RECT 128.400 339.600 129.450 349.950 ;
        RECT 136.950 346.950 139.050 349.050 ;
        RECT 128.400 337.350 129.600 339.600 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 131.400 333.900 132.600 334.650 ;
        RECT 130.950 331.800 133.050 333.900 ;
        RECT 137.400 325.050 138.450 346.950 ;
        RECT 139.950 338.100 142.050 340.200 ;
        RECT 140.400 334.050 141.450 338.100 ;
        RECT 139.950 331.950 142.050 334.050 ;
        RECT 136.950 322.950 139.050 325.050 ;
        RECT 118.950 307.950 121.050 310.050 ;
        RECT 119.400 288.900 120.450 307.950 ;
        RECT 124.950 293.100 127.050 295.200 ;
        RECT 130.950 293.100 133.050 295.200 ;
        RECT 125.400 292.350 126.600 293.100 ;
        RECT 131.400 292.350 132.600 293.100 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 118.950 286.800 121.050 288.900 ;
        RECT 128.400 287.400 129.600 289.650 ;
        RECT 134.400 287.400 135.600 289.650 ;
        RECT 115.950 280.950 118.050 283.050 ;
        RECT 128.400 274.050 129.450 287.400 ;
        RECT 134.400 286.050 135.450 287.400 ;
        RECT 133.950 283.950 136.050 286.050 ;
        RECT 127.950 271.950 130.050 274.050 ;
        RECT 115.950 262.950 118.050 265.050 ;
        RECT 112.950 253.950 115.050 256.050 ;
        RECT 109.950 238.950 112.050 241.050 ;
        RECT 116.400 232.050 117.450 262.950 ;
        RECT 118.950 260.100 121.050 262.200 ;
        RECT 127.950 260.100 130.050 262.200 ;
        RECT 119.400 235.050 120.450 260.100 ;
        RECT 128.400 259.350 129.600 260.100 ;
        RECT 122.100 256.950 124.200 259.050 ;
        RECT 127.500 256.950 129.600 259.050 ;
        RECT 130.800 256.950 132.900 259.050 ;
        RECT 122.400 254.400 123.600 256.650 ;
        RECT 131.400 254.400 132.600 256.650 ;
        RECT 118.950 232.950 121.050 235.050 ;
        RECT 115.950 229.950 118.050 232.050 ;
        RECT 122.400 229.050 123.450 254.400 ;
        RECT 127.950 244.950 130.050 247.050 ;
        RECT 121.950 226.950 124.050 229.050 ;
        RECT 124.950 220.950 127.050 223.050 ;
        RECT 112.950 215.100 115.050 217.200 ;
        RECT 120.000 216.600 124.050 217.050 ;
        RECT 113.400 214.350 114.600 215.100 ;
        RECT 119.400 214.950 124.050 216.600 ;
        RECT 119.400 214.350 120.600 214.950 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 116.400 210.900 117.600 211.650 ;
        RECT 125.400 211.050 126.450 220.950 ;
        RECT 115.950 208.800 118.050 210.900 ;
        RECT 121.950 208.950 124.050 211.050 ;
        RECT 124.950 208.950 127.050 211.050 ;
        RECT 122.400 205.050 123.450 208.950 ;
        RECT 115.950 202.950 118.050 205.050 ;
        RECT 121.950 202.950 124.050 205.050 ;
        RECT 116.400 183.600 117.450 202.950 ;
        RECT 116.400 181.350 117.600 183.600 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 113.400 176.400 114.600 178.650 ;
        RECT 119.400 176.400 120.600 178.650 ;
        RECT 109.950 172.950 112.050 175.050 ;
        RECT 106.950 166.950 109.050 169.050 ;
        RECT 100.950 145.950 103.050 148.050 ;
        RECT 97.950 137.100 100.050 139.200 ;
        RECT 105.000 138.600 109.050 139.050 ;
        RECT 98.400 136.350 99.600 137.100 ;
        RECT 104.400 136.950 109.050 138.600 ;
        RECT 104.400 136.350 105.600 136.950 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 101.400 132.900 102.600 133.650 ;
        RECT 100.950 130.800 103.050 132.900 ;
        RECT 110.400 129.450 111.450 172.950 ;
        RECT 113.400 133.050 114.450 176.400 ;
        RECT 119.400 157.050 120.450 176.400 ;
        RECT 128.400 175.050 129.450 244.950 ;
        RECT 131.400 244.050 132.450 254.400 ;
        RECT 134.400 247.050 135.450 283.950 ;
        RECT 136.950 277.950 139.050 280.050 ;
        RECT 137.400 256.050 138.450 277.950 ;
        RECT 136.950 253.950 139.050 256.050 ;
        RECT 133.950 244.950 136.050 247.050 ;
        RECT 130.950 241.950 133.050 244.050 ;
        RECT 133.950 235.950 136.050 238.050 ;
        RECT 130.950 226.950 133.050 229.050 ;
        RECT 131.400 205.050 132.450 226.950 ;
        RECT 134.400 217.050 135.450 235.950 ;
        RECT 140.400 223.050 141.450 331.950 ;
        RECT 143.400 256.050 144.450 361.950 ;
        RECT 148.950 338.100 151.050 340.200 ;
        RECT 156.000 339.600 160.050 340.050 ;
        RECT 149.400 337.350 150.600 338.100 ;
        RECT 155.400 337.950 160.050 339.600 ;
        RECT 155.400 337.350 156.600 337.950 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 152.400 333.900 153.600 334.650 ;
        RECT 161.400 334.050 162.450 365.400 ;
        RECT 167.400 365.400 168.600 367.650 ;
        RECT 173.400 366.900 174.600 367.650 ;
        RECT 167.400 361.050 168.450 365.400 ;
        RECT 172.950 364.800 175.050 366.900 ;
        RECT 179.400 361.050 180.450 410.400 ;
        RECT 182.400 410.400 183.600 412.650 ;
        RECT 188.400 411.900 189.600 412.650 ;
        RECT 182.400 391.050 183.450 410.400 ;
        RECT 187.950 409.800 190.050 411.900 ;
        RECT 187.950 403.950 190.050 406.050 ;
        RECT 190.950 403.950 193.050 406.050 ;
        RECT 184.950 397.950 187.050 400.050 ;
        RECT 181.950 388.950 184.050 391.050 ;
        RECT 185.400 384.450 186.450 397.950 ;
        RECT 188.400 385.050 189.450 403.950 ;
        RECT 182.400 383.400 186.450 384.450 ;
        RECT 166.950 358.950 169.050 361.050 ;
        RECT 172.950 358.950 175.050 361.050 ;
        RECT 178.950 358.950 181.050 361.050 ;
        RECT 173.400 340.200 174.450 358.950 ;
        RECT 182.400 346.050 183.450 383.400 ;
        RECT 187.950 382.950 190.050 385.050 ;
        RECT 184.950 370.950 187.050 373.050 ;
        RECT 191.400 372.600 192.450 403.950 ;
        RECT 197.400 373.050 198.450 451.950 ;
        RECT 185.400 366.900 186.450 370.950 ;
        RECT 191.400 370.350 192.600 372.600 ;
        RECT 196.950 370.950 199.050 373.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 184.950 364.800 187.050 366.900 ;
        RECT 194.400 365.400 195.600 367.650 ;
        RECT 194.400 364.050 195.450 365.400 ;
        RECT 200.400 364.050 201.450 466.950 ;
        RECT 212.400 460.050 213.450 472.950 ;
        RECT 224.400 469.050 225.450 484.950 ;
        RECT 223.950 466.950 226.050 469.050 ;
        RECT 211.950 457.950 214.050 460.050 ;
        RECT 217.950 449.100 220.050 451.200 ;
        RECT 223.950 449.100 226.050 451.200 ;
        RECT 218.400 448.350 219.600 449.100 ;
        RECT 212.100 445.950 214.200 448.050 ;
        RECT 218.100 445.950 220.200 448.050 ;
        RECT 220.950 439.950 223.050 442.050 ;
        RECT 217.950 433.950 220.050 436.050 ;
        RECT 208.950 427.950 211.050 430.050 ;
        RECT 209.400 417.600 210.450 427.950 ;
        RECT 214.950 424.950 217.050 427.050 ;
        RECT 215.400 417.600 216.450 424.950 ;
        RECT 218.400 418.050 219.450 433.950 ;
        RECT 209.400 415.350 210.600 417.600 ;
        RECT 215.400 415.350 216.600 417.600 ;
        RECT 217.950 415.950 220.050 418.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 208.950 412.950 211.050 415.050 ;
        RECT 211.950 412.950 214.050 415.050 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 206.400 410.400 207.600 412.650 ;
        RECT 212.400 411.900 213.600 412.650 ;
        RECT 206.400 406.050 207.450 410.400 ;
        RECT 211.950 409.800 214.050 411.900 ;
        RECT 217.950 409.950 220.050 412.050 ;
        RECT 205.950 403.950 208.050 406.050 ;
        RECT 211.950 379.950 214.050 382.050 ;
        RECT 205.950 370.950 208.050 373.050 ;
        RECT 212.400 372.600 213.450 379.950 ;
        RECT 218.400 373.050 219.450 409.950 ;
        RECT 193.950 361.950 196.050 364.050 ;
        RECT 199.950 361.950 202.050 364.050 ;
        RECT 181.950 343.950 184.050 346.050 ;
        RECT 163.950 337.950 166.050 340.050 ;
        RECT 166.950 337.950 169.050 340.050 ;
        RECT 172.950 338.100 175.050 340.200 ;
        RECT 151.950 331.800 154.050 333.900 ;
        RECT 160.950 331.950 163.050 334.050 ;
        RECT 154.950 301.950 157.050 304.050 ;
        RECT 155.400 294.600 156.450 301.950 ;
        RECT 164.400 300.450 165.450 337.950 ;
        RECT 167.400 334.050 168.450 337.950 ;
        RECT 173.400 337.350 174.600 338.100 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 166.950 333.450 169.050 334.050 ;
        RECT 176.400 333.900 177.600 334.650 ;
        RECT 166.950 332.400 171.450 333.450 ;
        RECT 166.950 331.950 169.050 332.400 ;
        RECT 164.400 299.400 168.450 300.450 ;
        RECT 155.400 292.350 156.600 294.600 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 157.950 289.950 160.050 292.050 ;
        RECT 152.400 287.400 153.600 289.650 ;
        RECT 158.400 288.000 159.600 289.650 ;
        RECT 152.400 277.050 153.450 287.400 ;
        RECT 157.950 283.950 160.050 288.000 ;
        RECT 151.950 274.950 154.050 277.050 ;
        RECT 148.950 261.000 151.050 265.050 ;
        RECT 149.400 259.350 150.600 261.000 ;
        RECT 154.950 260.100 157.050 262.200 ;
        RECT 155.400 259.350 156.600 260.100 ;
        RECT 160.950 259.950 163.050 262.050 ;
        RECT 163.950 260.100 166.050 262.200 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 142.950 253.950 145.050 256.050 ;
        RECT 145.950 253.950 148.050 256.050 ;
        RECT 152.400 255.900 153.600 256.650 ;
        RECT 139.950 220.950 142.050 223.050 ;
        RECT 146.400 220.050 147.450 253.950 ;
        RECT 151.950 253.800 154.050 255.900 ;
        RECT 161.400 235.050 162.450 259.950 ;
        RECT 160.950 232.950 163.050 235.050 ;
        RECT 148.950 229.950 151.050 232.050 ;
        RECT 164.400 231.450 165.450 260.100 ;
        RECT 161.400 230.400 165.450 231.450 ;
        RECT 145.950 217.950 148.050 220.050 ;
        RECT 133.950 214.950 136.050 217.050 ;
        RECT 139.950 215.100 142.050 217.200 ;
        RECT 146.400 216.450 147.600 216.600 ;
        RECT 149.400 216.450 150.450 229.950 ;
        RECT 154.950 220.950 157.050 223.050 ;
        RECT 157.950 220.950 160.050 223.050 ;
        RECT 146.400 215.400 150.450 216.450 ;
        RECT 140.400 214.350 141.600 215.100 ;
        RECT 146.400 214.350 147.600 215.400 ;
        RECT 151.950 215.100 154.050 217.200 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 145.950 211.950 148.050 214.050 ;
        RECT 137.400 210.900 138.600 211.650 ;
        RECT 136.950 208.800 139.050 210.900 ;
        RECT 143.400 209.400 144.600 211.650 ;
        RECT 152.400 210.450 153.450 215.100 ;
        RECT 149.400 209.400 153.450 210.450 ;
        RECT 143.400 205.050 144.450 209.400 ;
        RECT 130.950 202.950 133.050 205.050 ;
        RECT 142.950 202.950 145.050 205.050 ;
        RECT 131.400 175.050 132.450 202.950 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 140.400 183.600 141.450 196.950 ;
        RECT 140.400 181.350 141.600 183.600 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 137.400 177.000 138.600 178.650 ;
        RECT 143.400 177.000 144.600 178.650 ;
        RECT 121.950 172.950 124.050 175.050 ;
        RECT 127.950 172.950 130.050 175.050 ;
        RECT 130.950 172.950 133.050 175.050 ;
        RECT 136.950 172.950 139.050 177.000 ;
        RECT 142.950 172.950 145.050 177.000 ;
        RECT 118.950 154.950 121.050 157.050 ;
        RECT 118.950 145.950 121.050 148.050 ;
        RECT 115.950 136.950 118.050 139.050 ;
        RECT 116.400 133.050 117.450 136.950 ;
        RECT 112.800 130.950 114.900 133.050 ;
        RECT 115.950 130.950 118.050 133.050 ;
        RECT 110.400 128.400 114.450 129.450 ;
        RECT 91.950 124.950 94.050 127.050 ;
        RECT 100.950 124.950 103.050 127.050 ;
        RECT 94.950 109.950 97.050 112.050 ;
        RECT 95.400 105.600 96.450 109.950 ;
        RECT 101.400 105.600 102.450 124.950 ;
        RECT 109.950 109.950 112.050 112.050 ;
        RECT 95.400 103.350 96.600 105.600 ;
        RECT 101.400 103.350 102.600 105.600 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 92.400 99.900 93.600 100.650 ;
        RECT 91.950 97.800 94.050 99.900 ;
        RECT 98.400 99.000 99.600 100.650 ;
        RECT 92.400 64.050 93.450 97.800 ;
        RECT 97.950 94.950 100.050 99.000 ;
        RECT 91.950 61.950 94.050 64.050 ;
        RECT 88.950 58.950 91.050 61.050 ;
        RECT 94.950 60.000 97.050 64.050 ;
        RECT 100.950 60.000 103.050 64.050 ;
        RECT 85.950 49.950 88.050 52.050 ;
        RECT 64.950 31.950 67.050 34.050 ;
        RECT 65.400 27.600 66.450 31.950 ;
        RECT 82.950 28.950 85.050 31.050 ;
        RECT 65.400 25.350 66.600 27.600 ;
        RECT 65.400 22.950 67.500 25.050 ;
        RECT 70.800 22.950 72.900 25.050 ;
        RECT 83.400 22.050 84.450 28.950 ;
        RECT 89.400 27.600 90.450 58.950 ;
        RECT 95.400 58.350 96.600 60.000 ;
        RECT 101.400 58.350 102.600 60.000 ;
        RECT 94.950 55.950 97.050 58.050 ;
        RECT 97.950 55.950 100.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 98.400 53.400 99.600 55.650 ;
        RECT 104.400 54.900 105.600 55.650 ;
        RECT 98.400 49.050 99.450 53.400 ;
        RECT 103.950 52.800 106.050 54.900 ;
        RECT 97.950 46.950 100.050 49.050 ;
        RECT 110.400 46.050 111.450 109.950 ;
        RECT 113.400 55.050 114.450 128.400 ;
        RECT 119.400 127.050 120.450 145.950 ;
        RECT 122.400 138.600 123.450 172.950 ;
        RECT 139.950 169.950 142.050 172.050 ;
        RECT 122.400 136.350 123.600 138.600 ;
        RECT 130.950 138.450 133.050 139.200 ;
        RECT 130.950 137.400 135.450 138.450 ;
        RECT 130.950 137.100 133.050 137.400 ;
        RECT 131.400 136.350 132.600 137.100 ;
        RECT 122.100 133.950 124.200 136.050 ;
        RECT 125.400 133.950 127.500 136.050 ;
        RECT 130.800 133.950 132.900 136.050 ;
        RECT 125.400 132.900 126.600 133.650 ;
        RECT 134.400 133.050 135.450 137.400 ;
        RECT 124.950 130.800 127.050 132.900 ;
        RECT 133.950 130.950 136.050 133.050 ;
        RECT 118.950 124.950 121.050 127.050 ;
        RECT 125.400 112.050 126.450 130.800 ;
        RECT 140.400 130.050 141.450 169.950 ;
        RECT 127.950 127.950 130.050 130.050 ;
        RECT 139.950 127.950 142.050 130.050 ;
        RECT 124.950 109.950 127.050 112.050 ;
        RECT 128.400 111.450 129.450 127.950 ;
        RECT 128.400 109.200 129.600 111.450 ;
        RECT 123.900 105.900 126.000 107.700 ;
        RECT 127.800 106.800 129.900 108.900 ;
        RECT 131.100 108.300 133.200 110.400 ;
        RECT 122.400 104.700 131.100 105.900 ;
        RECT 119.100 100.950 121.200 103.050 ;
        RECT 119.400 99.900 120.600 100.650 ;
        RECT 118.950 97.800 121.050 99.900 ;
        RECT 122.400 95.700 123.300 104.700 ;
        RECT 129.000 103.800 131.100 104.700 ;
        RECT 132.000 102.900 132.900 108.300 ;
        RECT 133.950 104.100 136.050 106.200 ;
        RECT 139.950 104.100 142.050 106.200 ;
        RECT 134.400 103.350 135.600 104.100 ;
        RECT 126.000 101.700 132.900 102.900 ;
        RECT 126.000 99.300 126.900 101.700 ;
        RECT 124.800 97.200 126.900 99.300 ;
        RECT 127.800 97.950 129.900 100.050 ;
        RECT 121.500 93.600 123.600 95.700 ;
        RECT 128.400 95.400 129.600 97.650 ;
        RECT 131.700 94.500 132.900 101.700 ;
        RECT 133.800 100.950 135.900 103.050 ;
        RECT 131.100 92.400 133.200 94.500 ;
        RECT 115.950 67.950 118.050 70.050 ;
        RECT 136.950 67.950 139.050 70.050 ;
        RECT 112.800 52.950 114.900 55.050 ;
        RECT 116.400 54.900 117.450 67.950 ;
        RECT 124.950 59.100 127.050 61.200 ;
        RECT 125.400 58.350 126.600 59.100 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 122.400 54.900 123.600 55.650 ;
        RECT 115.950 52.800 118.050 54.900 ;
        RECT 121.950 52.800 124.050 54.900 ;
        RECT 128.400 54.000 129.600 55.650 ;
        RECT 127.950 49.950 130.050 54.000 ;
        RECT 112.950 46.950 115.050 49.050 ;
        RECT 94.950 43.950 97.050 46.050 ;
        RECT 109.950 43.950 112.050 46.050 ;
        RECT 95.400 27.600 96.450 43.950 ;
        RECT 109.950 28.950 112.050 31.050 ;
        RECT 89.400 25.350 90.600 27.600 ;
        RECT 95.400 25.350 96.600 27.600 ;
        RECT 103.950 25.950 106.050 28.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 97.950 22.950 100.050 25.050 ;
        RECT 52.950 19.800 55.050 21.900 ;
        RECT 82.950 19.950 85.050 22.050 ;
        RECT 92.400 21.900 93.600 22.650 ;
        RECT 98.400 21.900 99.600 22.650 ;
        RECT 104.400 21.900 105.450 25.950 ;
        RECT 110.400 21.900 111.450 28.950 ;
        RECT 91.950 19.800 94.050 21.900 ;
        RECT 97.950 19.800 100.050 21.900 ;
        RECT 103.950 19.800 106.050 21.900 ;
        RECT 109.950 19.800 112.050 21.900 ;
        RECT 113.400 21.450 114.450 46.950 ;
        RECT 118.950 26.100 121.050 28.200 ;
        RECT 119.400 25.350 120.600 26.100 ;
        RECT 116.100 22.950 118.200 25.050 ;
        RECT 119.400 22.950 121.500 25.050 ;
        RECT 124.800 22.950 126.900 25.050 ;
        RECT 116.400 21.450 117.600 22.650 ;
        RECT 125.400 21.900 126.600 22.650 ;
        RECT 137.400 21.900 138.450 67.950 ;
        RECT 140.400 67.050 141.450 104.100 ;
        RECT 143.400 70.050 144.450 172.950 ;
        RECT 149.400 172.050 150.450 209.400 ;
        RECT 155.400 175.050 156.450 220.950 ;
        RECT 158.400 210.900 159.450 220.950 ;
        RECT 161.400 217.050 162.450 230.400 ;
        RECT 167.400 229.050 168.450 299.400 ;
        RECT 170.400 262.050 171.450 332.400 ;
        RECT 175.950 331.800 178.050 333.900 ;
        RECT 182.400 316.050 183.450 343.950 ;
        RECT 194.400 340.200 195.450 361.950 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 187.950 338.100 190.050 340.200 ;
        RECT 193.950 338.100 196.050 340.200 ;
        RECT 200.400 339.600 201.450 343.950 ;
        RECT 188.400 333.450 189.450 338.100 ;
        RECT 194.400 337.350 195.600 338.100 ;
        RECT 200.400 337.350 201.600 339.600 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 188.400 332.400 192.450 333.450 ;
        RECT 181.950 313.950 184.050 316.050 ;
        RECT 178.950 293.100 181.050 295.200 ;
        RECT 184.950 293.100 187.050 295.200 ;
        RECT 179.400 292.350 180.600 293.100 ;
        RECT 185.400 292.350 186.600 293.100 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 176.400 288.900 177.600 289.650 ;
        RECT 175.950 286.800 178.050 288.900 ;
        RECT 182.400 287.400 183.600 289.650 ;
        RECT 175.950 280.950 178.050 283.050 ;
        RECT 169.950 259.950 172.050 262.050 ;
        RECT 176.400 261.600 177.450 280.950 ;
        RECT 182.400 280.050 183.450 287.400 ;
        RECT 181.950 277.950 184.050 280.050 ;
        RECT 191.400 265.050 192.450 332.400 ;
        RECT 197.400 332.400 198.600 334.650 ;
        RECT 206.400 334.050 207.450 370.950 ;
        RECT 212.400 370.350 213.600 372.600 ;
        RECT 217.950 370.950 220.050 373.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 215.400 365.400 216.600 367.650 ;
        RECT 215.400 339.450 216.450 365.400 ;
        RECT 221.400 349.050 222.450 439.950 ;
        RECT 224.400 421.050 225.450 449.100 ;
        RECT 223.950 418.950 226.050 421.050 ;
        RECT 223.950 415.800 226.050 417.900 ;
        RECT 224.400 373.050 225.450 415.800 ;
        RECT 223.950 370.950 226.050 373.050 ;
        RECT 223.950 367.800 226.050 369.900 ;
        RECT 224.400 358.050 225.450 367.800 ;
        RECT 223.950 355.950 226.050 358.050 ;
        RECT 220.950 346.950 223.050 349.050 ;
        RECT 212.400 338.400 216.450 339.450 ;
        RECT 221.400 339.600 222.450 346.950 ;
        RECT 227.400 343.050 228.450 487.950 ;
        RECT 230.400 487.050 231.450 502.950 ;
        RECT 229.950 484.950 232.050 487.050 ;
        RECT 229.950 460.950 232.050 463.050 ;
        RECT 230.400 418.050 231.450 460.950 ;
        RECT 233.400 421.050 234.450 508.950 ;
        RECT 236.400 496.200 237.450 521.400 ;
        RECT 242.400 499.050 243.450 521.400 ;
        RECT 241.950 496.950 244.050 499.050 ;
        RECT 235.950 494.100 238.050 496.200 ;
        RECT 244.950 494.100 247.050 496.200 ;
        RECT 251.400 496.050 252.450 526.950 ;
        RECT 254.400 502.050 255.450 628.950 ;
        RECT 262.950 616.950 265.050 619.050 ;
        RECT 256.950 607.950 259.050 610.050 ;
        RECT 257.400 600.900 258.450 607.950 ;
        RECT 263.400 606.600 264.450 616.950 ;
        RECT 269.400 610.200 270.450 649.950 ;
        RECT 278.400 649.350 279.600 650.100 ;
        RECT 284.400 649.350 285.600 651.600 ;
        RECT 289.950 649.950 292.050 653.400 ;
        RECT 277.950 646.950 280.050 649.050 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 281.400 645.000 282.600 646.650 ;
        RECT 287.400 645.900 288.600 646.650 ;
        RECT 293.400 645.900 294.450 655.950 ;
        RECT 295.950 649.950 298.050 652.050 ;
        RECT 280.950 640.950 283.050 645.000 ;
        RECT 286.950 643.800 289.050 645.900 ;
        RECT 292.950 643.800 295.050 645.900 ;
        RECT 283.950 610.950 286.050 613.050 ;
        RECT 268.950 608.100 271.050 610.200 ;
        RECT 263.400 604.350 264.600 606.600 ;
        RECT 268.950 604.950 271.050 607.050 ;
        RECT 280.950 605.100 283.050 607.200 ;
        RECT 269.400 604.350 270.600 604.950 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 266.400 600.900 267.600 601.650 ;
        RECT 256.950 598.800 259.050 600.900 ;
        RECT 265.950 598.800 268.050 600.900 ;
        RECT 272.400 599.400 273.600 601.650 ;
        RECT 266.400 573.600 267.450 598.800 ;
        RECT 272.400 586.050 273.450 599.400 ;
        RECT 271.950 583.950 274.050 586.050 ;
        RECT 266.400 571.350 267.600 573.600 ;
        RECT 271.950 573.000 274.050 577.050 ;
        RECT 277.950 574.950 280.050 577.050 ;
        RECT 272.400 571.350 273.600 573.000 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 263.400 567.900 264.600 568.650 ;
        RECT 269.400 567.900 270.600 568.650 ;
        RECT 262.950 565.800 265.050 567.900 ;
        RECT 268.950 565.800 271.050 567.900 ;
        RECT 259.950 562.950 262.050 565.050 ;
        RECT 260.400 547.050 261.450 562.950 ;
        RECT 278.400 553.050 279.450 574.950 ;
        RECT 281.400 574.200 282.450 605.100 ;
        RECT 280.950 572.100 283.050 574.200 ;
        RECT 274.950 550.950 277.050 553.050 ;
        RECT 277.950 550.950 280.050 553.050 ;
        RECT 259.950 544.950 262.050 547.050 ;
        RECT 256.950 541.950 259.050 544.050 ;
        RECT 257.400 532.050 258.450 541.950 ;
        RECT 271.950 538.950 274.050 541.050 ;
        RECT 262.950 535.950 265.050 538.050 ;
        RECT 256.950 529.950 259.050 532.050 ;
        RECT 263.400 528.600 264.450 535.950 ;
        RECT 263.400 526.350 264.600 528.600 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 260.400 521.400 261.600 523.650 ;
        RECT 266.400 521.400 267.600 523.650 ;
        RECT 272.400 523.050 273.450 538.950 ;
        RECT 260.400 517.050 261.450 521.400 ;
        RECT 259.950 514.950 262.050 517.050 ;
        RECT 266.400 505.050 267.450 521.400 ;
        RECT 271.950 520.950 274.050 523.050 ;
        RECT 271.950 508.950 274.050 511.050 ;
        RECT 265.950 502.950 268.050 505.050 ;
        RECT 253.950 499.950 256.050 502.050 ;
        RECT 265.950 499.800 268.050 501.900 ;
        RECT 253.950 496.800 256.050 498.900 ;
        RECT 245.400 493.350 246.600 494.100 ;
        RECT 250.950 493.950 253.050 496.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 242.400 489.900 243.600 490.650 ;
        RECT 241.950 487.800 244.050 489.900 ;
        RECT 248.400 488.400 249.600 490.650 ;
        RECT 254.400 489.900 255.450 496.800 ;
        RECT 266.400 496.200 267.450 499.800 ;
        RECT 259.950 493.950 262.050 496.050 ;
        RECT 265.950 494.100 268.050 496.200 ;
        RECT 272.400 495.600 273.450 508.950 ;
        RECT 248.400 481.050 249.450 488.400 ;
        RECT 253.950 487.800 256.050 489.900 ;
        RECT 247.950 478.950 250.050 481.050 ;
        RECT 241.950 449.100 244.050 451.200 ;
        RECT 247.950 449.100 250.050 451.200 ;
        RECT 242.400 448.350 243.600 449.100 ;
        RECT 248.400 448.350 249.600 449.100 ;
        RECT 238.950 445.950 241.050 448.050 ;
        RECT 241.950 445.950 244.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 239.400 443.400 240.600 445.650 ;
        RECT 245.400 443.400 246.600 445.650 ;
        RECT 235.950 423.450 238.050 424.050 ;
        RECT 239.400 423.450 240.450 443.400 ;
        RECT 245.400 427.050 246.450 443.400 ;
        RECT 250.950 442.950 253.050 445.050 ;
        RECT 247.950 427.950 250.050 430.050 ;
        RECT 241.950 424.950 244.050 427.050 ;
        RECT 244.950 424.950 247.050 427.050 ;
        RECT 235.950 422.400 240.450 423.450 ;
        RECT 235.950 421.950 238.050 422.400 ;
        RECT 232.950 418.950 235.050 421.050 ;
        RECT 229.950 415.950 232.050 418.050 ;
        RECT 236.400 417.600 237.450 421.950 ;
        RECT 242.400 417.600 243.450 424.950 ;
        RECT 236.400 415.350 237.600 417.600 ;
        RECT 242.400 415.350 243.600 417.600 ;
        RECT 232.950 412.950 235.050 415.050 ;
        RECT 235.950 412.950 238.050 415.050 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 233.400 411.900 234.600 412.650 ;
        RECT 239.400 411.900 240.600 412.650 ;
        RECT 230.400 373.050 231.450 409.950 ;
        RECT 232.950 409.800 235.050 411.900 ;
        RECT 238.950 409.800 241.050 411.900 ;
        RECT 233.400 400.050 234.450 409.800 ;
        RECT 232.950 397.950 235.050 400.050 ;
        RECT 248.400 391.050 249.450 427.950 ;
        RECT 251.400 412.050 252.450 442.950 ;
        RECT 254.400 427.050 255.450 487.800 ;
        RECT 260.400 484.050 261.450 493.950 ;
        RECT 266.400 493.350 267.600 494.100 ;
        RECT 272.400 493.350 273.600 495.600 ;
        RECT 275.400 495.450 276.450 550.950 ;
        RECT 281.400 541.050 282.450 572.100 ;
        RECT 284.400 553.050 285.450 610.950 ;
        RECT 296.400 607.200 297.450 649.950 ;
        RECT 299.400 613.050 300.450 683.400 ;
        RECT 313.950 683.100 316.050 685.200 ;
        RECT 320.400 684.600 321.450 727.950 ;
        RECT 326.400 727.350 327.600 729.000 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 329.400 723.900 330.600 724.650 ;
        RECT 328.950 721.800 331.050 723.900 ;
        RECT 335.400 723.450 336.450 775.950 ;
        RECT 337.950 762.000 340.050 766.050 ;
        RECT 347.400 765.450 348.450 811.950 ;
        RECT 355.950 806.100 358.050 808.200 ;
        RECT 362.400 807.600 363.450 817.950 ;
        RECT 368.400 814.050 369.450 820.950 ;
        RECT 367.950 811.950 370.050 814.050 ;
        RECT 391.950 811.950 394.050 814.050 ;
        RECT 373.950 808.950 376.050 811.050 ;
        RECT 356.400 805.350 357.600 806.100 ;
        RECT 362.400 805.350 363.600 807.600 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 361.950 802.950 364.050 805.050 ;
        RECT 353.400 800.400 354.600 802.650 ;
        RECT 359.400 801.900 360.600 802.650 ;
        RECT 353.400 796.050 354.450 800.400 ;
        RECT 358.950 799.800 361.050 801.900 ;
        RECT 367.950 799.800 370.050 801.900 ;
        RECT 359.400 798.450 360.450 799.800 ;
        RECT 359.400 797.400 363.450 798.450 ;
        RECT 352.950 793.950 355.050 796.050 ;
        RECT 358.950 793.950 361.050 796.050 ;
        RECT 353.400 790.050 354.450 793.950 ;
        RECT 352.950 787.950 355.050 790.050 ;
        RECT 347.400 764.400 351.450 765.450 ;
        RECT 338.400 760.350 339.600 762.000 ;
        RECT 346.950 761.100 349.050 763.200 ;
        RECT 347.400 760.350 348.600 761.100 ;
        RECT 338.100 757.950 340.200 760.050 ;
        RECT 343.500 757.950 345.600 760.050 ;
        RECT 346.800 757.950 348.900 760.050 ;
        RECT 344.400 755.400 345.600 757.650 ;
        RECT 344.400 745.050 345.450 755.400 ;
        RECT 343.950 742.950 346.050 745.050 ;
        RECT 350.400 736.050 351.450 764.400 ;
        RECT 355.950 763.950 358.050 766.050 ;
        RECT 352.950 761.100 355.050 763.200 ;
        RECT 353.400 748.050 354.450 761.100 ;
        RECT 356.400 756.900 357.450 763.950 ;
        RECT 355.950 754.800 358.050 756.900 ;
        RECT 352.950 745.950 355.050 748.050 ;
        RECT 352.950 739.950 355.050 742.050 ;
        RECT 340.950 733.950 343.050 736.050 ;
        RECT 349.950 733.950 352.050 736.050 ;
        RECT 337.950 728.100 340.050 730.200 ;
        RECT 332.400 722.400 336.450 723.450 ;
        RECT 325.950 697.950 328.050 700.050 ;
        RECT 322.950 691.950 325.050 694.050 ;
        RECT 323.400 685.050 324.450 691.950 ;
        RECT 314.400 682.350 315.600 683.100 ;
        RECT 320.400 682.350 321.600 684.600 ;
        RECT 322.950 682.950 325.050 685.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 311.400 677.400 312.600 679.650 ;
        RECT 317.400 678.900 318.600 679.650 ;
        RECT 311.400 661.050 312.450 677.400 ;
        RECT 316.950 676.800 319.050 678.900 ;
        RECT 310.950 658.950 313.050 661.050 ;
        RECT 319.950 658.950 322.050 661.050 ;
        RECT 304.950 650.100 307.050 652.200 ;
        RECT 310.950 651.000 313.050 655.050 ;
        RECT 305.400 649.350 306.600 650.100 ;
        RECT 311.400 649.350 312.600 651.000 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 307.950 646.950 310.050 649.050 ;
        RECT 310.950 646.950 313.050 649.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 308.400 645.000 309.600 646.650 ;
        RECT 314.400 645.900 315.600 646.650 ;
        RECT 307.950 640.950 310.050 645.000 ;
        RECT 313.950 643.800 316.050 645.900 ;
        RECT 310.950 634.950 313.050 637.050 ;
        RECT 298.950 610.950 301.050 613.050 ;
        RECT 289.950 605.100 292.050 607.200 ;
        RECT 295.950 605.100 298.050 607.200 ;
        RECT 290.400 604.350 291.600 605.100 ;
        RECT 296.400 604.350 297.600 605.100 ;
        RECT 304.950 604.950 307.050 607.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 293.400 600.000 294.600 601.650 ;
        RECT 292.950 595.950 295.050 600.000 ;
        RECT 299.400 599.400 300.600 601.650 ;
        RECT 292.950 572.100 295.050 574.200 ;
        RECT 293.400 571.350 294.600 572.100 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 290.400 567.900 291.600 568.650 ;
        RECT 289.950 565.800 292.050 567.900 ;
        RECT 289.950 556.950 292.050 559.050 ;
        RECT 283.950 550.950 286.050 553.050 ;
        RECT 280.950 538.950 283.050 541.050 ;
        RECT 277.950 529.950 280.050 532.050 ;
        RECT 278.400 499.050 279.450 529.950 ;
        RECT 283.950 528.000 286.050 532.050 ;
        RECT 290.400 528.600 291.450 556.950 ;
        RECT 295.950 547.950 298.050 550.050 ;
        RECT 296.400 528.600 297.450 547.950 ;
        RECT 299.400 532.050 300.450 599.400 ;
        RECT 305.400 565.050 306.450 604.950 ;
        RECT 311.400 600.900 312.450 634.950 ;
        RECT 320.400 606.600 321.450 658.950 ;
        RECT 326.400 655.050 327.450 697.950 ;
        RECT 328.950 684.450 331.050 685.050 ;
        RECT 332.400 684.450 333.450 722.400 ;
        RECT 338.400 712.050 339.450 728.100 ;
        RECT 337.950 711.450 340.050 712.050 ;
        RECT 328.950 683.400 333.450 684.450 ;
        RECT 335.400 710.400 340.050 711.450 ;
        RECT 328.950 682.950 331.050 683.400 ;
        RECT 329.400 658.050 330.450 682.950 ;
        RECT 335.400 678.900 336.450 710.400 ;
        RECT 337.950 709.950 340.050 710.400 ;
        RECT 341.400 688.050 342.450 733.950 ;
        RECT 346.950 728.100 349.050 730.200 ;
        RECT 353.400 729.600 354.450 739.950 ;
        RECT 359.400 730.050 360.450 793.950 ;
        RECT 362.400 787.050 363.450 797.400 ;
        RECT 364.950 796.950 367.050 799.050 ;
        RECT 365.400 790.050 366.450 796.950 ;
        RECT 364.950 787.950 367.050 790.050 ;
        RECT 361.950 784.950 364.050 787.050 ;
        RECT 368.400 762.600 369.450 799.800 ;
        RECT 374.400 778.050 375.450 808.950 ;
        RECT 382.950 807.000 385.050 811.050 ;
        RECT 388.950 807.000 391.050 811.050 ;
        RECT 392.400 808.050 393.450 811.950 ;
        RECT 383.400 805.350 384.600 807.000 ;
        RECT 389.400 805.350 390.600 807.000 ;
        RECT 391.950 805.950 394.050 808.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 382.950 802.950 385.050 805.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 380.400 801.900 381.600 802.650 ;
        RECT 386.400 801.900 387.600 802.650 ;
        RECT 379.950 799.800 382.050 801.900 ;
        RECT 385.950 799.800 388.050 801.900 ;
        RECT 373.950 775.950 376.050 778.050 ;
        RECT 379.950 772.950 382.050 775.050 ;
        RECT 368.400 760.350 369.600 762.600 ;
        RECT 364.950 757.950 367.050 760.050 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 365.400 756.900 366.600 757.650 ;
        RECT 371.400 756.900 372.600 757.650 ;
        RECT 364.950 751.950 367.050 756.900 ;
        RECT 370.950 754.800 373.050 756.900 ;
        RECT 367.950 742.950 370.050 745.050 ;
        RECT 361.950 730.950 364.050 733.050 ;
        RECT 347.400 727.350 348.600 728.100 ;
        RECT 353.400 727.350 354.600 729.600 ;
        RECT 358.950 727.950 361.050 730.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 350.400 723.900 351.600 724.650 ;
        RECT 356.400 723.900 357.600 724.650 ;
        RECT 349.950 721.800 352.050 723.900 ;
        RECT 355.950 721.800 358.050 723.900 ;
        RECT 356.400 718.050 357.450 721.800 ;
        RECT 355.950 715.950 358.050 718.050 ;
        RECT 349.950 703.950 352.050 706.050 ;
        RECT 346.950 691.950 349.050 694.050 ;
        RECT 340.950 685.950 343.050 688.050 ;
        RECT 337.950 683.100 340.050 685.200 ;
        RECT 347.400 684.600 348.450 691.950 ;
        RECT 338.400 682.350 339.600 683.100 ;
        RECT 347.400 682.350 348.600 684.600 ;
        RECT 338.100 679.950 340.200 682.050 ;
        RECT 341.400 679.950 343.500 682.050 ;
        RECT 346.800 679.950 348.900 682.050 ;
        RECT 341.400 678.900 342.600 679.650 ;
        RECT 350.400 678.900 351.450 703.950 ;
        RECT 352.950 685.950 355.050 688.050 ;
        RECT 334.950 676.800 337.050 678.900 ;
        RECT 340.950 676.800 343.050 678.900 ;
        RECT 349.950 676.800 352.050 678.900 ;
        RECT 334.950 661.950 337.050 664.050 ;
        RECT 328.950 655.950 331.050 658.050 ;
        RECT 325.950 652.950 328.050 655.050 ;
        RECT 326.400 645.900 327.450 652.950 ;
        RECT 335.400 652.200 336.450 661.950 ;
        RECT 334.950 650.100 337.050 652.200 ;
        RECT 340.950 650.100 343.050 652.200 ;
        RECT 335.400 649.350 336.600 650.100 ;
        RECT 341.400 649.350 342.600 650.100 ;
        RECT 346.950 649.950 349.050 652.050 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 340.950 646.950 343.050 649.050 ;
        RECT 332.400 645.900 333.600 646.650 ;
        RECT 325.950 643.800 328.050 645.900 ;
        RECT 331.950 643.800 334.050 645.900 ;
        RECT 338.400 644.400 339.600 646.650 ;
        RECT 338.400 643.050 339.450 644.400 ;
        RECT 343.950 643.950 346.050 646.050 ;
        RECT 337.950 642.450 340.050 643.050 ;
        RECT 337.950 641.400 342.450 642.450 ;
        RECT 337.950 640.950 340.050 641.400 ;
        RECT 325.950 631.950 328.050 634.050 ;
        RECT 341.400 633.450 342.450 641.400 ;
        RECT 344.400 637.050 345.450 643.950 ;
        RECT 343.950 634.950 346.050 637.050 ;
        RECT 347.400 633.450 348.450 649.950 ;
        RECT 341.400 632.400 348.450 633.450 ;
        RECT 326.400 625.050 327.450 631.950 ;
        RECT 331.950 625.950 334.050 628.050 ;
        RECT 325.950 622.950 328.050 625.050 ;
        RECT 326.400 606.600 327.450 622.950 ;
        RECT 320.400 604.350 321.600 606.600 ;
        RECT 326.400 604.350 327.600 606.600 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 310.950 598.800 313.050 600.900 ;
        RECT 317.400 599.400 318.600 601.650 ;
        RECT 323.400 600.900 324.600 601.650 ;
        RECT 317.400 598.050 318.450 599.400 ;
        RECT 322.950 598.800 325.050 600.900 ;
        RECT 316.950 595.950 319.050 598.050 ;
        RECT 317.400 576.450 318.450 595.950 ;
        RECT 332.400 583.050 333.450 625.950 ;
        RECT 346.950 613.950 349.050 616.050 ;
        RECT 347.400 606.600 348.450 613.950 ;
        RECT 353.400 607.050 354.450 685.950 ;
        RECT 355.950 682.950 358.050 685.050 ;
        RECT 362.400 684.450 363.450 730.950 ;
        RECT 364.950 727.950 367.050 730.050 ;
        RECT 365.400 723.900 366.450 727.950 ;
        RECT 364.950 721.800 367.050 723.900 ;
        RECT 368.400 706.050 369.450 742.950 ;
        RECT 380.400 733.050 381.450 772.950 ;
        RECT 395.400 772.050 396.450 823.950 ;
        RECT 398.400 814.050 399.450 844.950 ;
        RECT 401.400 826.050 402.450 847.950 ;
        RECT 409.950 839.100 412.050 844.050 ;
        RECT 418.950 841.950 421.050 844.050 ;
        RECT 437.400 843.450 438.450 859.950 ;
        RECT 442.950 850.950 445.050 853.050 ;
        RECT 443.400 847.050 444.450 850.950 ;
        RECT 458.400 850.050 459.450 877.800 ;
        RECT 457.950 847.950 460.050 850.050 ;
        RECT 442.950 844.950 445.050 847.050 ;
        RECT 434.400 842.400 438.450 843.450 ;
        RECT 410.400 838.350 411.600 839.100 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 407.400 833.400 408.600 835.650 ;
        RECT 400.950 823.950 403.050 826.050 ;
        RECT 407.400 817.050 408.450 833.400 ;
        RECT 419.400 826.050 420.450 841.950 ;
        RECT 421.950 839.100 424.050 841.200 ;
        RECT 427.950 839.100 430.050 841.200 ;
        RECT 434.400 840.600 435.450 842.400 ;
        RECT 418.950 823.950 421.050 826.050 ;
        RECT 400.950 814.950 403.050 817.050 ;
        RECT 406.950 814.950 409.050 817.050 ;
        RECT 397.950 811.950 400.050 814.050 ;
        RECT 397.950 808.800 400.050 810.900 ;
        RECT 398.400 801.900 399.450 808.800 ;
        RECT 397.950 799.800 400.050 801.900 ;
        RECT 401.400 793.050 402.450 814.950 ;
        RECT 409.950 811.950 412.050 814.050 ;
        RECT 410.400 807.600 411.450 811.950 ;
        RECT 410.400 805.350 411.600 807.600 ;
        RECT 415.950 806.100 418.050 808.200 ;
        RECT 416.400 805.350 417.600 806.100 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 407.400 801.900 408.600 802.650 ;
        RECT 406.950 799.800 409.050 801.900 ;
        RECT 413.400 800.400 414.600 802.650 ;
        RECT 422.400 802.050 423.450 839.100 ;
        RECT 428.400 838.350 429.600 839.100 ;
        RECT 434.400 838.350 435.600 840.600 ;
        RECT 427.950 835.950 430.050 838.050 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 431.400 834.000 432.600 835.650 ;
        RECT 430.950 829.950 433.050 834.000 ;
        RECT 437.400 833.400 438.600 835.650 ;
        RECT 424.950 826.950 427.050 829.050 ;
        RECT 413.400 799.050 414.450 800.400 ;
        RECT 421.950 799.950 424.050 802.050 ;
        RECT 412.950 796.950 415.050 799.050 ;
        RECT 403.950 793.950 406.050 796.050 ;
        RECT 400.950 790.950 403.050 793.050 ;
        RECT 400.950 784.950 403.050 787.050 ;
        RECT 382.950 769.950 385.050 772.050 ;
        RECT 394.950 769.950 397.050 772.050 ;
        RECT 379.950 730.950 382.050 733.050 ;
        RECT 376.950 728.100 379.050 730.200 ;
        RECT 383.400 730.050 384.450 769.950 ;
        RECT 388.950 768.450 391.050 769.050 ;
        RECT 386.400 767.400 391.050 768.450 ;
        RECT 386.400 756.900 387.450 767.400 ;
        RECT 388.950 766.950 391.050 767.400 ;
        RECT 389.400 762.600 390.450 766.950 ;
        RECT 389.400 760.350 390.600 762.600 ;
        RECT 397.950 761.100 400.050 763.200 ;
        RECT 398.400 760.350 399.600 761.100 ;
        RECT 389.100 757.950 391.200 760.050 ;
        RECT 392.400 757.950 394.500 760.050 ;
        RECT 397.800 757.950 399.900 760.050 ;
        RECT 385.950 754.800 388.050 756.900 ;
        RECT 392.400 756.000 393.600 757.650 ;
        RECT 391.950 751.950 394.050 756.000 ;
        RECT 388.950 748.950 391.050 751.050 ;
        RECT 385.950 745.950 388.050 748.050 ;
        RECT 377.400 727.350 378.600 728.100 ;
        RECT 382.950 727.950 385.050 730.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 374.400 722.400 375.600 724.650 ;
        RECT 380.400 723.000 381.600 724.650 ;
        RECT 374.400 715.050 375.450 722.400 ;
        RECT 379.950 718.950 382.050 723.000 ;
        RECT 373.950 712.950 376.050 715.050 ;
        RECT 379.950 712.950 382.050 715.050 ;
        RECT 367.950 703.950 370.050 706.050 ;
        RECT 376.950 691.950 379.050 694.050 ;
        RECT 359.400 683.400 363.450 684.450 ;
        RECT 356.400 652.050 357.450 682.950 ;
        RECT 359.400 652.200 360.450 683.400 ;
        RECT 367.950 683.100 370.050 685.200 ;
        RECT 368.400 682.350 369.600 683.100 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 370.950 679.950 373.050 682.050 ;
        RECT 365.400 678.900 366.600 679.650 ;
        RECT 371.400 678.900 372.600 679.650 ;
        RECT 364.950 676.800 367.050 678.900 ;
        RECT 370.950 676.800 373.050 678.900 ;
        RECT 364.950 664.950 367.050 667.050 ;
        RECT 355.950 649.950 358.050 652.050 ;
        RECT 358.950 650.100 361.050 652.200 ;
        RECT 365.400 651.600 366.450 664.950 ;
        RECT 377.400 654.450 378.450 691.950 ;
        RECT 380.400 667.050 381.450 712.950 ;
        RECT 386.400 684.450 387.450 745.950 ;
        RECT 389.400 742.050 390.450 748.950 ;
        RECT 401.400 745.050 402.450 784.950 ;
        RECT 400.950 742.950 403.050 745.050 ;
        RECT 388.950 739.950 391.050 742.050 ;
        RECT 388.950 727.950 391.050 730.050 ;
        RECT 391.950 727.950 394.050 730.050 ;
        RECT 401.400 729.450 402.600 729.600 ;
        RECT 404.400 729.450 405.450 793.950 ;
        RECT 413.400 793.050 414.450 796.950 ;
        RECT 406.950 790.950 409.050 793.050 ;
        RECT 412.950 790.950 415.050 793.050 ;
        RECT 401.400 728.400 405.450 729.450 ;
        RECT 389.400 712.050 390.450 727.950 ;
        RECT 392.400 715.050 393.450 727.950 ;
        RECT 401.400 727.350 402.600 728.400 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 398.400 722.400 399.600 724.650 ;
        RECT 391.950 712.950 394.050 715.050 ;
        RECT 388.950 709.950 391.050 712.050 ;
        RECT 391.950 703.950 394.050 706.050 ;
        RECT 383.400 683.400 387.450 684.450 ;
        RECT 392.400 684.600 393.450 703.950 ;
        RECT 398.400 688.050 399.450 722.400 ;
        RECT 400.950 718.950 403.050 721.050 ;
        RECT 401.400 712.050 402.450 718.950 ;
        RECT 400.950 709.950 403.050 712.050 ;
        RECT 397.950 685.950 400.050 688.050 ;
        RECT 403.950 685.950 406.050 688.050 ;
        RECT 399.000 684.600 403.050 685.050 ;
        RECT 383.400 678.900 384.450 683.400 ;
        RECT 392.400 682.350 393.600 684.600 ;
        RECT 398.400 682.950 403.050 684.600 ;
        RECT 398.400 682.350 399.600 682.950 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 394.950 679.950 397.050 682.050 ;
        RECT 397.950 679.950 400.050 682.050 ;
        RECT 389.400 678.900 390.600 679.650 ;
        RECT 382.950 676.800 385.050 678.900 ;
        RECT 388.950 676.800 391.050 678.900 ;
        RECT 395.400 677.400 396.600 679.650 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 379.950 658.950 382.050 661.050 ;
        RECT 374.400 653.400 378.450 654.450 ;
        RECT 359.400 649.350 360.600 650.100 ;
        RECT 365.400 649.350 366.600 651.600 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 362.400 644.400 363.600 646.650 ;
        RECT 362.400 607.200 363.450 644.400 ;
        RECT 374.400 628.050 375.450 653.400 ;
        RECT 380.400 652.050 381.450 658.950 ;
        RECT 376.800 649.950 378.900 652.050 ;
        RECT 379.950 649.950 382.050 652.050 ;
        RECT 385.950 650.100 388.050 652.200 ;
        RECT 373.950 625.950 376.050 628.050 ;
        RECT 377.400 622.050 378.450 649.950 ;
        RECT 386.400 649.350 387.600 650.100 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 383.400 645.900 384.600 646.650 ;
        RECT 389.400 645.900 390.600 646.650 ;
        RECT 382.950 643.800 385.050 645.900 ;
        RECT 388.950 643.800 391.050 645.900 ;
        RECT 395.400 625.050 396.450 677.400 ;
        RECT 400.950 652.950 403.050 655.050 ;
        RECT 397.950 649.950 400.050 652.050 ;
        RECT 394.950 622.950 397.050 625.050 ;
        RECT 376.950 619.950 379.050 622.050 ;
        RECT 379.950 613.950 382.050 616.050 ;
        RECT 394.950 613.950 397.050 616.050 ;
        RECT 347.400 604.350 348.600 606.600 ;
        RECT 352.950 604.950 355.050 607.050 ;
        RECT 358.950 604.950 361.050 607.050 ;
        RECT 361.950 605.100 364.050 607.200 ;
        RECT 367.950 605.100 370.050 607.200 ;
        RECT 376.950 606.000 379.050 610.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 344.400 599.400 345.600 601.650 ;
        RECT 350.400 600.900 351.600 601.650 ;
        RECT 359.400 600.900 360.450 604.950 ;
        RECT 368.400 604.350 369.600 605.100 ;
        RECT 377.400 604.350 378.600 606.000 ;
        RECT 368.100 601.950 370.200 604.050 ;
        RECT 373.500 601.950 375.600 604.050 ;
        RECT 376.800 601.950 378.900 604.050 ;
        RECT 374.400 600.900 375.600 601.650 ;
        RECT 380.400 600.900 381.450 613.950 ;
        RECT 382.950 610.950 385.050 613.050 ;
        RECT 344.400 592.050 345.450 599.400 ;
        RECT 349.950 598.800 352.050 600.900 ;
        RECT 358.950 598.800 361.050 600.900 ;
        RECT 373.950 598.800 376.050 600.900 ;
        RECT 379.950 598.800 382.050 600.900 ;
        RECT 343.950 589.950 346.050 592.050 ;
        RECT 361.950 583.950 364.050 586.050 ;
        RECT 331.950 580.950 334.050 583.050 ;
        RECT 314.400 575.400 318.450 576.450 ;
        RECT 314.400 573.600 315.450 575.400 ;
        RECT 321.000 573.600 325.050 574.050 ;
        RECT 314.400 571.350 315.600 573.600 ;
        RECT 320.400 571.950 325.050 573.600 ;
        RECT 331.950 571.950 334.050 574.050 ;
        RECT 340.950 572.100 343.050 574.200 ;
        RECT 320.400 571.350 321.600 571.950 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 319.950 568.950 322.050 571.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 311.400 568.050 312.600 568.650 ;
        RECT 307.950 566.400 312.600 568.050 ;
        RECT 317.400 567.000 318.600 568.650 ;
        RECT 307.950 565.950 312.000 566.400 ;
        RECT 304.950 562.950 307.050 565.050 ;
        RECT 316.950 562.950 319.050 567.000 ;
        RECT 304.950 559.800 307.050 561.900 ;
        RECT 298.950 529.950 301.050 532.050 ;
        RECT 284.400 526.350 285.600 528.000 ;
        RECT 290.400 526.350 291.600 528.600 ;
        RECT 296.400 526.350 297.600 528.600 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 280.950 520.950 283.050 523.050 ;
        RECT 287.400 521.400 288.600 523.650 ;
        RECT 293.400 521.400 294.600 523.650 ;
        RECT 305.400 523.050 306.450 559.800 ;
        RECT 326.400 550.050 327.450 568.950 ;
        RECT 332.400 567.900 333.450 571.950 ;
        RECT 341.400 571.350 342.600 572.100 ;
        RECT 352.800 571.950 354.900 574.050 ;
        RECT 355.950 572.100 358.050 574.200 ;
        RECT 362.400 573.600 363.450 583.950 ;
        RECT 367.950 577.950 370.050 580.050 ;
        RECT 368.400 573.600 369.450 577.950 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 340.950 568.950 343.050 571.050 ;
        RECT 343.950 568.950 346.050 571.050 ;
        RECT 331.950 565.800 334.050 567.900 ;
        RECT 338.400 566.400 339.600 568.650 ;
        RECT 344.400 567.900 345.600 568.650 ;
        RECT 353.400 567.900 354.450 571.950 ;
        RECT 331.950 559.950 334.050 562.050 ;
        RECT 325.950 547.950 328.050 550.050 ;
        RECT 319.950 532.950 322.050 538.050 ;
        RECT 316.950 527.100 319.050 529.200 ;
        RECT 323.400 528.450 324.600 528.600 ;
        RECT 323.400 527.400 330.450 528.450 ;
        RECT 317.400 526.350 318.600 527.100 ;
        RECT 323.400 526.350 324.600 527.400 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 277.950 496.950 280.050 499.050 ;
        RECT 275.400 494.400 279.450 495.450 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 268.950 490.950 271.050 493.050 ;
        RECT 271.950 490.950 274.050 493.050 ;
        RECT 262.950 487.950 265.050 490.050 ;
        RECT 269.400 489.900 270.600 490.650 ;
        RECT 259.950 481.950 262.050 484.050 ;
        RECT 256.950 469.950 259.050 472.050 ;
        RECT 257.400 451.200 258.450 469.950 ;
        RECT 256.950 449.100 259.050 451.200 ;
        RECT 263.400 451.050 264.450 487.950 ;
        RECT 268.950 487.800 271.050 489.900 ;
        RECT 268.950 478.950 271.050 481.050 ;
        RECT 269.400 454.050 270.450 478.950 ;
        RECT 278.400 478.050 279.450 494.400 ;
        RECT 281.400 481.050 282.450 520.950 ;
        RECT 287.400 495.450 288.450 521.400 ;
        RECT 293.400 514.050 294.450 521.400 ;
        RECT 304.950 520.950 307.050 523.050 ;
        RECT 310.950 520.950 313.050 523.050 ;
        RECT 314.400 522.900 315.600 523.650 ;
        RECT 292.950 511.950 295.050 514.050 ;
        RECT 284.400 494.400 288.450 495.450 ;
        RECT 280.950 478.950 283.050 481.050 ;
        RECT 277.950 475.950 280.050 478.050 ;
        RECT 284.400 454.050 285.450 494.400 ;
        RECT 289.950 494.100 292.050 496.200 ;
        RECT 295.950 495.000 298.050 499.050 ;
        RECT 304.950 496.950 307.050 499.050 ;
        RECT 290.400 493.350 291.600 494.100 ;
        RECT 296.400 493.350 297.600 495.000 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 295.950 490.950 298.050 493.050 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 293.400 488.400 294.600 490.650 ;
        RECT 299.400 488.400 300.600 490.650 ;
        RECT 293.400 484.050 294.450 488.400 ;
        RECT 292.950 481.950 295.050 484.050 ;
        RECT 292.950 478.800 295.050 480.900 ;
        RECT 257.400 442.050 258.450 449.100 ;
        RECT 262.950 448.950 265.050 451.050 ;
        RECT 268.950 450.000 271.050 454.050 ;
        RECT 283.950 451.950 286.050 454.050 ;
        RECT 269.400 448.350 270.600 450.000 ;
        RECT 283.950 448.800 286.050 450.900 ;
        RECT 293.400 450.600 294.450 478.800 ;
        RECT 299.400 478.050 300.450 488.400 ;
        RECT 298.950 475.950 301.050 478.050 ;
        RECT 305.400 453.450 306.450 496.950 ;
        RECT 307.950 493.950 310.050 496.050 ;
        RECT 302.400 452.400 306.450 453.450 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 266.400 444.900 267.600 445.650 ;
        RECT 265.950 442.800 268.050 444.900 ;
        RECT 272.400 443.400 273.600 445.650 ;
        RECT 256.950 439.950 259.050 442.050 ;
        RECT 266.400 433.050 267.450 442.800 ;
        RECT 265.950 430.950 268.050 433.050 ;
        RECT 272.400 430.050 273.450 443.400 ;
        RECT 277.950 439.950 280.050 442.050 ;
        RECT 253.950 424.950 256.050 427.050 ;
        RECT 256.950 424.950 259.050 430.050 ;
        RECT 271.950 427.950 274.050 430.050 ;
        RECT 253.950 421.800 256.050 423.900 ;
        RECT 259.950 421.950 262.050 424.050 ;
        RECT 250.950 409.950 253.050 412.050 ;
        RECT 254.400 406.050 255.450 421.800 ;
        RECT 260.400 417.600 261.450 421.950 ;
        RECT 271.950 418.950 274.050 421.050 ;
        RECT 260.400 415.350 261.600 417.600 ;
        RECT 265.950 416.100 268.050 418.200 ;
        RECT 266.400 415.350 267.600 416.100 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 263.400 411.900 264.600 412.650 ;
        RECT 262.950 409.800 265.050 411.900 ;
        RECT 253.950 403.950 256.050 406.050 ;
        RECT 250.950 394.950 253.050 397.050 ;
        RECT 247.950 388.950 250.050 391.050 ;
        RECT 251.400 382.050 252.450 394.950 ;
        RECT 250.950 379.950 253.050 382.050 ;
        RECT 229.950 370.950 232.050 373.050 ;
        RECT 235.950 372.000 238.050 376.050 ;
        RECT 236.400 370.350 237.600 372.000 ;
        RECT 241.950 371.100 244.050 373.200 ;
        RECT 250.950 371.100 253.050 373.200 ;
        RECT 242.400 370.350 243.600 371.100 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 238.950 367.950 241.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 247.950 367.950 250.050 370.050 ;
        RECT 229.950 364.950 232.050 367.050 ;
        RECT 233.400 366.000 234.600 367.650 ;
        RECT 230.400 346.050 231.450 364.950 ;
        RECT 232.950 361.950 235.050 366.000 ;
        RECT 239.400 365.400 240.600 367.650 ;
        RECT 232.950 355.950 235.050 358.050 ;
        RECT 229.950 343.950 232.050 346.050 ;
        RECT 226.950 340.950 229.050 343.050 ;
        RECT 233.400 342.450 234.450 355.950 ;
        RECT 230.400 341.400 234.450 342.450 ;
        RECT 212.400 334.050 213.450 338.400 ;
        RECT 221.400 337.350 222.600 339.600 ;
        RECT 227.400 339.450 228.600 339.600 ;
        RECT 230.400 339.450 231.450 341.400 ;
        RECT 227.400 338.400 231.450 339.450 ;
        RECT 227.400 337.350 228.600 338.400 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 239.400 339.450 240.450 365.400 ;
        RECT 244.950 364.950 247.050 367.050 ;
        RECT 245.400 351.450 246.450 364.950 ;
        RECT 248.400 355.050 249.450 367.950 ;
        RECT 251.400 364.050 252.450 371.100 ;
        RECT 250.950 361.950 253.050 364.050 ;
        RECT 247.950 352.950 250.050 355.050 ;
        RECT 245.400 350.400 249.450 351.450 ;
        RECT 236.400 338.400 240.450 339.450 ;
        RECT 217.950 334.950 220.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 218.400 334.050 219.600 334.650 ;
        RECT 197.400 322.050 198.450 332.400 ;
        RECT 205.950 331.950 208.050 334.050 ;
        RECT 211.950 331.950 214.050 334.050 ;
        RECT 214.950 332.400 219.600 334.050 ;
        RECT 224.400 332.400 225.600 334.650 ;
        RECT 214.950 331.950 219.000 332.400 ;
        RECT 217.950 328.950 220.050 331.050 ;
        RECT 214.950 325.950 217.050 328.050 ;
        RECT 196.950 319.950 199.050 322.050 ;
        RECT 196.950 313.950 199.050 316.050 ;
        RECT 193.950 283.950 196.050 286.050 ;
        RECT 190.950 262.950 193.050 265.050 ;
        RECT 176.400 259.350 177.600 261.600 ;
        RECT 181.950 260.100 184.050 262.200 ;
        RECT 187.950 260.100 190.050 262.200 ;
        RECT 194.400 262.050 195.450 283.950 ;
        RECT 197.400 283.050 198.450 313.950 ;
        RECT 205.950 293.100 208.050 295.200 ;
        RECT 206.400 292.350 207.600 293.100 ;
        RECT 211.950 292.950 214.050 298.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 203.400 288.000 204.600 289.650 ;
        RECT 202.950 283.950 205.050 288.000 ;
        RECT 209.400 287.400 210.600 289.650 ;
        RECT 197.400 281.400 202.050 283.050 ;
        RECT 198.000 280.950 202.050 281.400 ;
        RECT 209.400 271.050 210.450 287.400 ;
        RECT 211.950 277.950 214.050 280.050 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 182.400 259.350 183.600 260.100 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 173.400 254.400 174.600 256.650 ;
        RECT 179.400 255.900 180.600 256.650 ;
        RECT 173.400 249.450 174.450 254.400 ;
        RECT 178.950 253.800 181.050 255.900 ;
        RECT 175.950 249.450 178.050 253.050 ;
        RECT 173.400 249.000 178.050 249.450 ;
        RECT 173.400 248.400 177.450 249.000 ;
        RECT 166.950 226.950 169.050 229.050 ;
        RECT 160.950 214.950 163.050 217.050 ;
        RECT 166.950 216.000 169.050 220.050 ;
        RECT 167.400 214.350 168.600 216.000 ;
        RECT 163.950 211.950 166.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 164.400 210.900 165.600 211.650 ;
        RECT 157.950 208.800 160.050 210.900 ;
        RECT 163.950 208.800 166.050 210.900 ;
        RECT 170.400 209.400 171.600 211.650 ;
        RECT 176.400 211.050 177.450 248.400 ;
        RECT 188.400 247.050 189.450 260.100 ;
        RECT 193.950 259.950 196.050 262.050 ;
        RECT 202.950 260.100 205.050 262.200 ;
        RECT 212.400 262.050 213.450 277.950 ;
        RECT 194.400 255.900 195.450 259.950 ;
        RECT 203.400 259.350 204.600 260.100 ;
        RECT 211.950 259.950 214.050 262.050 ;
        RECT 199.950 256.950 202.050 259.050 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 193.950 253.800 196.050 255.900 ;
        RECT 200.400 255.000 201.600 256.650 ;
        RECT 199.950 250.950 202.050 255.000 ;
        RECT 206.400 254.400 207.600 256.650 ;
        RECT 187.950 244.950 190.050 247.050 ;
        RECT 196.950 235.950 199.050 238.050 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 178.950 215.100 181.050 217.200 ;
        RECT 188.400 216.600 189.450 232.950 ;
        RECT 197.400 229.050 198.450 235.950 ;
        RECT 196.950 226.950 199.050 229.050 ;
        RECT 199.950 217.950 202.050 220.050 ;
        RECT 170.400 199.050 171.450 209.400 ;
        RECT 175.950 208.950 178.050 211.050 ;
        RECT 169.950 196.950 172.050 199.050 ;
        RECT 172.950 190.950 175.050 193.050 ;
        RECT 163.950 183.000 166.050 187.050 ;
        RECT 164.400 181.350 165.600 183.000 ;
        RECT 161.100 178.950 163.200 181.050 ;
        RECT 164.400 178.950 166.500 181.050 ;
        RECT 169.800 178.950 171.900 181.050 ;
        RECT 161.400 176.400 162.600 178.650 ;
        RECT 170.400 177.900 171.600 178.650 ;
        RECT 169.950 177.450 172.050 177.900 ;
        RECT 173.400 177.450 174.450 190.950 ;
        RECT 175.950 184.950 178.050 187.050 ;
        RECT 169.950 176.400 174.450 177.450 ;
        RECT 154.950 172.950 157.050 175.050 ;
        RECT 148.950 169.950 151.050 172.050 ;
        RECT 161.400 166.050 162.450 176.400 ;
        RECT 169.950 175.800 172.050 176.400 ;
        RECT 176.400 175.050 177.450 184.950 ;
        RECT 175.950 172.950 178.050 175.050 ;
        RECT 160.950 163.950 163.050 166.050 ;
        RECT 169.950 163.950 172.050 166.050 ;
        RECT 151.800 142.500 153.900 144.600 ;
        RECT 149.100 133.950 151.200 136.050 ;
        RECT 152.100 135.300 153.300 142.500 ;
        RECT 155.400 139.350 156.600 141.600 ;
        RECT 161.400 141.300 163.500 143.400 ;
        RECT 155.100 136.950 157.200 139.050 ;
        RECT 158.100 137.700 160.200 139.800 ;
        RECT 158.100 135.300 159.000 137.700 ;
        RECT 152.100 134.100 159.000 135.300 ;
        RECT 149.400 132.450 150.600 133.650 ;
        RECT 146.400 131.400 150.600 132.450 ;
        RECT 146.400 121.050 147.450 131.400 ;
        RECT 152.100 128.700 153.000 134.100 ;
        RECT 153.900 132.300 156.000 133.200 ;
        RECT 161.700 132.300 162.600 141.300 ;
        RECT 164.400 138.450 165.600 138.600 ;
        RECT 164.400 137.400 168.450 138.450 ;
        RECT 164.400 136.350 165.600 137.400 ;
        RECT 163.800 133.950 165.900 136.050 ;
        RECT 153.900 131.100 162.600 132.300 ;
        RECT 151.800 126.600 153.900 128.700 ;
        RECT 155.100 128.100 157.200 130.200 ;
        RECT 159.000 129.300 161.100 131.100 ;
        RECT 155.400 127.050 156.600 127.800 ;
        RECT 167.400 127.050 168.450 137.400 ;
        RECT 154.950 124.950 157.050 127.050 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 145.950 118.950 148.050 121.050 ;
        RECT 170.400 118.050 171.450 163.950 ;
        RECT 179.400 163.050 180.450 215.100 ;
        RECT 188.400 214.350 189.600 216.600 ;
        RECT 193.950 215.100 196.050 217.200 ;
        RECT 194.400 214.350 195.600 215.100 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 191.400 210.900 192.600 211.650 ;
        RECT 190.950 208.800 193.050 210.900 ;
        RECT 181.950 181.950 184.050 184.050 ;
        RECT 190.950 182.100 193.050 184.200 ;
        RECT 182.400 175.050 183.450 181.950 ;
        RECT 191.400 181.350 192.600 182.100 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 188.400 177.000 189.600 178.650 ;
        RECT 181.950 172.950 184.050 175.050 ;
        RECT 187.950 172.950 190.050 177.000 ;
        RECT 194.400 176.400 195.600 178.650 ;
        RECT 187.950 169.800 190.050 171.900 ;
        RECT 178.950 160.950 181.050 163.050 ;
        RECT 188.400 138.600 189.450 169.800 ;
        RECT 194.400 166.050 195.450 176.400 ;
        RECT 193.950 163.950 196.050 166.050 ;
        RECT 196.950 160.950 199.050 163.050 ;
        RECT 182.400 138.450 183.600 138.600 ;
        RECT 176.400 137.400 183.600 138.450 ;
        RECT 157.950 115.950 160.050 118.050 ;
        RECT 169.950 115.950 172.050 118.050 ;
        RECT 145.950 109.950 148.050 112.050 ;
        RECT 158.400 111.450 159.450 115.950 ;
        RECT 146.400 106.050 147.450 109.950 ;
        RECT 154.800 108.300 156.900 110.400 ;
        RECT 158.400 109.200 159.600 111.450 ;
        RECT 145.950 103.950 148.050 106.050 ;
        RECT 152.400 105.450 153.600 105.600 ;
        RECT 149.400 104.400 153.600 105.450 ;
        RECT 146.400 99.900 147.450 103.950 ;
        RECT 145.950 97.800 148.050 99.900 ;
        RECT 145.950 91.950 148.050 94.050 ;
        RECT 142.950 67.950 145.050 70.050 ;
        RECT 139.950 64.950 142.050 67.050 ;
        RECT 140.400 55.050 141.450 64.950 ;
        RECT 146.400 61.200 147.450 91.950 ;
        RECT 149.400 76.050 150.450 104.400 ;
        RECT 152.400 103.350 153.600 104.400 ;
        RECT 152.100 100.950 154.200 103.050 ;
        RECT 155.100 102.900 156.000 108.300 ;
        RECT 158.100 106.800 160.200 108.900 ;
        RECT 162.000 105.900 164.100 107.700 ;
        RECT 156.900 104.700 165.600 105.900 ;
        RECT 156.900 103.800 159.000 104.700 ;
        RECT 155.100 101.700 162.000 102.900 ;
        RECT 155.100 94.500 156.300 101.700 ;
        RECT 158.100 97.950 160.200 100.050 ;
        RECT 161.100 99.300 162.000 101.700 ;
        RECT 158.400 95.400 159.600 97.650 ;
        RECT 161.100 97.200 163.200 99.300 ;
        RECT 164.700 95.700 165.600 104.700 ;
        RECT 166.800 100.950 168.900 103.050 ;
        RECT 167.400 99.900 168.600 100.650 ;
        RECT 166.950 97.800 169.050 99.900 ;
        RECT 154.800 92.400 156.900 94.500 ;
        RECT 164.400 93.600 166.500 95.700 ;
        RECT 148.950 73.950 151.050 76.050 ;
        RECT 149.400 70.050 150.450 73.950 ;
        RECT 148.950 67.950 151.050 70.050 ;
        RECT 176.400 64.050 177.450 137.400 ;
        RECT 182.400 136.350 183.600 137.400 ;
        RECT 188.400 136.350 189.600 138.600 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 184.950 133.950 187.050 136.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 190.950 133.950 193.050 136.050 ;
        RECT 185.400 132.900 186.600 133.650 ;
        RECT 191.400 132.900 192.600 133.650 ;
        RECT 184.950 130.800 187.050 132.900 ;
        RECT 190.950 130.800 193.050 132.900 ;
        RECT 197.400 118.050 198.450 160.950 ;
        RECT 196.950 115.950 199.050 118.050 ;
        RECT 187.950 104.100 190.050 106.200 ;
        RECT 196.950 104.100 199.050 106.200 ;
        RECT 188.400 103.350 189.600 104.100 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 185.400 99.900 186.600 100.650 ;
        RECT 184.950 97.800 187.050 99.900 ;
        RECT 191.400 98.400 192.600 100.650 ;
        RECT 191.400 97.050 192.450 98.400 ;
        RECT 197.400 97.050 198.450 104.100 ;
        RECT 190.950 94.950 193.050 97.050 ;
        RECT 196.950 94.950 199.050 97.050 ;
        RECT 181.950 67.950 184.050 70.050 ;
        RECT 145.950 59.100 148.050 61.200 ;
        RECT 169.950 60.000 172.050 64.050 ;
        RECT 175.950 61.950 178.050 64.050 ;
        RECT 146.400 58.350 147.600 59.100 ;
        RECT 170.400 58.350 171.600 60.000 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 139.950 52.950 142.050 55.050 ;
        RECT 149.400 54.900 150.600 55.650 ;
        RECT 148.950 52.800 151.050 54.900 ;
        RECT 167.400 54.000 168.600 55.650 ;
        RECT 182.400 54.900 183.450 67.950 ;
        RECT 191.400 60.600 192.450 94.950 ;
        RECT 200.400 82.050 201.450 217.950 ;
        RECT 206.400 205.050 207.450 254.400 ;
        RECT 211.950 229.950 214.050 232.050 ;
        RECT 212.400 216.600 213.450 229.950 ;
        RECT 215.400 220.050 216.450 325.950 ;
        RECT 218.400 271.050 219.450 328.950 ;
        RECT 220.950 325.950 223.050 328.050 ;
        RECT 221.400 316.050 222.450 325.950 ;
        RECT 224.400 322.050 225.450 332.400 ;
        RECT 226.950 328.950 229.050 331.050 ;
        RECT 223.950 319.950 226.050 322.050 ;
        RECT 220.950 313.950 223.050 316.050 ;
        RECT 227.400 310.050 228.450 328.950 ;
        RECT 226.950 307.950 229.050 310.050 ;
        RECT 233.400 301.050 234.450 337.950 ;
        RECT 220.950 298.950 223.050 301.050 ;
        RECT 232.950 298.950 235.050 301.050 ;
        RECT 217.950 268.950 220.050 271.050 ;
        RECT 221.400 261.450 222.450 298.950 ;
        RECT 236.400 298.050 237.450 338.400 ;
        RECT 241.950 338.100 244.050 340.200 ;
        RECT 248.400 339.600 249.450 350.400 ;
        RECT 242.400 337.350 243.600 338.100 ;
        RECT 248.400 337.350 249.600 339.600 ;
        RECT 254.400 339.450 255.450 403.950 ;
        RECT 272.400 403.050 273.450 418.950 ;
        RECT 274.950 416.100 277.050 418.200 ;
        RECT 275.400 412.050 276.450 416.100 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 274.950 403.950 277.050 406.050 ;
        RECT 265.950 400.950 268.050 403.050 ;
        RECT 271.950 400.950 274.050 403.050 ;
        RECT 266.400 379.050 267.450 400.950 ;
        RECT 265.950 376.950 268.050 379.050 ;
        RECT 271.950 376.950 274.050 379.050 ;
        RECT 259.950 371.100 262.050 373.200 ;
        RECT 266.400 372.600 267.450 376.950 ;
        RECT 260.400 370.350 261.600 371.100 ;
        RECT 266.400 370.350 267.600 372.600 ;
        RECT 272.400 370.050 273.450 376.950 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 263.400 365.400 264.600 367.650 ;
        RECT 263.400 349.050 264.450 365.400 ;
        RECT 275.400 364.050 276.450 403.950 ;
        RECT 265.950 361.950 268.050 364.050 ;
        RECT 274.950 361.950 277.050 364.050 ;
        RECT 262.950 346.950 265.050 349.050 ;
        RECT 259.950 343.950 262.050 346.050 ;
        RECT 266.400 345.450 267.450 361.950 ;
        RECT 263.400 344.400 267.450 345.450 ;
        RECT 254.400 338.400 258.450 339.450 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 238.950 331.950 241.050 334.050 ;
        RECT 245.400 333.900 246.600 334.650 ;
        RECT 251.400 333.900 252.600 334.650 ;
        RECT 239.400 319.050 240.450 331.950 ;
        RECT 244.950 331.800 247.050 333.900 ;
        RECT 250.950 331.800 253.050 333.900 ;
        RECT 247.950 325.950 250.050 328.050 ;
        RECT 238.950 316.950 241.050 319.050 ;
        RECT 244.950 307.950 247.050 310.050 ;
        RECT 226.950 294.000 229.050 298.050 ;
        RECT 235.950 295.950 238.050 298.050 ;
        RECT 241.950 295.950 244.050 298.050 ;
        RECT 227.400 292.350 228.600 294.000 ;
        RECT 232.950 293.100 235.050 295.200 ;
        RECT 233.400 292.350 234.600 293.100 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 223.950 286.950 226.050 289.050 ;
        RECT 230.400 287.400 231.600 289.650 ;
        RECT 236.400 287.400 237.600 289.650 ;
        RECT 224.400 283.050 225.450 286.950 ;
        RECT 223.950 280.950 226.050 283.050 ;
        RECT 230.400 277.050 231.450 287.400 ;
        RECT 236.400 286.050 237.450 287.400 ;
        RECT 235.950 283.950 238.050 286.050 ;
        RECT 229.950 274.950 232.050 277.050 ;
        RECT 226.950 268.950 229.050 271.050 ;
        RECT 218.400 260.400 222.450 261.450 ;
        RECT 227.400 261.600 228.450 268.950 ;
        RECT 218.400 223.050 219.450 260.400 ;
        RECT 227.400 259.350 228.600 261.600 ;
        RECT 232.950 259.950 235.050 262.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 224.400 254.400 225.600 256.650 ;
        RECT 230.400 255.900 231.600 256.650 ;
        RECT 224.400 247.050 225.450 254.400 ;
        RECT 229.950 253.800 232.050 255.900 ;
        RECT 236.400 253.050 237.450 283.950 ;
        RECT 238.950 262.950 241.050 265.050 ;
        RECT 229.950 250.650 232.050 252.750 ;
        RECT 235.950 250.950 238.050 253.050 ;
        RECT 223.950 244.950 226.050 247.050 ;
        RECT 217.950 220.950 220.050 223.050 ;
        RECT 226.950 220.950 229.050 223.050 ;
        RECT 214.950 217.950 217.050 220.050 ;
        RECT 212.400 214.350 213.600 216.600 ;
        RECT 221.400 216.450 222.600 216.600 ;
        RECT 221.400 215.400 225.450 216.450 ;
        RECT 221.400 214.350 222.600 215.400 ;
        RECT 212.100 211.950 214.200 214.050 ;
        RECT 215.400 211.950 217.500 214.050 ;
        RECT 220.800 211.950 222.900 214.050 ;
        RECT 215.400 209.400 216.600 211.650 ;
        RECT 205.950 202.950 208.050 205.050 ;
        RECT 211.950 196.950 214.050 199.050 ;
        RECT 212.400 183.600 213.450 196.950 ;
        RECT 215.400 187.050 216.450 209.400 ;
        RECT 224.400 202.050 225.450 215.400 ;
        RECT 223.950 199.950 226.050 202.050 ;
        RECT 214.950 184.950 217.050 187.050 ;
        RECT 212.400 181.350 213.600 183.600 ;
        RECT 217.950 182.100 220.050 184.200 ;
        RECT 218.400 181.350 219.600 182.100 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 215.400 177.900 216.600 178.650 ;
        RECT 214.950 175.800 217.050 177.900 ;
        RECT 221.400 177.000 222.600 178.650 ;
        RECT 220.950 172.950 223.050 177.000 ;
        RECT 223.950 175.950 226.050 178.050 ;
        RECT 224.400 166.050 225.450 175.950 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 223.950 163.950 226.050 166.050 ;
        RECT 212.400 138.600 213.450 163.950 ;
        RECT 212.400 136.350 213.600 138.600 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 202.950 130.800 205.050 132.900 ;
        RECT 209.400 131.400 210.600 133.650 ;
        RECT 215.400 131.400 216.600 133.650 ;
        RECT 203.400 127.050 204.450 130.800 ;
        RECT 209.400 127.050 210.450 131.400 ;
        RECT 202.950 124.950 205.050 127.050 ;
        RECT 208.950 124.950 211.050 127.050 ;
        RECT 199.950 79.950 202.050 82.050 ;
        RECT 199.950 73.950 202.050 76.050 ;
        RECT 200.400 64.050 201.450 73.950 ;
        RECT 203.400 70.050 204.450 124.950 ;
        RECT 215.400 118.050 216.450 131.400 ;
        RECT 217.950 124.950 220.050 127.050 ;
        RECT 214.950 115.950 217.050 118.050 ;
        RECT 211.950 104.100 214.050 106.200 ;
        RECT 218.400 105.600 219.450 124.950 ;
        RECT 212.400 103.350 213.600 104.100 ;
        RECT 218.400 103.350 219.600 105.600 ;
        RECT 223.950 103.950 226.050 106.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 209.400 98.400 210.600 100.650 ;
        RECT 215.400 99.900 216.600 100.650 ;
        RECT 224.400 99.900 225.450 103.950 ;
        RECT 202.950 67.950 205.050 70.050 ;
        RECT 199.950 61.950 202.050 64.050 ;
        RECT 191.400 58.350 192.600 60.600 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 188.400 54.900 189.600 55.650 ;
        RECT 194.400 54.900 195.600 55.650 ;
        RECT 200.400 54.900 201.450 61.950 ;
        RECT 209.400 61.200 210.450 98.400 ;
        RECT 214.950 97.800 217.050 99.900 ;
        RECT 223.950 97.800 226.050 99.900 ;
        RECT 223.950 79.950 226.050 82.050 ;
        RECT 208.950 60.450 211.050 61.200 ;
        RECT 206.400 59.400 211.050 60.450 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 154.950 49.950 157.050 52.050 ;
        RECT 166.950 49.950 169.050 54.000 ;
        RECT 181.950 52.800 184.050 54.900 ;
        RECT 187.950 52.800 190.050 54.900 ;
        RECT 193.950 52.800 196.050 54.900 ;
        RECT 199.950 52.800 202.050 54.900 ;
        RECT 145.950 26.100 148.050 28.200 ;
        RECT 146.400 25.350 147.600 26.100 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 143.400 21.900 144.600 22.650 ;
        RECT 113.400 20.400 117.600 21.450 ;
        RECT 124.950 19.800 127.050 21.900 ;
        RECT 136.950 19.800 139.050 21.900 ;
        RECT 142.950 19.800 145.050 21.900 ;
        RECT 149.400 21.450 150.600 22.650 ;
        RECT 155.400 21.450 156.450 49.950 ;
        RECT 203.400 34.050 204.450 55.950 ;
        RECT 202.950 31.950 205.050 34.050 ;
        RECT 173.400 27.450 174.600 27.600 ;
        RECT 178.950 27.450 181.050 28.050 ;
        RECT 173.400 26.400 181.050 27.450 ;
        RECT 173.400 25.350 174.600 26.400 ;
        RECT 178.950 25.950 181.050 26.400 ;
        RECT 190.950 26.100 193.050 28.200 ;
        RECT 191.400 25.350 192.600 26.100 ;
        RECT 167.100 22.950 169.200 25.050 ;
        RECT 172.500 22.950 174.600 25.050 ;
        RECT 191.400 22.950 193.500 25.050 ;
        RECT 196.800 22.950 198.900 25.050 ;
        RECT 149.400 20.400 156.450 21.450 ;
        RECT 206.400 13.050 207.450 59.400 ;
        RECT 208.950 59.100 211.050 59.400 ;
        RECT 214.950 59.100 217.050 61.200 ;
        RECT 215.400 58.350 216.600 59.100 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 212.400 53.400 213.600 55.650 ;
        RECT 218.400 54.900 219.600 55.650 ;
        RECT 212.400 46.050 213.450 53.400 ;
        RECT 217.950 52.800 220.050 54.900 ;
        RECT 211.950 43.950 214.050 46.050 ;
        RECT 218.400 27.600 219.450 52.800 ;
        RECT 224.400 46.050 225.450 79.950 ;
        RECT 227.400 54.900 228.450 220.950 ;
        RECT 230.400 139.050 231.450 250.650 ;
        RECT 232.950 235.950 235.050 238.050 ;
        RECT 233.400 175.050 234.450 235.950 ;
        RECT 239.400 216.600 240.450 262.950 ;
        RECT 242.400 226.050 243.450 295.950 ;
        RECT 245.400 262.050 246.450 307.950 ;
        RECT 248.400 283.050 249.450 325.950 ;
        RECT 253.950 301.950 256.050 304.050 ;
        RECT 254.400 294.600 255.450 301.950 ;
        RECT 257.400 301.050 258.450 338.400 ;
        RECT 260.400 328.050 261.450 343.950 ;
        RECT 259.950 325.950 262.050 328.050 ;
        RECT 263.400 325.050 264.450 344.400 ;
        RECT 268.950 338.100 271.050 340.200 ;
        RECT 274.950 339.000 277.050 343.050 ;
        RECT 278.400 340.050 279.450 439.950 ;
        RECT 284.400 421.050 285.450 448.800 ;
        RECT 293.400 448.350 294.600 450.600 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 295.950 445.950 298.050 448.050 ;
        RECT 290.400 444.000 291.600 445.650 ;
        RECT 289.950 439.950 292.050 444.000 ;
        RECT 296.400 443.400 297.600 445.650 ;
        RECT 290.400 427.050 291.450 439.950 ;
        RECT 289.950 424.950 292.050 427.050 ;
        RECT 283.950 417.000 286.050 421.050 ;
        RECT 284.400 415.350 285.600 417.000 ;
        RECT 292.950 416.100 295.050 418.200 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 287.400 411.900 288.600 412.650 ;
        RECT 286.950 409.800 289.050 411.900 ;
        RECT 287.400 400.050 288.450 409.800 ;
        RECT 286.950 397.950 289.050 400.050 ;
        RECT 293.400 397.050 294.450 416.100 ;
        RECT 292.950 394.950 295.050 397.050 ;
        RECT 286.950 379.950 289.050 382.050 ;
        RECT 287.400 372.600 288.450 379.950 ;
        RECT 287.400 370.350 288.600 372.600 ;
        RECT 292.950 372.000 295.050 376.050 ;
        RECT 296.400 373.050 297.450 443.400 ;
        RECT 298.950 442.800 301.050 444.900 ;
        RECT 299.400 439.050 300.450 442.800 ;
        RECT 298.950 436.950 301.050 439.050 ;
        RECT 298.950 409.800 301.050 411.900 ;
        RECT 299.400 406.050 300.450 409.800 ;
        RECT 298.950 403.950 301.050 406.050 ;
        RECT 302.400 400.050 303.450 452.400 ;
        RECT 308.400 444.900 309.450 493.950 ;
        RECT 311.400 484.050 312.450 520.950 ;
        RECT 313.950 520.800 316.050 522.900 ;
        RECT 320.400 521.400 321.600 523.650 ;
        RECT 320.400 511.050 321.450 521.400 ;
        RECT 329.400 520.050 330.450 527.400 ;
        RECT 332.400 526.050 333.450 559.950 ;
        RECT 338.400 559.050 339.450 566.400 ;
        RECT 343.950 565.800 346.050 567.900 ;
        RECT 352.950 565.800 355.050 567.900 ;
        RECT 337.950 556.950 340.050 559.050 ;
        RECT 343.950 556.950 346.050 559.050 ;
        RECT 337.950 529.950 340.050 535.050 ;
        RECT 344.400 528.600 345.450 556.950 ;
        RECT 352.950 553.950 355.050 556.050 ;
        RECT 344.400 526.350 345.600 528.600 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 343.950 523.950 346.050 526.050 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 341.400 522.000 342.600 523.650 ;
        RECT 328.950 517.950 331.050 520.050 ;
        RECT 340.950 517.950 343.050 522.000 ;
        RECT 347.400 521.400 348.600 523.650 ;
        RECT 325.950 514.950 328.050 517.050 ;
        RECT 319.950 508.950 322.050 511.050 ;
        RECT 321.000 495.600 325.050 496.050 ;
        RECT 320.400 493.950 325.050 495.600 ;
        RECT 320.400 493.350 321.600 493.950 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 317.400 488.400 318.600 490.650 ;
        RECT 317.400 484.050 318.450 488.400 ;
        RECT 326.400 487.050 327.450 514.950 ;
        RECT 325.950 484.950 328.050 487.050 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 316.950 481.950 319.050 484.050 ;
        RECT 322.950 481.950 325.050 484.050 ;
        RECT 318.000 453.450 322.050 454.050 ;
        RECT 317.400 451.950 322.050 453.450 ;
        RECT 317.400 450.600 318.450 451.950 ;
        RECT 323.400 451.050 324.450 481.950 ;
        RECT 325.950 451.950 328.050 454.050 ;
        RECT 317.400 448.350 318.600 450.600 ;
        RECT 322.950 448.950 325.050 451.050 ;
        RECT 326.400 448.050 327.450 451.950 ;
        RECT 313.950 445.950 316.050 448.050 ;
        RECT 316.950 445.950 319.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 314.400 444.900 315.600 445.650 ;
        RECT 307.950 442.800 310.050 444.900 ;
        RECT 313.950 442.800 316.050 444.900 ;
        RECT 320.400 443.400 321.600 445.650 ;
        RECT 320.400 436.050 321.450 443.400 ;
        RECT 322.950 442.950 325.050 445.050 ;
        RECT 319.950 433.950 322.050 436.050 ;
        RECT 313.950 430.950 316.050 433.050 ;
        RECT 314.400 423.450 315.450 430.950 ;
        RECT 314.400 421.200 315.600 423.450 ;
        RECT 309.900 417.900 312.000 419.700 ;
        RECT 313.800 418.800 315.900 420.900 ;
        RECT 317.100 420.300 319.200 422.400 ;
        RECT 308.400 416.700 317.100 417.900 ;
        RECT 305.100 412.950 307.200 415.050 ;
        RECT 305.400 411.900 306.600 412.650 ;
        RECT 304.950 409.800 307.050 411.900 ;
        RECT 308.400 407.700 309.300 416.700 ;
        RECT 315.000 415.800 317.100 416.700 ;
        RECT 318.000 414.900 318.900 420.300 ;
        RECT 319.950 416.100 322.050 418.200 ;
        RECT 320.400 415.350 321.600 416.100 ;
        RECT 312.000 413.700 318.900 414.900 ;
        RECT 312.000 411.300 312.900 413.700 ;
        RECT 310.800 409.200 312.900 411.300 ;
        RECT 313.800 409.950 315.900 412.050 ;
        RECT 307.500 405.600 309.600 407.700 ;
        RECT 314.400 407.400 315.600 409.650 ;
        RECT 317.700 406.500 318.900 413.700 ;
        RECT 319.800 412.950 321.900 415.050 ;
        RECT 317.100 404.400 319.200 406.500 ;
        RECT 301.950 397.950 304.050 400.050 ;
        RECT 304.950 394.950 307.050 397.050 ;
        RECT 305.400 382.050 306.450 394.950 ;
        RECT 323.400 382.050 324.450 442.950 ;
        RECT 329.400 433.050 330.450 517.950 ;
        RECT 347.400 511.050 348.450 521.400 ;
        RECT 331.950 508.950 334.050 511.050 ;
        RECT 346.950 508.950 349.050 511.050 ;
        RECT 332.400 445.050 333.450 508.950 ;
        RECT 334.950 499.950 337.050 502.050 ;
        RECT 340.950 499.950 343.050 502.050 ;
        RECT 335.400 496.050 336.450 499.950 ;
        RECT 334.950 493.950 337.050 496.050 ;
        RECT 341.400 495.600 342.450 499.950 ;
        RECT 341.400 493.350 342.600 495.600 ;
        RECT 346.950 494.100 349.050 496.200 ;
        RECT 347.400 493.350 348.600 494.100 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 338.400 488.400 339.600 490.650 ;
        RECT 344.400 489.000 345.600 490.650 ;
        RECT 338.400 478.050 339.450 488.400 ;
        RECT 343.950 484.950 346.050 489.000 ;
        RECT 337.950 475.950 340.050 478.050 ;
        RECT 349.950 451.950 352.050 454.050 ;
        RECT 340.950 449.100 343.050 451.200 ;
        RECT 341.400 448.350 342.600 449.100 ;
        RECT 350.400 448.050 351.450 451.950 ;
        RECT 337.950 445.950 340.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 349.950 445.950 352.050 448.050 ;
        RECT 331.950 442.950 334.050 445.050 ;
        RECT 338.400 443.400 339.600 445.650 ;
        RECT 338.400 439.050 339.450 443.400 ;
        RECT 343.950 442.950 346.050 445.050 ;
        RECT 353.400 444.450 354.450 553.950 ;
        RECT 356.400 553.050 357.450 572.100 ;
        RECT 362.400 571.350 363.600 573.600 ;
        RECT 368.400 571.350 369.600 573.600 ;
        RECT 373.950 572.100 376.050 574.200 ;
        RECT 374.400 571.350 375.600 572.100 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 365.400 566.400 366.600 568.650 ;
        RECT 371.400 567.900 372.600 568.650 ;
        RECT 365.400 562.050 366.450 566.400 ;
        RECT 370.950 565.800 373.050 567.900 ;
        RECT 364.950 559.950 367.050 562.050 ;
        RECT 361.950 556.950 364.050 559.050 ;
        RECT 355.950 550.950 358.050 553.050 ;
        RECT 358.950 499.950 361.050 502.050 ;
        RECT 355.950 493.950 358.050 496.050 ;
        RECT 356.400 489.900 357.450 493.950 ;
        RECT 355.950 487.800 358.050 489.900 ;
        RECT 359.400 472.050 360.450 499.950 ;
        RECT 358.950 469.950 361.050 472.050 ;
        RECT 362.400 463.050 363.450 556.950 ;
        RECT 376.950 544.950 379.050 547.050 ;
        RECT 364.950 528.000 367.050 532.050 ;
        RECT 365.400 526.350 366.600 528.000 ;
        RECT 373.950 527.100 376.050 529.200 ;
        RECT 374.400 526.350 375.600 527.100 ;
        RECT 365.100 523.950 367.200 526.050 ;
        RECT 370.500 523.950 372.600 526.050 ;
        RECT 373.800 523.950 375.900 526.050 ;
        RECT 371.400 521.400 372.600 523.650 ;
        RECT 371.400 517.050 372.450 521.400 ;
        RECT 370.950 514.950 373.050 517.050 ;
        RECT 367.950 494.100 370.050 496.200 ;
        RECT 368.400 493.350 369.600 494.100 ;
        RECT 365.100 490.950 367.200 493.050 ;
        RECT 368.400 490.950 370.500 493.050 ;
        RECT 373.800 490.950 375.900 493.050 ;
        RECT 365.400 489.900 366.600 490.650 ;
        RECT 364.950 487.800 367.050 489.900 ;
        RECT 374.400 488.400 375.600 490.650 ;
        RECT 370.950 484.950 373.050 487.050 ;
        RECT 361.950 460.950 364.050 463.050 ;
        RECT 358.950 450.000 361.050 454.050 ;
        RECT 359.400 448.350 360.600 450.000 ;
        RECT 364.950 449.100 367.050 451.200 ;
        RECT 365.400 448.350 366.600 449.100 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 361.950 445.950 364.050 448.050 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 362.400 444.900 363.600 445.650 ;
        RECT 371.400 445.050 372.450 484.950 ;
        RECT 374.400 463.050 375.450 488.400 ;
        RECT 373.950 460.950 376.050 463.050 ;
        RECT 373.950 454.950 376.050 457.050 ;
        RECT 353.400 443.400 357.450 444.450 ;
        RECT 337.950 436.950 340.050 439.050 ;
        RECT 328.950 430.950 331.050 433.050 ;
        RECT 334.950 424.950 337.050 427.050 ;
        RECT 325.950 418.950 328.050 424.050 ;
        RECT 331.950 415.950 334.050 421.050 ;
        RECT 335.400 417.450 336.450 424.950 ;
        RECT 344.400 423.450 345.450 442.950 ;
        RECT 340.800 420.300 342.900 422.400 ;
        RECT 344.400 421.200 345.600 423.450 ;
        RECT 338.400 417.450 339.600 417.600 ;
        RECT 335.400 416.400 339.600 417.450 ;
        RECT 338.400 415.350 339.600 416.400 ;
        RECT 338.100 412.950 340.200 415.050 ;
        RECT 341.100 414.900 342.000 420.300 ;
        RECT 344.100 418.800 346.200 420.900 ;
        RECT 348.000 417.900 350.100 419.700 ;
        RECT 342.900 416.700 351.600 417.900 ;
        RECT 342.900 415.800 345.000 416.700 ;
        RECT 341.100 413.700 348.000 414.900 ;
        RECT 331.950 406.950 334.050 409.050 ;
        RECT 332.400 397.050 333.450 406.950 ;
        RECT 341.100 406.500 342.300 413.700 ;
        RECT 344.100 409.950 346.200 412.050 ;
        RECT 347.100 411.300 348.000 413.700 ;
        RECT 344.400 407.400 345.600 409.650 ;
        RECT 347.100 409.200 349.200 411.300 ;
        RECT 350.700 407.700 351.600 416.700 ;
        RECT 352.800 412.950 354.900 415.050 ;
        RECT 353.400 411.900 354.600 412.650 ;
        RECT 352.950 409.800 355.050 411.900 ;
        RECT 334.950 403.950 337.050 406.050 ;
        RECT 340.800 404.400 342.900 406.500 ;
        RECT 350.400 405.600 352.500 407.700 ;
        RECT 331.950 394.950 334.050 397.050 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 310.950 379.950 313.050 382.050 ;
        RECT 322.950 379.950 325.050 382.050 ;
        RECT 301.950 373.950 304.050 376.050 ;
        RECT 293.400 370.350 294.600 372.000 ;
        RECT 295.950 370.950 298.050 373.050 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 280.950 364.950 283.050 367.050 ;
        RECT 284.400 365.400 285.600 367.650 ;
        RECT 290.400 366.000 291.600 367.650 ;
        RECT 281.400 346.050 282.450 364.950 ;
        RECT 280.950 343.950 283.050 346.050 ;
        RECT 269.400 337.350 270.600 338.100 ;
        RECT 275.400 337.350 276.600 339.000 ;
        RECT 277.950 337.950 280.050 340.050 ;
        RECT 268.950 334.950 271.050 337.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 272.400 332.400 273.600 334.650 ;
        RECT 262.950 322.950 265.050 325.050 ;
        RECT 272.400 301.050 273.450 332.400 ;
        RECT 277.950 331.950 280.050 334.050 ;
        RECT 278.400 310.050 279.450 331.950 ;
        RECT 277.950 307.950 280.050 310.050 ;
        RECT 256.950 298.950 259.050 301.050 ;
        RECT 259.950 298.950 262.050 301.050 ;
        RECT 271.950 298.950 274.050 301.050 ;
        RECT 260.400 294.600 261.450 298.950 ;
        RECT 271.950 295.800 274.050 297.900 ;
        RECT 254.400 292.350 255.600 294.600 ;
        RECT 260.400 292.350 261.600 294.600 ;
        RECT 265.950 293.100 268.050 295.200 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 250.950 286.950 253.050 289.050 ;
        RECT 257.400 288.900 258.600 289.650 ;
        RECT 247.950 280.950 250.050 283.050 ;
        RECT 251.400 262.200 252.450 286.950 ;
        RECT 256.950 286.800 259.050 288.900 ;
        RECT 256.950 280.950 259.050 283.050 ;
        RECT 262.950 282.450 265.050 283.050 ;
        RECT 266.400 282.450 267.450 293.100 ;
        RECT 272.400 289.050 273.450 295.800 ;
        RECT 281.400 294.600 282.450 343.950 ;
        RECT 284.400 340.200 285.450 365.400 ;
        RECT 289.950 361.950 292.050 366.000 ;
        RECT 286.950 349.950 289.050 352.050 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 283.950 338.100 286.050 340.200 ;
        RECT 284.400 333.900 285.450 338.100 ;
        RECT 287.400 334.050 288.450 349.950 ;
        RECT 292.950 343.950 295.050 346.050 ;
        RECT 293.400 339.600 294.450 343.950 ;
        RECT 299.400 339.600 300.450 349.950 ;
        RECT 302.400 349.050 303.450 373.950 ;
        RECT 301.950 346.950 304.050 349.050 ;
        RECT 305.400 343.050 306.450 379.950 ;
        RECT 311.400 372.600 312.450 379.950 ;
        RECT 311.400 370.350 312.600 372.600 ;
        RECT 316.950 372.000 319.050 376.050 ;
        RECT 317.400 370.350 318.600 372.000 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 314.400 366.900 315.600 367.650 ;
        RECT 313.950 364.800 316.050 366.900 ;
        RECT 323.400 361.050 324.450 379.950 ;
        RECT 328.950 371.100 331.050 373.200 ;
        RECT 335.400 372.600 336.450 403.950 ;
        RECT 356.400 402.450 357.450 443.400 ;
        RECT 361.950 442.800 364.050 444.900 ;
        RECT 370.800 442.950 372.900 445.050 ;
        RECT 374.400 444.900 375.450 454.950 ;
        RECT 373.950 442.800 376.050 444.900 ;
        RECT 377.400 444.450 378.450 544.950 ;
        RECT 383.400 531.450 384.450 610.950 ;
        RECT 395.400 606.600 396.450 613.950 ;
        RECT 398.400 613.050 399.450 649.950 ;
        RECT 401.400 616.050 402.450 652.950 ;
        RECT 404.400 652.050 405.450 685.950 ;
        RECT 407.400 655.050 408.450 790.950 ;
        RECT 425.400 787.050 426.450 826.950 ;
        RECT 433.950 811.950 436.050 814.050 ;
        RECT 427.950 806.100 430.050 808.200 ;
        RECT 434.400 807.600 435.450 811.950 ;
        RECT 437.400 810.450 438.450 833.400 ;
        RECT 443.400 832.050 444.450 844.950 ;
        RECT 457.950 839.100 460.050 841.200 ;
        RECT 458.400 838.350 459.600 839.100 ;
        RECT 463.950 838.950 466.050 841.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 455.400 833.400 456.600 835.650 ;
        RECT 461.400 834.900 462.600 835.650 ;
        RECT 442.950 829.950 445.050 832.050 ;
        RECT 455.400 829.050 456.450 833.400 ;
        RECT 460.950 832.800 463.050 834.900 ;
        RECT 463.950 832.950 466.050 835.050 ;
        RECT 454.950 826.950 457.050 829.050 ;
        RECT 445.950 823.950 448.050 826.050 ;
        RECT 437.400 809.400 441.450 810.450 ;
        RECT 440.400 807.600 441.450 809.400 ;
        RECT 424.950 784.950 427.050 787.050 ;
        RECT 428.400 784.050 429.450 806.100 ;
        RECT 434.400 805.350 435.600 807.600 ;
        RECT 440.400 805.350 441.600 807.600 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 430.950 799.950 433.050 802.050 ;
        RECT 437.400 800.400 438.600 802.650 ;
        RECT 427.950 781.950 430.050 784.050 ;
        RECT 409.950 769.950 412.050 772.050 ;
        RECT 410.400 738.450 411.450 769.950 ;
        RECT 418.950 761.100 421.050 763.200 ;
        RECT 424.950 761.100 427.050 763.200 ;
        RECT 419.400 760.350 420.600 761.100 ;
        RECT 425.400 760.350 426.600 761.100 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 418.950 757.950 421.050 760.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 416.400 755.400 417.600 757.650 ;
        RECT 422.400 756.900 423.600 757.650 ;
        RECT 431.400 757.050 432.450 799.950 ;
        RECT 433.950 761.100 436.050 763.200 ;
        RECT 434.400 757.050 435.450 761.100 ;
        RECT 416.400 751.050 417.450 755.400 ;
        RECT 421.950 754.800 424.050 756.900 ;
        RECT 430.800 754.950 432.900 757.050 ;
        RECT 433.950 754.950 436.050 757.050 ;
        RECT 430.950 751.800 433.050 753.900 ;
        RECT 415.950 748.950 418.050 751.050 ;
        RECT 410.400 737.400 414.450 738.450 ;
        RECT 409.950 733.950 412.050 736.050 ;
        RECT 410.400 658.050 411.450 733.950 ;
        RECT 413.400 694.050 414.450 737.400 ;
        RECT 421.950 728.100 424.050 730.200 ;
        RECT 422.400 727.350 423.600 728.100 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 419.400 723.900 420.600 724.650 ;
        RECT 418.950 721.800 421.050 723.900 ;
        RECT 425.400 722.400 426.600 724.650 ;
        RECT 419.400 709.050 420.450 721.800 ;
        RECT 421.950 712.950 424.050 715.050 ;
        RECT 418.950 706.950 421.050 709.050 ;
        RECT 415.950 700.950 418.050 703.050 ;
        RECT 412.950 691.950 415.050 694.050 ;
        RECT 416.400 684.600 417.450 700.950 ;
        RECT 422.400 691.050 423.450 712.950 ;
        RECT 425.400 697.050 426.450 722.400 ;
        RECT 424.950 694.950 427.050 697.050 ;
        RECT 427.950 691.950 430.050 694.050 ;
        RECT 421.950 688.950 424.050 691.050 ;
        RECT 422.400 684.600 423.450 688.950 ;
        RECT 428.400 688.050 429.450 691.950 ;
        RECT 427.950 685.950 430.050 688.050 ;
        RECT 416.400 682.350 417.600 684.600 ;
        RECT 422.400 682.350 423.600 684.600 ;
        RECT 415.950 679.950 418.050 682.050 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 419.400 678.900 420.600 679.650 ;
        RECT 425.400 678.900 426.600 679.650 ;
        RECT 418.950 676.800 421.050 678.900 ;
        RECT 424.950 676.800 427.050 678.900 ;
        RECT 409.950 655.950 412.050 658.050 ;
        RECT 418.950 655.950 421.050 658.050 ;
        RECT 406.950 652.950 409.050 655.050 ;
        RECT 403.950 649.950 406.050 652.050 ;
        RECT 409.950 650.100 412.050 652.200 ;
        RECT 410.400 649.350 411.600 650.100 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 407.400 645.900 408.600 646.650 ;
        RECT 406.950 643.800 409.050 645.900 ;
        RECT 413.400 644.400 414.600 646.650 ;
        RECT 413.400 640.050 414.450 644.400 ;
        RECT 403.950 637.950 406.050 640.050 ;
        RECT 412.950 637.950 415.050 640.050 ;
        RECT 400.950 613.950 403.050 616.050 ;
        RECT 397.950 610.950 400.050 613.050 ;
        RECT 400.950 607.950 403.050 610.050 ;
        RECT 395.400 604.350 396.600 606.600 ;
        RECT 401.400 606.450 402.600 606.600 ;
        RECT 404.400 606.450 405.450 637.950 ;
        RECT 406.950 613.950 409.050 616.050 ;
        RECT 415.950 613.950 418.050 616.050 ;
        RECT 401.400 605.400 405.450 606.450 ;
        RECT 401.400 604.350 402.600 605.400 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 392.400 599.400 393.600 601.650 ;
        RECT 398.400 599.400 399.600 601.650 ;
        RECT 392.400 577.050 393.450 599.400 ;
        RECT 398.400 583.050 399.450 599.400 ;
        RECT 397.950 580.950 400.050 583.050 ;
        RECT 400.950 577.950 403.050 580.050 ;
        RECT 385.950 574.950 388.050 577.050 ;
        RECT 391.950 574.950 394.050 577.050 ;
        RECT 380.400 530.400 384.450 531.450 ;
        RECT 380.400 502.050 381.450 530.400 ;
        RECT 382.950 526.950 385.050 529.050 ;
        RECT 379.950 499.950 382.050 502.050 ;
        RECT 383.400 474.450 384.450 526.950 ;
        RECT 386.400 496.200 387.450 574.950 ;
        RECT 391.950 571.800 394.050 573.900 ;
        RECT 401.400 573.600 402.450 577.950 ;
        RECT 407.400 574.050 408.450 613.950 ;
        RECT 412.950 610.950 415.050 613.050 ;
        RECT 409.950 607.950 412.050 610.050 ;
        RECT 392.400 538.050 393.450 571.800 ;
        RECT 401.400 571.350 402.600 573.600 ;
        RECT 406.950 571.950 409.050 574.050 ;
        RECT 410.400 573.600 411.450 607.950 ;
        RECT 410.400 571.350 411.600 573.600 ;
        RECT 413.400 573.450 414.450 610.950 ;
        RECT 416.400 606.450 417.450 613.950 ;
        RECT 419.400 610.050 420.450 655.950 ;
        RECT 431.400 655.200 432.450 751.800 ;
        RECT 433.950 742.950 436.050 745.050 ;
        RECT 434.400 721.050 435.450 742.950 ;
        RECT 437.400 736.050 438.450 800.400 ;
        RECT 439.950 784.950 442.050 787.050 ;
        RECT 440.400 763.050 441.450 784.950 ;
        RECT 446.400 780.450 447.450 823.950 ;
        RECT 461.400 823.050 462.450 832.800 ;
        RECT 460.950 820.950 463.050 823.050 ;
        RECT 451.950 808.950 454.050 811.050 ;
        RECT 448.950 806.100 451.050 808.200 ;
        RECT 449.400 790.050 450.450 806.100 ;
        RECT 448.950 787.950 451.050 790.050 ;
        RECT 452.400 787.050 453.450 808.950 ;
        RECT 457.950 807.000 460.050 811.050 ;
        RECT 464.400 807.600 465.450 832.950 ;
        RECT 467.400 829.050 468.450 895.950 ;
        RECT 469.950 871.950 472.050 874.050 ;
        RECT 470.400 834.900 471.450 871.950 ;
        RECT 469.950 832.800 472.050 834.900 ;
        RECT 466.950 826.950 469.050 829.050 ;
        RECT 469.950 823.950 472.050 826.050 ;
        RECT 458.400 805.350 459.600 807.000 ;
        RECT 464.400 805.350 465.600 807.600 ;
        RECT 470.400 807.450 471.450 823.950 ;
        RECT 473.400 817.050 474.450 949.950 ;
        RECT 475.950 937.950 478.050 940.050 ;
        RECT 476.400 912.900 477.450 937.950 ;
        RECT 479.400 934.050 480.450 953.400 ;
        RECT 478.950 931.950 481.050 934.050 ;
        RECT 479.400 913.050 480.450 931.950 ;
        RECT 484.950 918.000 487.050 922.050 ;
        RECT 491.400 919.200 492.450 967.950 ;
        RECT 499.950 962.100 502.050 964.200 ;
        RECT 505.950 962.100 508.050 964.200 ;
        RECT 520.950 963.000 523.050 967.050 ;
        RECT 500.400 961.350 501.600 962.100 ;
        RECT 496.950 958.950 499.050 961.050 ;
        RECT 499.950 958.950 502.050 961.050 ;
        RECT 497.400 957.900 498.600 958.650 ;
        RECT 496.950 955.800 499.050 957.900 ;
        RECT 497.400 925.050 498.450 955.800 ;
        RECT 506.400 940.050 507.450 962.100 ;
        RECT 521.400 961.350 522.600 963.000 ;
        RECT 541.950 962.100 544.050 964.200 ;
        RECT 562.950 962.100 565.050 964.200 ;
        RECT 568.950 962.100 571.050 964.200 ;
        RECT 542.400 961.350 543.600 962.100 ;
        RECT 563.400 961.350 564.600 962.100 ;
        RECT 569.400 961.350 570.600 962.100 ;
        RECT 580.950 961.950 583.050 964.050 ;
        RECT 586.950 962.100 589.050 964.200 ;
        RECT 592.950 963.000 595.050 967.050 ;
        RECT 598.950 964.950 601.050 967.050 ;
        RECT 517.950 958.950 520.050 961.050 ;
        RECT 520.950 958.950 523.050 961.050 ;
        RECT 526.950 958.950 529.050 961.050 ;
        RECT 538.950 958.950 541.050 961.050 ;
        RECT 541.950 958.950 544.050 961.050 ;
        RECT 544.950 958.950 547.050 961.050 ;
        RECT 559.950 958.950 562.050 961.050 ;
        RECT 562.950 958.950 565.050 961.050 ;
        RECT 565.950 958.950 568.050 961.050 ;
        RECT 568.950 958.950 571.050 961.050 ;
        RECT 518.400 956.400 519.600 958.650 ;
        RECT 518.400 949.050 519.450 956.400 ;
        RECT 517.950 946.950 520.050 949.050 ;
        RECT 505.950 937.950 508.050 940.050 ;
        RECT 499.950 925.950 502.050 928.050 ;
        RECT 496.950 922.950 499.050 925.050 ;
        RECT 485.400 916.350 486.600 918.000 ;
        RECT 490.950 917.100 493.050 919.200 ;
        RECT 496.950 917.100 499.050 919.200 ;
        RECT 491.400 916.350 492.600 917.100 ;
        RECT 484.950 913.950 487.050 916.050 ;
        RECT 487.950 913.950 490.050 916.050 ;
        RECT 490.950 913.950 493.050 916.050 ;
        RECT 475.800 910.800 477.900 912.900 ;
        RECT 478.950 910.950 481.050 913.050 ;
        RECT 488.400 912.900 489.600 913.650 ;
        RECT 487.950 910.800 490.050 912.900 ;
        RECT 493.950 901.950 496.050 904.050 ;
        RECT 481.950 884.100 484.050 886.200 ;
        RECT 482.400 883.350 483.600 884.100 ;
        RECT 490.950 883.950 493.050 886.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 481.950 880.950 484.050 883.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 479.400 879.900 480.600 880.650 ;
        RECT 478.950 877.800 481.050 879.900 ;
        RECT 485.400 878.400 486.600 880.650 ;
        RECT 485.400 868.050 486.450 878.400 ;
        RECT 484.950 865.950 487.050 868.050 ;
        RECT 491.400 843.450 492.450 883.950 ;
        RECT 494.400 871.050 495.450 901.950 ;
        RECT 497.400 879.450 498.450 917.100 ;
        RECT 500.400 886.050 501.450 925.950 ;
        RECT 511.950 917.100 514.050 919.200 ;
        RECT 512.400 916.350 513.600 917.100 ;
        RECT 508.950 913.950 511.050 916.050 ;
        RECT 511.950 913.950 514.050 916.050 ;
        RECT 514.950 913.950 517.050 916.050 ;
        RECT 509.400 911.400 510.600 913.650 ;
        RECT 515.400 911.400 516.600 913.650 ;
        RECT 509.400 892.050 510.450 911.400 ;
        RECT 508.950 889.950 511.050 892.050 ;
        RECT 515.400 889.050 516.450 911.400 ;
        RECT 527.400 898.050 528.450 958.950 ;
        RECT 539.400 957.900 540.600 958.650 ;
        RECT 538.950 955.800 541.050 957.900 ;
        RECT 545.400 957.000 546.600 958.650 ;
        RECT 544.950 952.950 547.050 957.000 ;
        RECT 560.400 956.400 561.600 958.650 ;
        RECT 566.400 957.900 567.600 958.650 ;
        RECT 560.400 952.050 561.450 956.400 ;
        RECT 565.950 955.800 568.050 957.900 ;
        RECT 581.400 952.050 582.450 961.950 ;
        RECT 587.400 961.350 588.600 962.100 ;
        RECT 593.400 961.350 594.600 963.000 ;
        RECT 586.950 958.950 589.050 961.050 ;
        RECT 589.950 958.950 592.050 961.050 ;
        RECT 592.950 958.950 595.050 961.050 ;
        RECT 590.400 957.900 591.600 958.650 ;
        RECT 589.950 955.800 592.050 957.900 ;
        RECT 599.400 955.050 600.450 964.950 ;
        RECT 604.950 961.950 607.050 964.050 ;
        RECT 613.950 962.100 616.050 964.200 ;
        RECT 620.400 963.600 621.450 967.950 ;
        RECT 559.950 949.950 562.050 952.050 ;
        RECT 580.950 949.950 583.050 952.050 ;
        RECT 595.950 949.950 598.050 955.050 ;
        RECT 598.950 952.950 601.050 955.050 ;
        RECT 595.950 928.950 598.050 931.050 ;
        RECT 583.950 922.950 586.050 925.050 ;
        RECT 532.950 917.100 535.050 919.200 ;
        RECT 538.950 917.100 541.050 919.200 ;
        RECT 547.950 917.100 550.050 919.200 ;
        RECT 533.400 916.350 534.600 917.100 ;
        RECT 539.400 916.350 540.600 917.100 ;
        RECT 532.950 913.950 535.050 916.050 ;
        RECT 535.950 913.950 538.050 916.050 ;
        RECT 538.950 913.950 541.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 536.400 911.400 537.600 913.650 ;
        RECT 542.400 912.900 543.600 913.650 ;
        RECT 526.950 895.950 529.050 898.050 ;
        RECT 499.950 883.950 502.050 886.050 ;
        RECT 502.950 884.100 505.050 886.200 ;
        RECT 508.950 885.000 511.050 888.900 ;
        RECT 514.950 886.950 517.050 889.050 ;
        RECT 503.400 883.350 504.600 884.100 ;
        RECT 509.400 883.350 510.600 885.000 ;
        RECT 511.950 883.950 514.050 886.050 ;
        RECT 502.950 880.950 505.050 883.050 ;
        RECT 505.950 880.950 508.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 506.400 879.900 507.600 880.650 ;
        RECT 497.400 878.400 501.450 879.450 ;
        RECT 493.950 868.950 496.050 871.050 ;
        RECT 488.400 842.400 492.450 843.450 ;
        RECT 481.950 839.100 484.050 841.200 ;
        RECT 488.400 840.600 489.450 842.400 ;
        RECT 482.400 838.350 483.600 839.100 ;
        RECT 488.400 838.350 489.600 840.600 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 487.950 835.950 490.050 838.050 ;
        RECT 490.950 835.950 493.050 838.050 ;
        RECT 475.950 832.950 478.050 835.050 ;
        RECT 479.400 833.400 480.600 835.650 ;
        RECT 485.400 833.400 486.600 835.650 ;
        RECT 491.400 834.900 492.600 835.650 ;
        RECT 476.400 817.050 477.450 832.950 ;
        RECT 479.400 823.050 480.450 833.400 ;
        RECT 485.400 826.050 486.450 833.400 ;
        RECT 490.950 832.800 493.050 834.900 ;
        RECT 496.950 826.950 499.050 829.050 ;
        RECT 484.950 823.950 487.050 826.050 ;
        RECT 478.950 820.950 481.050 823.050 ;
        RECT 484.950 820.800 487.050 822.900 ;
        RECT 472.950 814.950 475.050 817.050 ;
        RECT 475.950 814.950 478.050 817.050 ;
        RECT 478.950 814.950 481.050 817.050 ;
        RECT 470.400 806.400 474.450 807.450 ;
        RECT 457.950 802.950 460.050 805.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 461.400 800.400 462.600 802.650 ;
        RECT 467.400 801.900 468.600 802.650 ;
        RECT 461.400 793.050 462.450 800.400 ;
        RECT 466.950 799.800 469.050 801.900 ;
        RECT 460.950 790.950 463.050 793.050 ;
        RECT 451.950 784.950 454.050 787.050 ;
        RECT 457.950 781.950 460.050 784.050 ;
        RECT 446.400 779.400 450.450 780.450 ;
        RECT 445.950 775.950 448.050 778.050 ;
        RECT 439.950 760.950 442.050 763.050 ;
        RECT 446.400 762.600 447.450 775.950 ;
        RECT 449.400 766.050 450.450 779.400 ;
        RECT 448.950 763.950 451.050 766.050 ;
        RECT 446.400 760.350 447.600 762.600 ;
        RECT 451.950 761.100 454.050 763.200 ;
        RECT 452.400 760.350 453.600 761.100 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 443.400 756.900 444.600 757.650 ;
        RECT 442.950 754.800 445.050 756.900 ;
        RECT 449.400 755.400 450.600 757.650 ;
        RECT 449.400 748.050 450.450 755.400 ;
        RECT 448.950 745.950 451.050 748.050 ;
        RECT 436.950 733.950 439.050 736.050 ;
        RECT 454.950 733.950 457.050 736.050 ;
        RECT 436.950 728.100 439.050 730.200 ;
        RECT 445.950 728.100 448.050 730.200 ;
        RECT 433.950 718.950 436.050 721.050 ;
        RECT 433.950 709.950 436.050 712.050 ;
        RECT 434.400 688.050 435.450 709.950 ;
        RECT 433.950 685.950 436.050 688.050 ;
        RECT 433.950 682.800 436.050 684.900 ;
        RECT 434.400 673.050 435.450 682.800 ;
        RECT 437.400 676.050 438.450 728.100 ;
        RECT 446.400 727.350 447.600 728.100 ;
        RECT 451.950 727.950 454.050 730.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 443.400 723.000 444.600 724.650 ;
        RECT 442.950 718.950 445.050 723.000 ;
        RECT 448.950 706.950 451.050 709.050 ;
        RECT 449.400 703.050 450.450 706.950 ;
        RECT 448.950 700.950 451.050 703.050 ;
        RECT 445.950 683.100 448.050 685.200 ;
        RECT 452.400 685.050 453.450 727.950 ;
        RECT 455.400 709.050 456.450 733.950 ;
        RECT 454.950 706.950 457.050 709.050 ;
        RECT 446.400 682.350 447.600 683.100 ;
        RECT 451.950 682.950 454.050 685.050 ;
        RECT 442.950 679.950 445.050 682.050 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 448.950 679.950 451.050 682.050 ;
        RECT 443.400 678.450 444.600 679.650 ;
        RECT 449.400 678.900 450.600 679.650 ;
        RECT 440.400 677.400 444.600 678.450 ;
        RECT 436.950 673.950 439.050 676.050 ;
        RECT 433.950 670.950 436.050 673.050 ;
        RECT 440.400 658.050 441.450 677.400 ;
        RECT 448.950 676.800 451.050 678.900 ;
        RECT 451.950 676.950 454.050 679.050 ;
        RECT 442.950 673.950 445.050 676.050 ;
        RECT 439.950 655.950 442.050 658.050 ;
        RECT 421.950 652.950 424.050 655.050 ;
        RECT 430.950 653.100 433.050 655.200 ;
        RECT 422.400 613.050 423.450 652.950 ;
        RECT 430.950 649.950 433.050 652.050 ;
        RECT 436.950 650.100 439.050 652.200 ;
        RECT 431.400 649.350 432.600 649.950 ;
        RECT 437.400 649.350 438.600 650.100 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 434.400 644.400 435.600 646.650 ;
        RECT 421.950 610.950 424.050 613.050 ;
        RECT 418.950 607.950 421.050 610.050 ;
        RECT 419.400 606.450 420.600 606.600 ;
        RECT 416.400 605.400 420.600 606.450 ;
        RECT 424.950 606.000 427.050 610.050 ;
        RECT 419.400 604.350 420.600 605.400 ;
        RECT 425.400 604.350 426.600 606.000 ;
        RECT 418.950 601.950 421.050 604.050 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 422.400 600.900 423.600 601.650 ;
        RECT 421.950 598.800 424.050 600.900 ;
        RECT 428.400 599.400 429.600 601.650 ;
        RECT 434.400 600.900 435.450 644.400 ;
        RECT 443.400 640.050 444.450 673.950 ;
        RECT 445.950 664.950 448.050 667.050 ;
        RECT 442.950 637.950 445.050 640.050 ;
        RECT 439.950 619.950 442.050 622.050 ;
        RECT 436.950 607.950 439.050 610.050 ;
        RECT 418.950 589.950 421.050 592.050 ;
        RECT 413.400 572.400 417.450 573.450 ;
        RECT 395.400 568.950 397.500 571.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 403.950 568.950 406.050 571.050 ;
        RECT 410.100 568.950 412.200 571.050 ;
        RECT 395.400 566.400 396.600 568.650 ;
        RECT 404.400 566.400 405.600 568.650 ;
        RECT 395.400 550.050 396.450 566.400 ;
        RECT 404.400 556.050 405.450 566.400 ;
        RECT 403.950 553.950 406.050 556.050 ;
        RECT 416.400 550.050 417.450 572.400 ;
        RECT 394.950 547.950 397.050 550.050 ;
        RECT 415.950 547.950 418.050 550.050 ;
        RECT 406.950 541.950 409.050 544.050 ;
        RECT 391.950 535.950 394.050 538.050 ;
        RECT 400.950 535.950 403.050 538.050 ;
        RECT 394.950 528.000 397.050 532.050 ;
        RECT 401.400 528.600 402.450 535.950 ;
        RECT 395.400 526.350 396.600 528.000 ;
        RECT 401.400 526.350 402.600 528.600 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 397.950 523.950 400.050 526.050 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 392.400 521.400 393.600 523.650 ;
        RECT 398.400 522.000 399.600 523.650 ;
        RECT 407.400 523.050 408.450 541.950 ;
        RECT 419.400 535.050 420.450 589.950 ;
        RECT 428.400 586.050 429.450 599.400 ;
        RECT 433.950 598.800 436.050 600.900 ;
        RECT 437.400 592.050 438.450 607.950 ;
        RECT 440.400 600.900 441.450 619.950 ;
        RECT 446.400 613.050 447.450 664.950 ;
        RECT 452.400 651.450 453.450 676.950 ;
        RECT 455.400 658.050 456.450 706.950 ;
        RECT 458.400 703.050 459.450 781.950 ;
        RECT 473.400 772.050 474.450 806.400 ;
        RECT 472.950 769.950 475.050 772.050 ;
        RECT 460.950 763.950 463.050 766.050 ;
        RECT 461.400 730.050 462.450 763.950 ;
        RECT 469.950 761.100 472.050 763.200 ;
        RECT 470.400 760.350 471.600 761.100 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 473.400 756.900 474.600 757.650 ;
        RECT 472.950 754.800 475.050 756.900 ;
        RECT 479.400 754.050 480.450 814.950 ;
        RECT 485.400 807.600 486.450 820.800 ;
        RECT 485.400 805.350 486.600 807.600 ;
        RECT 490.950 806.100 493.050 808.200 ;
        RECT 491.400 805.350 492.600 806.100 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 488.400 801.900 489.600 802.650 ;
        RECT 487.950 799.800 490.050 801.900 ;
        RECT 497.400 799.050 498.450 826.950 ;
        RECT 500.400 808.050 501.450 878.400 ;
        RECT 505.950 877.800 508.050 879.900 ;
        RECT 511.950 877.950 514.050 880.050 ;
        RECT 515.400 876.450 516.450 886.950 ;
        RECT 517.950 884.100 520.050 889.050 ;
        RECT 523.950 884.100 526.050 886.200 ;
        RECT 529.950 885.000 532.050 889.050 ;
        RECT 518.400 879.450 519.450 884.100 ;
        RECT 524.400 883.350 525.600 884.100 ;
        RECT 530.400 883.350 531.600 885.000 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 529.950 880.950 532.050 883.050 ;
        RECT 518.400 878.400 522.450 879.450 ;
        RECT 512.400 875.400 516.450 876.450 ;
        RECT 512.400 840.600 513.450 875.400 ;
        RECT 512.400 838.350 513.600 840.600 ;
        RECT 508.950 835.950 511.050 838.050 ;
        RECT 511.950 835.950 514.050 838.050 ;
        RECT 514.950 835.950 517.050 838.050 ;
        RECT 509.400 833.400 510.600 835.650 ;
        RECT 515.400 833.400 516.600 835.650 ;
        RECT 502.950 820.950 505.050 823.050 ;
        RECT 499.950 805.950 502.050 808.050 ;
        RECT 496.950 796.950 499.050 799.050 ;
        RECT 500.400 796.050 501.450 805.950 ;
        RECT 499.950 793.950 502.050 796.050 ;
        RECT 487.950 784.950 490.050 787.050 ;
        RECT 484.950 778.950 487.050 781.050 ;
        RECT 481.950 760.950 484.050 763.050 ;
        RECT 472.950 751.650 475.050 753.750 ;
        RECT 478.950 751.950 481.050 754.050 ;
        RECT 460.950 727.950 463.050 730.050 ;
        RECT 466.950 728.100 469.050 730.200 ;
        RECT 473.400 729.600 474.450 751.650 ;
        RECT 482.400 748.050 483.450 760.950 ;
        RECT 481.950 745.950 484.050 748.050 ;
        RECT 467.400 727.350 468.600 728.100 ;
        RECT 473.400 727.350 474.600 729.600 ;
        RECT 478.950 727.950 481.050 730.050 ;
        RECT 485.400 729.450 486.450 778.950 ;
        RECT 488.400 736.050 489.450 784.950 ;
        RECT 499.950 775.950 502.050 778.050 ;
        RECT 500.400 772.050 501.450 775.950 ;
        RECT 503.400 775.050 504.450 820.950 ;
        RECT 509.400 814.050 510.450 833.400 ;
        RECT 515.400 823.050 516.450 833.400 ;
        RECT 514.950 820.950 517.050 823.050 ;
        RECT 508.950 811.950 511.050 814.050 ;
        RECT 505.950 807.600 510.000 808.050 ;
        RECT 505.950 805.950 510.600 807.600 ;
        RECT 514.950 806.100 517.050 808.200 ;
        RECT 509.400 805.350 510.600 805.950 ;
        RECT 515.400 805.350 516.600 806.100 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 512.400 800.400 513.600 802.650 ;
        RECT 508.950 796.950 511.050 799.050 ;
        RECT 502.950 772.950 505.050 775.050 ;
        RECT 499.950 769.950 502.050 772.050 ;
        RECT 490.950 766.950 493.050 769.050 ;
        RECT 491.400 762.600 492.450 766.950 ;
        RECT 500.400 762.600 501.450 769.950 ;
        RECT 491.400 760.350 492.600 762.600 ;
        RECT 500.400 760.350 501.600 762.600 ;
        RECT 491.100 757.950 493.200 760.050 ;
        RECT 496.500 757.950 498.600 760.050 ;
        RECT 499.800 757.950 501.900 760.050 ;
        RECT 497.400 756.900 498.600 757.650 ;
        RECT 496.950 754.800 499.050 756.900 ;
        RECT 487.950 733.950 490.050 736.050 ;
        RECT 497.400 733.050 498.450 754.800 ;
        RECT 505.950 745.950 508.050 748.050 ;
        RECT 496.950 730.950 499.050 733.050 ;
        RECT 482.400 728.400 486.450 729.450 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 460.950 721.800 463.050 723.900 ;
        RECT 464.400 722.400 465.600 724.650 ;
        RECT 470.400 723.900 471.600 724.650 ;
        RECT 461.400 709.050 462.450 721.800 ;
        RECT 464.400 718.050 465.450 722.400 ;
        RECT 469.950 721.800 472.050 723.900 ;
        RECT 479.400 718.050 480.450 727.950 ;
        RECT 463.950 715.950 466.050 718.050 ;
        RECT 478.950 715.950 481.050 718.050 ;
        RECT 460.950 706.950 463.050 709.050 ;
        RECT 457.950 700.950 460.050 703.050 ;
        RECT 457.950 688.950 460.050 691.050 ;
        RECT 458.400 676.050 459.450 688.950 ;
        RECT 457.950 673.950 460.050 676.050 ;
        RECT 461.400 673.050 462.450 706.950 ;
        RECT 482.400 688.050 483.450 728.400 ;
        RECT 493.950 728.100 496.050 730.200 ;
        RECT 494.400 727.350 495.600 728.100 ;
        RECT 502.950 727.950 505.050 730.050 ;
        RECT 484.950 724.950 487.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 485.400 700.050 486.450 724.950 ;
        RECT 491.400 723.900 492.600 724.650 ;
        RECT 490.950 721.800 493.050 723.900 ;
        RECT 497.400 722.400 498.600 724.650 ;
        RECT 491.400 712.050 492.450 721.800 ;
        RECT 497.400 718.050 498.450 722.400 ;
        RECT 503.400 721.050 504.450 727.950 ;
        RECT 506.400 723.900 507.450 745.950 ;
        RECT 505.950 721.800 508.050 723.900 ;
        RECT 502.950 718.950 505.050 721.050 ;
        RECT 496.950 715.950 499.050 718.050 ;
        RECT 505.950 715.950 508.050 718.050 ;
        RECT 490.950 709.950 493.050 712.050 ;
        RECT 502.950 709.950 505.050 712.050 ;
        RECT 484.950 697.950 487.050 700.050 ;
        RECT 481.950 685.950 484.050 688.050 ;
        RECT 466.950 683.100 469.050 685.200 ;
        RECT 472.950 683.100 475.050 685.200 ;
        RECT 467.400 682.350 468.600 683.100 ;
        RECT 473.400 682.350 474.600 683.100 ;
        RECT 481.950 682.800 484.050 684.900 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 472.950 679.950 475.050 682.050 ;
        RECT 475.950 679.950 478.050 682.050 ;
        RECT 470.400 677.400 471.600 679.650 ;
        RECT 476.400 677.400 477.600 679.650 ;
        RECT 482.400 678.450 483.450 682.800 ;
        RECT 479.400 677.400 483.450 678.450 ;
        RECT 470.400 673.050 471.450 677.400 ;
        RECT 476.400 675.450 477.450 677.400 ;
        RECT 473.400 674.400 477.450 675.450 ;
        RECT 460.950 670.950 463.050 673.050 ;
        RECT 469.950 670.950 472.050 673.050 ;
        RECT 461.400 664.050 462.450 670.950 ;
        RECT 460.950 661.950 463.050 664.050 ;
        RECT 466.950 658.950 469.050 661.050 ;
        RECT 454.950 655.950 457.050 658.050 ;
        RECT 449.400 650.400 453.450 651.450 ;
        RECT 449.400 637.050 450.450 650.400 ;
        RECT 457.950 650.100 460.050 652.200 ;
        RECT 458.400 649.350 459.600 650.100 ;
        RECT 454.950 646.950 457.050 649.050 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 455.400 645.000 456.600 646.650 ;
        RECT 461.400 645.900 462.600 646.650 ;
        RECT 467.400 645.900 468.450 658.950 ;
        RECT 469.950 652.950 472.050 655.050 ;
        RECT 454.950 640.950 457.050 645.000 ;
        RECT 460.950 643.800 463.050 645.900 ;
        RECT 466.950 643.800 469.050 645.900 ;
        RECT 470.400 643.050 471.450 652.950 ;
        RECT 473.400 646.050 474.450 674.400 ;
        RECT 479.400 661.050 480.450 677.400 ;
        RECT 485.400 675.450 486.450 697.950 ;
        RECT 503.400 694.050 504.450 709.950 ;
        RECT 506.400 697.050 507.450 715.950 ;
        RECT 505.950 694.950 508.050 697.050 ;
        RECT 502.950 691.950 505.050 694.050 ;
        RECT 487.950 685.950 490.050 688.050 ;
        RECT 502.950 685.950 505.050 688.050 ;
        RECT 482.400 674.400 486.450 675.450 ;
        RECT 478.950 658.950 481.050 661.050 ;
        RECT 482.400 651.600 483.450 674.400 ;
        RECT 482.400 649.350 483.600 651.600 ;
        RECT 488.400 651.450 489.450 685.950 ;
        RECT 493.950 683.100 496.050 685.200 ;
        RECT 494.400 682.350 495.600 683.100 ;
        RECT 493.950 679.950 496.050 682.050 ;
        RECT 496.950 679.950 499.050 682.050 ;
        RECT 497.400 678.000 498.600 679.650 ;
        RECT 496.950 673.950 499.050 678.000 ;
        RECT 503.400 676.050 504.450 685.950 ;
        RECT 506.400 678.900 507.450 694.950 ;
        RECT 505.950 676.800 508.050 678.900 ;
        RECT 502.950 673.950 505.050 676.050 ;
        RECT 509.400 673.050 510.450 796.950 ;
        RECT 512.400 793.050 513.450 800.400 ;
        RECT 521.400 799.050 522.450 878.400 ;
        RECT 527.400 878.400 528.600 880.650 ;
        RECT 527.400 877.050 528.450 878.400 ;
        RECT 527.400 875.400 532.050 877.050 ;
        RECT 528.000 874.950 532.050 875.400 ;
        RECT 536.400 862.050 537.450 911.400 ;
        RECT 541.950 910.800 544.050 912.900 ;
        RECT 548.400 904.050 549.450 917.100 ;
        RECT 553.950 916.950 556.050 919.050 ;
        RECT 562.950 917.100 565.050 919.200 ;
        RECT 584.400 918.600 585.450 922.950 ;
        RECT 547.950 901.950 550.050 904.050 ;
        RECT 554.400 898.050 555.450 916.950 ;
        RECT 563.400 916.350 564.600 917.100 ;
        RECT 584.400 916.350 585.600 918.600 ;
        RECT 589.950 917.100 592.050 919.200 ;
        RECT 590.400 916.350 591.600 917.100 ;
        RECT 559.950 913.950 562.050 916.050 ;
        RECT 562.950 913.950 565.050 916.050 ;
        RECT 565.950 913.950 568.050 916.050 ;
        RECT 583.950 913.950 586.050 916.050 ;
        RECT 586.950 913.950 589.050 916.050 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 556.950 912.450 559.050 912.900 ;
        RECT 560.400 912.450 561.600 913.650 ;
        RECT 566.400 912.900 567.600 913.650 ;
        RECT 587.400 912.900 588.600 913.650 ;
        RECT 556.950 911.400 561.600 912.450 ;
        RECT 556.950 910.800 559.050 911.400 ;
        RECT 565.950 910.800 568.050 912.900 ;
        RECT 586.950 910.800 589.050 912.900 ;
        RECT 592.950 910.950 595.050 913.050 ;
        RECT 538.950 895.950 541.050 898.050 ;
        RECT 553.950 895.950 556.050 898.050 ;
        RECT 535.950 859.950 538.050 862.050 ;
        RECT 539.400 853.050 540.450 895.950 ;
        RECT 550.950 884.100 553.050 886.200 ;
        RECT 557.400 885.600 558.450 910.800 ;
        RECT 589.950 907.950 592.050 910.050 ;
        RECT 551.400 883.350 552.600 884.100 ;
        RECT 557.400 883.350 558.600 885.600 ;
        RECT 577.950 884.100 580.050 886.200 ;
        RECT 578.400 883.350 579.600 884.100 ;
        RECT 547.950 880.950 550.050 883.050 ;
        RECT 550.950 880.950 553.050 883.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 548.400 879.900 549.600 880.650 ;
        RECT 547.950 877.800 550.050 879.900 ;
        RECT 554.400 879.000 555.600 880.650 ;
        RECT 553.950 874.950 556.050 879.000 ;
        RECT 575.400 878.400 576.600 880.650 ;
        RECT 581.400 879.000 582.600 880.650 ;
        RECT 575.400 871.050 576.450 878.400 ;
        RECT 580.950 874.950 583.050 879.000 ;
        RECT 590.400 877.050 591.450 907.950 ;
        RECT 593.400 880.050 594.450 910.950 ;
        RECT 596.400 910.050 597.450 928.950 ;
        RECT 595.950 907.950 598.050 910.050 ;
        RECT 595.950 901.950 598.050 904.050 ;
        RECT 596.400 888.450 597.450 901.950 ;
        RECT 599.400 892.050 600.450 952.950 ;
        RECT 605.400 949.050 606.450 961.950 ;
        RECT 614.400 961.350 615.600 962.100 ;
        RECT 620.400 961.350 621.600 963.600 ;
        RECT 610.950 958.950 613.050 961.050 ;
        RECT 613.950 958.950 616.050 961.050 ;
        RECT 616.950 958.950 619.050 961.050 ;
        RECT 619.950 958.950 622.050 961.050 ;
        RECT 611.400 957.000 612.600 958.650 ;
        RECT 610.950 952.950 613.050 957.000 ;
        RECT 617.400 956.400 618.600 958.650 ;
        RECT 617.400 954.450 618.450 956.400 ;
        RECT 632.400 955.050 633.450 967.950 ;
        RECT 640.950 962.100 643.050 964.200 ;
        RECT 641.400 961.350 642.600 962.100 ;
        RECT 655.950 961.950 658.050 964.050 ;
        RECT 665.400 963.600 666.450 967.950 ;
        RECT 637.950 958.950 640.050 961.050 ;
        RECT 640.950 958.950 643.050 961.050 ;
        RECT 643.950 958.950 646.050 961.050 ;
        RECT 638.400 957.000 639.600 958.650 ;
        RECT 617.400 953.400 621.450 954.450 ;
        RECT 604.950 946.950 607.050 949.050 ;
        RECT 620.400 946.050 621.450 953.400 ;
        RECT 631.950 952.950 634.050 955.050 ;
        RECT 637.950 952.950 640.050 957.000 ;
        RECT 644.400 956.400 645.600 958.650 ;
        RECT 656.400 957.900 657.450 961.950 ;
        RECT 665.400 961.350 666.600 963.600 ;
        RECT 670.950 962.100 673.050 964.200 ;
        RECT 671.400 961.350 672.600 962.100 ;
        RECT 676.950 961.950 679.050 964.050 ;
        RECT 691.950 962.100 694.050 964.200 ;
        RECT 661.950 958.950 664.050 961.050 ;
        RECT 664.950 958.950 667.050 961.050 ;
        RECT 667.950 958.950 670.050 961.050 ;
        RECT 670.950 958.950 673.050 961.050 ;
        RECT 662.400 957.900 663.600 958.650 ;
        RECT 644.400 946.050 645.450 956.400 ;
        RECT 655.950 955.800 658.050 957.900 ;
        RECT 661.950 955.800 664.050 957.900 ;
        RECT 668.400 956.400 669.600 958.650 ;
        RECT 668.400 949.050 669.450 956.400 ;
        RECT 667.950 946.950 670.050 949.050 ;
        RECT 619.950 943.950 622.050 946.050 ;
        RECT 643.950 943.950 646.050 946.050 ;
        RECT 601.950 937.950 604.050 940.050 ;
        RECT 602.400 907.050 603.450 937.950 ;
        RECT 610.950 917.100 613.050 919.200 ;
        RECT 611.400 916.350 612.600 917.100 ;
        RECT 607.950 913.950 610.050 916.050 ;
        RECT 610.950 913.950 613.050 916.050 ;
        RECT 613.950 913.950 616.050 916.050 ;
        RECT 604.950 910.950 607.050 913.050 ;
        RECT 608.400 911.400 609.600 913.650 ;
        RECT 614.400 911.400 615.600 913.650 ;
        RECT 620.400 912.450 621.450 943.950 ;
        RECT 649.950 925.950 652.050 928.050 ;
        RECT 634.950 922.950 637.050 925.050 ;
        RECT 643.950 922.950 646.050 925.050 ;
        RECT 625.950 916.950 628.050 919.050 ;
        RECT 635.400 918.600 636.450 922.950 ;
        RECT 626.400 912.900 627.450 916.950 ;
        RECT 635.400 916.350 636.600 918.600 ;
        RECT 631.950 913.950 634.050 916.050 ;
        RECT 634.950 913.950 637.050 916.050 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 632.400 912.900 633.600 913.650 ;
        RECT 638.400 912.900 639.600 913.650 ;
        RECT 644.400 912.900 645.450 922.950 ;
        RECT 646.950 917.100 649.050 919.200 ;
        RECT 617.400 911.400 621.450 912.450 ;
        RECT 601.950 904.950 604.050 907.050 ;
        RECT 598.950 889.950 601.050 892.050 ;
        RECT 596.400 887.400 600.450 888.450 ;
        RECT 599.400 885.600 600.450 887.400 ;
        RECT 605.400 885.600 606.450 910.950 ;
        RECT 608.400 901.050 609.450 911.400 ;
        RECT 614.400 907.050 615.450 911.400 ;
        RECT 613.950 904.950 616.050 907.050 ;
        RECT 607.950 898.950 610.050 901.050 ;
        RECT 599.400 883.350 600.600 885.600 ;
        RECT 605.400 883.350 606.600 885.600 ;
        RECT 613.950 883.950 616.050 886.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 604.950 880.950 607.050 883.050 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 592.950 877.950 595.050 880.050 ;
        RECT 602.400 879.000 603.600 880.650 ;
        RECT 608.400 879.900 609.600 880.650 ;
        RECT 589.950 874.950 592.050 877.050 ;
        RECT 601.950 874.950 604.050 879.000 ;
        RECT 607.950 877.800 610.050 879.900 ;
        RECT 614.400 877.050 615.450 883.950 ;
        RECT 613.950 874.950 616.050 877.050 ;
        RECT 604.950 871.950 607.050 874.050 ;
        RECT 574.950 868.950 577.050 871.050 ;
        RECT 547.950 862.950 550.050 865.050 ;
        RECT 538.950 850.950 541.050 853.050 ;
        RECT 535.950 839.100 538.050 841.200 ;
        RECT 541.950 839.100 544.050 841.200 ;
        RECT 536.400 838.350 537.600 839.100 ;
        RECT 542.400 838.350 543.600 839.100 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 535.950 835.950 538.050 838.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 533.400 833.400 534.600 835.650 ;
        RECT 539.400 834.900 540.600 835.650 ;
        RECT 533.400 829.050 534.450 833.400 ;
        RECT 538.950 832.800 541.050 834.900 ;
        RECT 544.950 832.950 547.050 835.050 ;
        RECT 532.950 826.950 535.050 829.050 ;
        RECT 545.400 826.050 546.450 832.950 ;
        RECT 544.950 823.950 547.050 826.050 ;
        RECT 541.950 820.950 544.050 823.050 ;
        RECT 526.950 805.950 529.050 808.050 ;
        RECT 535.950 806.100 538.050 808.200 ;
        RECT 542.400 808.050 543.450 820.950 ;
        RECT 527.400 801.900 528.450 805.950 ;
        RECT 536.400 805.350 537.600 806.100 ;
        RECT 541.950 805.950 544.050 808.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 533.400 801.900 534.600 802.650 ;
        RECT 545.400 802.050 546.450 823.950 ;
        RECT 526.950 799.800 529.050 801.900 ;
        RECT 532.950 799.800 535.050 801.900 ;
        RECT 538.950 799.950 541.050 802.050 ;
        RECT 544.950 799.950 547.050 802.050 ;
        RECT 520.950 796.950 523.050 799.050 ;
        RECT 529.950 793.950 532.050 796.050 ;
        RECT 511.950 790.950 514.050 793.050 ;
        RECT 514.950 787.950 517.050 790.050 ;
        RECT 515.400 781.050 516.450 787.950 ;
        RECT 514.950 778.950 517.050 781.050 ;
        RECT 520.950 761.100 523.050 763.200 ;
        RECT 521.400 760.350 522.600 761.100 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 518.400 755.400 519.600 757.650 ;
        RECT 524.400 755.400 525.600 757.650 ;
        RECT 518.400 742.050 519.450 755.400 ;
        RECT 524.400 751.050 525.450 755.400 ;
        RECT 530.400 754.050 531.450 793.950 ;
        RECT 529.950 751.950 532.050 754.050 ;
        RECT 523.950 748.950 526.050 751.050 ;
        RECT 533.400 742.050 534.450 799.800 ;
        RECT 539.400 787.050 540.450 799.950 ;
        RECT 538.950 784.950 541.050 787.050 ;
        RECT 544.950 769.950 547.050 772.050 ;
        RECT 535.950 763.950 538.050 766.050 ;
        RECT 536.400 756.900 537.450 763.950 ;
        RECT 545.400 762.600 546.450 769.950 ;
        RECT 548.400 766.050 549.450 862.950 ;
        RECT 575.400 862.050 576.450 868.950 ;
        RECT 574.950 859.950 577.050 862.050 ;
        RECT 565.950 856.950 568.050 859.050 ;
        RECT 550.950 839.100 553.050 841.200 ;
        RECT 559.950 839.100 562.050 841.200 ;
        RECT 566.400 840.600 567.450 856.950 ;
        RECT 571.950 853.950 574.050 856.050 ;
        RECT 572.400 841.200 573.450 853.950 ;
        RECT 551.400 835.050 552.450 839.100 ;
        RECT 560.400 838.350 561.600 839.100 ;
        RECT 566.400 838.350 567.600 840.600 ;
        RECT 571.950 839.100 574.050 841.200 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 550.950 832.950 553.050 835.050 ;
        RECT 563.400 834.900 564.600 835.650 ;
        RECT 562.950 832.800 565.050 834.900 ;
        RECT 556.950 826.950 559.050 829.050 ;
        RECT 557.400 817.050 558.450 826.950 ;
        RECT 572.400 819.450 573.450 839.100 ;
        RECT 575.400 823.050 576.450 859.950 ;
        RECT 592.950 847.950 595.050 850.050 ;
        RECT 586.950 839.100 589.050 841.200 ;
        RECT 593.400 840.600 594.450 847.950 ;
        RECT 587.400 838.350 588.600 839.100 ;
        RECT 593.400 838.350 594.600 840.600 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 592.950 835.950 595.050 838.050 ;
        RECT 584.400 833.400 585.600 835.650 ;
        RECT 590.400 834.000 591.600 835.650 ;
        RECT 574.950 820.950 577.050 823.050 ;
        RECT 572.400 818.400 576.450 819.450 ;
        RECT 556.950 814.950 559.050 817.050 ;
        RECT 568.950 814.950 571.050 817.050 ;
        RECT 557.400 807.600 558.450 814.950 ;
        RECT 562.950 808.950 565.050 811.050 ;
        RECT 557.400 805.350 558.600 807.600 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 554.400 801.900 555.600 802.650 ;
        RECT 563.400 802.050 564.450 808.950 ;
        RECT 565.950 805.950 568.050 808.050 ;
        RECT 553.950 799.800 556.050 801.900 ;
        RECT 562.950 799.950 565.050 802.050 ;
        RECT 559.950 778.950 562.050 781.050 ;
        RECT 547.950 763.950 550.050 766.050 ;
        RECT 545.400 760.350 546.600 762.600 ;
        RECT 553.950 761.100 556.050 763.200 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 547.950 757.950 550.050 760.050 ;
        RECT 535.950 754.800 538.050 756.900 ;
        RECT 542.400 755.400 543.600 757.650 ;
        RECT 548.400 756.900 549.600 757.650 ;
        RECT 542.400 754.050 543.450 755.400 ;
        RECT 547.950 754.800 550.050 756.900 ;
        RECT 541.950 751.950 544.050 754.050 ;
        RECT 517.950 739.950 520.050 742.050 ;
        RECT 532.950 739.950 535.050 742.050 ;
        RECT 542.400 733.050 543.450 751.950 ;
        RECT 550.950 739.950 553.050 742.050 ;
        RECT 514.950 729.000 517.050 733.050 ;
        RECT 532.950 730.950 535.050 733.050 ;
        RECT 541.950 730.950 544.050 733.050 ;
        RECT 515.400 727.350 516.600 729.000 ;
        RECT 520.950 728.100 523.050 730.200 ;
        RECT 526.950 728.100 529.050 730.200 ;
        RECT 521.400 727.350 522.600 728.100 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 518.400 723.900 519.600 724.650 ;
        RECT 517.950 721.800 520.050 723.900 ;
        RECT 527.400 712.050 528.450 728.100 ;
        RECT 529.950 727.950 532.050 730.050 ;
        RECT 526.950 709.950 529.050 712.050 ;
        RECT 517.950 703.950 520.050 706.050 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 512.400 688.050 513.450 700.950 ;
        RECT 511.950 685.950 514.050 688.050 ;
        RECT 518.400 684.600 519.450 703.950 ;
        RECT 526.950 691.950 529.050 694.050 ;
        RECT 518.400 682.350 519.600 684.600 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 517.950 679.950 520.050 682.050 ;
        RECT 520.950 679.950 523.050 682.050 ;
        RECT 515.400 677.400 516.600 679.650 ;
        RECT 521.400 678.900 522.600 679.650 ;
        RECT 508.950 670.950 511.050 673.050 ;
        RECT 515.400 664.050 516.450 677.400 ;
        RECT 520.950 676.800 523.050 678.900 ;
        RECT 527.400 678.450 528.450 691.950 ;
        RECT 530.400 679.050 531.450 727.950 ;
        RECT 533.400 706.050 534.450 730.950 ;
        RECT 535.950 729.600 540.000 730.050 ;
        RECT 535.950 727.950 540.600 729.600 ;
        RECT 544.950 728.100 547.050 730.200 ;
        RECT 551.400 729.450 552.450 739.950 ;
        RECT 554.400 739.050 555.450 761.100 ;
        RECT 560.400 756.900 561.450 778.950 ;
        RECT 566.400 769.050 567.450 805.950 ;
        RECT 569.400 781.050 570.450 814.950 ;
        RECT 575.400 808.200 576.450 818.400 ;
        RECT 584.400 817.050 585.450 833.400 ;
        RECT 589.950 829.950 592.050 834.000 ;
        RECT 595.950 832.950 598.050 835.050 ;
        RECT 605.400 834.900 606.450 871.950 ;
        RECT 613.950 868.950 616.050 871.050 ;
        RECT 614.400 856.050 615.450 868.950 ;
        RECT 613.950 853.950 616.050 856.050 ;
        RECT 617.400 853.050 618.450 911.400 ;
        RECT 625.950 910.800 628.050 912.900 ;
        RECT 631.950 910.800 634.050 912.900 ;
        RECT 637.950 910.800 640.050 912.900 ;
        RECT 643.950 910.800 646.050 912.900 ;
        RECT 647.400 910.050 648.450 917.100 ;
        RECT 650.400 912.450 651.450 925.950 ;
        RECT 677.400 922.050 678.450 961.950 ;
        RECT 692.400 961.350 693.600 962.100 ;
        RECT 703.950 961.950 706.050 964.050 ;
        RECT 712.950 962.100 715.050 964.200 ;
        RECT 737.400 963.600 738.450 967.950 ;
        RECT 743.400 963.600 744.450 967.950 ;
        RECT 767.400 964.200 768.450 967.950 ;
        RECT 835.950 964.950 838.050 967.050 ;
        RECT 688.950 958.950 691.050 961.050 ;
        RECT 691.950 958.950 694.050 961.050 ;
        RECT 694.950 958.950 697.050 961.050 ;
        RECT 689.400 957.900 690.600 958.650 ;
        RECT 688.950 955.800 691.050 957.900 ;
        RECT 695.400 956.400 696.600 958.650 ;
        RECT 695.400 946.050 696.450 956.400 ;
        RECT 694.950 943.950 697.050 946.050 ;
        RECT 700.950 934.950 703.050 937.050 ;
        RECT 658.950 917.100 661.050 919.200 ;
        RECT 664.950 918.000 667.050 922.050 ;
        RECT 676.950 919.950 679.050 922.050 ;
        RECT 659.400 916.350 660.600 917.100 ;
        RECT 665.400 916.350 666.600 918.000 ;
        RECT 676.950 916.800 679.050 918.900 ;
        RECT 682.950 917.100 685.050 919.200 ;
        RECT 688.950 917.100 691.050 919.200 ;
        RECT 694.950 917.100 697.050 919.200 ;
        RECT 655.950 913.950 658.050 916.050 ;
        RECT 658.950 913.950 661.050 916.050 ;
        RECT 661.950 913.950 664.050 916.050 ;
        RECT 664.950 913.950 667.050 916.050 ;
        RECT 656.400 912.450 657.600 913.650 ;
        RECT 662.400 912.900 663.600 913.650 ;
        RECT 650.400 911.400 657.600 912.450 ;
        RECT 661.950 910.800 664.050 912.900 ;
        RECT 670.950 910.800 673.050 912.900 ;
        RECT 646.950 907.950 649.050 910.050 ;
        RECT 655.950 907.950 658.050 910.050 ;
        RECT 619.950 898.950 622.050 901.050 ;
        RECT 620.400 856.050 621.450 898.950 ;
        RECT 625.950 895.950 628.050 898.050 ;
        RECT 626.400 886.200 627.450 895.950 ;
        RECT 637.950 889.950 640.050 892.050 ;
        RECT 643.950 889.950 646.050 892.050 ;
        RECT 625.950 884.100 628.050 886.200 ;
        RECT 633.000 885.600 637.050 886.050 ;
        RECT 626.400 883.350 627.600 884.100 ;
        RECT 632.400 883.950 637.050 885.600 ;
        RECT 632.400 883.350 633.600 883.950 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 629.400 879.900 630.600 880.650 ;
        RECT 628.950 877.800 631.050 879.900 ;
        RECT 631.950 874.950 634.050 877.050 ;
        RECT 622.950 865.950 625.050 868.050 ;
        RECT 619.950 853.950 622.050 856.050 ;
        RECT 616.950 850.950 619.050 853.050 ;
        RECT 613.950 839.100 616.050 841.200 ;
        RECT 614.400 838.350 615.600 839.100 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 611.400 834.900 612.600 835.650 ;
        RECT 589.950 820.950 592.050 823.050 ;
        RECT 583.950 814.950 586.050 817.050 ;
        RECT 586.950 808.950 589.050 811.050 ;
        RECT 574.950 806.100 577.050 808.200 ;
        RECT 580.950 806.100 583.050 808.200 ;
        RECT 575.400 805.350 576.600 806.100 ;
        RECT 581.400 805.350 582.600 806.100 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 571.950 799.950 574.050 802.050 ;
        RECT 578.400 800.400 579.600 802.650 ;
        RECT 568.950 778.950 571.050 781.050 ;
        RECT 572.400 775.050 573.450 799.950 ;
        RECT 578.400 778.050 579.450 800.400 ;
        RECT 583.950 799.950 586.050 802.050 ;
        RECT 584.400 787.050 585.450 799.950 ;
        RECT 583.950 784.950 586.050 787.050 ;
        RECT 577.950 775.950 580.050 778.050 ;
        RECT 571.950 772.950 574.050 775.050 ;
        RECT 565.950 766.950 568.050 769.050 ;
        RECT 580.950 766.950 583.050 769.050 ;
        RECT 568.950 761.100 571.050 763.200 ;
        RECT 574.950 761.100 577.050 763.200 ;
        RECT 569.400 760.350 570.600 761.100 ;
        RECT 575.400 760.350 576.600 761.100 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 566.400 756.900 567.600 757.650 ;
        RECT 559.950 754.800 562.050 756.900 ;
        RECT 565.950 754.800 568.050 756.900 ;
        RECT 572.400 755.400 573.600 757.650 ;
        RECT 572.400 742.050 573.450 755.400 ;
        RECT 577.950 748.950 580.050 751.050 ;
        RECT 571.950 739.950 574.050 742.050 ;
        RECT 553.950 736.950 556.050 739.050 ;
        RECT 571.950 736.800 574.050 738.900 ;
        RECT 565.950 733.950 568.050 736.050 ;
        RECT 566.400 729.600 567.450 733.950 ;
        RECT 572.400 729.600 573.450 736.800 ;
        RECT 551.400 728.400 555.450 729.450 ;
        RECT 539.400 727.350 540.600 727.950 ;
        RECT 545.400 727.350 546.600 728.100 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 541.950 724.950 544.050 727.050 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 542.400 723.000 543.600 724.650 ;
        RECT 541.950 718.950 544.050 723.000 ;
        RECT 548.400 722.400 549.600 724.650 ;
        RECT 548.400 706.050 549.450 722.400 ;
        RECT 550.950 715.950 553.050 718.050 ;
        RECT 532.950 703.950 535.050 706.050 ;
        RECT 547.950 703.950 550.050 706.050 ;
        RECT 551.400 703.050 552.450 715.950 ;
        RECT 550.950 700.950 553.050 703.050 ;
        RECT 541.950 694.950 544.050 697.050 ;
        RECT 532.950 685.950 535.050 688.050 ;
        RECT 524.400 677.400 528.450 678.450 ;
        RECT 517.950 670.950 520.050 673.050 ;
        RECT 493.950 661.950 496.050 664.050 ;
        RECT 514.950 661.950 517.050 664.050 ;
        RECT 488.400 650.400 492.450 651.450 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 481.950 646.950 484.050 649.050 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 472.950 643.950 475.050 646.050 ;
        RECT 479.400 645.900 480.600 646.650 ;
        RECT 485.400 645.900 486.600 646.650 ;
        RECT 478.950 643.800 481.050 645.900 ;
        RECT 484.950 643.800 487.050 645.900 ;
        RECT 469.950 640.950 472.050 643.050 ;
        RECT 448.950 634.950 451.050 637.050 ;
        RECT 457.950 634.950 460.050 637.050 ;
        RECT 445.950 610.950 448.050 613.050 ;
        RECT 448.950 605.100 451.050 607.200 ;
        RECT 454.950 605.100 457.050 607.200 ;
        RECT 449.400 604.350 450.600 605.100 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 446.400 600.900 447.600 601.650 ;
        RECT 439.950 598.800 442.050 600.900 ;
        RECT 445.950 598.800 448.050 600.900 ;
        RECT 436.950 589.950 439.050 592.050 ;
        RECT 448.950 589.950 451.050 592.050 ;
        RECT 427.950 583.950 430.050 586.050 ;
        RECT 421.950 577.950 424.050 580.050 ;
        RECT 422.400 535.050 423.450 577.950 ;
        RECT 430.950 572.100 433.050 574.200 ;
        RECT 436.950 572.100 439.050 574.200 ;
        RECT 442.950 572.100 445.050 574.200 ;
        RECT 431.400 571.350 432.600 572.100 ;
        RECT 437.400 571.350 438.600 572.100 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 428.400 566.400 429.600 568.650 ;
        RECT 434.400 567.900 435.600 568.650 ;
        RECT 428.400 544.050 429.450 566.400 ;
        RECT 433.950 565.800 436.050 567.900 ;
        RECT 436.950 562.950 439.050 565.050 ;
        RECT 437.400 559.050 438.450 562.950 ;
        RECT 443.400 559.050 444.450 572.100 ;
        RECT 449.400 565.050 450.450 589.950 ;
        RECT 455.400 583.050 456.450 605.100 ;
        RECT 454.950 580.950 457.050 583.050 ;
        RECT 458.400 577.050 459.450 634.950 ;
        RECT 466.950 628.950 469.050 631.050 ;
        RECT 460.950 616.950 463.050 619.050 ;
        RECT 461.400 601.050 462.450 616.950 ;
        RECT 467.400 606.600 468.450 628.950 ;
        RECT 470.400 610.050 471.450 640.950 ;
        RECT 479.400 622.050 480.450 643.800 ;
        RECT 481.950 634.950 484.050 637.050 ;
        RECT 478.950 619.950 481.050 622.050 ;
        RECT 469.950 609.450 472.050 610.050 ;
        RECT 469.950 608.400 474.450 609.450 ;
        RECT 469.950 607.950 472.050 608.400 ;
        RECT 473.400 606.600 474.450 608.400 ;
        RECT 467.400 604.350 468.600 606.600 ;
        RECT 473.400 604.350 474.600 606.600 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 460.950 598.950 463.050 601.050 ;
        RECT 470.400 600.900 471.600 601.650 ;
        RECT 469.950 598.800 472.050 600.900 ;
        RECT 476.400 600.450 477.600 601.650 ;
        RECT 482.400 600.450 483.450 634.950 ;
        RECT 491.400 606.450 492.450 650.400 ;
        RECT 494.400 640.050 495.450 661.950 ;
        RECT 496.950 658.950 499.050 661.050 ;
        RECT 497.400 646.050 498.450 658.950 ;
        RECT 505.950 651.000 508.050 655.050 ;
        RECT 506.400 649.350 507.600 651.000 ;
        RECT 511.950 650.100 514.050 652.200 ;
        RECT 512.400 649.350 513.600 650.100 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 496.950 643.950 499.050 646.050 ;
        RECT 503.400 644.400 504.600 646.650 ;
        RECT 509.400 644.400 510.600 646.650 ;
        RECT 493.950 637.950 496.050 640.050 ;
        RECT 503.400 637.050 504.450 644.400 ;
        RECT 509.400 640.050 510.450 644.400 ;
        RECT 514.950 643.950 517.050 646.050 ;
        RECT 508.950 637.950 511.050 640.050 ;
        RECT 502.950 634.950 505.050 637.050 ;
        RECT 515.400 631.050 516.450 643.950 ;
        RECT 514.950 628.950 517.050 631.050 ;
        RECT 518.400 628.050 519.450 670.950 ;
        RECT 521.400 642.450 522.450 676.800 ;
        RECT 524.400 646.050 525.450 677.400 ;
        RECT 529.950 676.950 532.050 679.050 ;
        RECT 533.400 673.050 534.450 685.950 ;
        RECT 542.400 684.600 543.450 694.950 ;
        RECT 554.400 688.050 555.450 728.400 ;
        RECT 566.400 727.350 567.600 729.600 ;
        RECT 572.400 727.350 573.600 729.600 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 571.950 724.950 574.050 727.050 ;
        RECT 556.950 721.950 559.050 724.050 ;
        RECT 569.400 723.900 570.600 724.650 ;
        RECT 578.400 724.050 579.450 748.950 ;
        RECT 581.400 747.450 582.450 766.950 ;
        RECT 584.400 766.050 585.450 784.950 ;
        RECT 583.950 763.950 586.050 766.050 ;
        RECT 583.950 760.800 586.050 762.900 ;
        RECT 584.400 754.050 585.450 760.800 ;
        RECT 583.950 751.950 586.050 754.050 ;
        RECT 581.400 746.400 585.450 747.450 ;
        RECT 580.950 739.950 583.050 742.050 ;
        RECT 553.950 685.950 556.050 688.050 ;
        RECT 542.400 682.350 543.600 684.600 ;
        RECT 547.950 683.100 550.050 685.200 ;
        RECT 548.400 682.350 549.600 683.100 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 541.950 679.950 544.050 682.050 ;
        RECT 544.950 679.950 547.050 682.050 ;
        RECT 547.950 679.950 550.050 682.050 ;
        RECT 539.400 677.400 540.600 679.650 ;
        RECT 545.400 678.000 546.600 679.650 ;
        RECT 532.950 670.950 535.050 673.050 ;
        RECT 529.950 650.100 532.050 652.200 ;
        RECT 535.950 651.000 538.050 655.050 ;
        RECT 539.400 652.050 540.450 677.400 ;
        RECT 544.950 673.950 547.050 678.000 ;
        RECT 557.400 676.050 558.450 721.950 ;
        RECT 568.950 721.800 571.050 723.900 ;
        RECT 577.950 721.950 580.050 724.050 ;
        RECT 559.950 709.950 562.050 712.050 ;
        RECT 560.400 678.900 561.450 709.950 ;
        RECT 581.400 697.050 582.450 739.950 ;
        RECT 584.400 723.900 585.450 746.400 ;
        RECT 587.400 736.050 588.450 808.950 ;
        RECT 590.400 772.050 591.450 820.950 ;
        RECT 592.950 814.950 595.050 817.050 ;
        RECT 593.400 790.050 594.450 814.950 ;
        RECT 596.400 808.050 597.450 832.950 ;
        RECT 604.950 832.800 607.050 834.900 ;
        RECT 610.950 832.800 613.050 834.900 ;
        RECT 617.400 834.000 618.600 835.650 ;
        RECT 601.950 829.950 604.050 832.050 ;
        RECT 616.950 831.450 619.050 834.000 ;
        RECT 616.950 830.400 621.450 831.450 ;
        RECT 616.950 829.950 619.050 830.400 ;
        RECT 598.950 823.950 601.050 826.050 ;
        RECT 599.400 811.050 600.450 823.950 ;
        RECT 602.400 814.050 603.450 829.950 ;
        RECT 604.950 826.950 607.050 829.050 ;
        RECT 601.950 811.950 604.050 814.050 ;
        RECT 598.950 808.950 601.050 811.050 ;
        RECT 595.950 805.950 598.050 808.050 ;
        RECT 602.400 807.600 603.450 811.950 ;
        RECT 605.400 811.050 606.450 826.950 ;
        RECT 613.950 820.950 616.050 823.050 ;
        RECT 604.950 808.950 607.050 811.050 ;
        RECT 614.400 808.050 615.450 820.950 ;
        RECT 602.400 805.350 603.600 807.600 ;
        RECT 613.950 805.950 616.050 808.050 ;
        RECT 620.400 807.450 621.450 830.400 ;
        RECT 623.400 823.050 624.450 865.950 ;
        RECT 632.400 865.050 633.450 874.950 ;
        RECT 638.400 865.050 639.450 889.950 ;
        RECT 640.950 883.950 643.050 886.050 ;
        RECT 641.400 871.050 642.450 883.950 ;
        RECT 640.950 868.950 643.050 871.050 ;
        RECT 631.950 862.950 634.050 865.050 ;
        RECT 637.950 862.950 640.050 865.050 ;
        RECT 644.400 859.050 645.450 889.950 ;
        RECT 649.950 884.100 652.050 886.200 ;
        RECT 656.400 885.600 657.450 907.950 ;
        RECT 667.950 901.950 670.050 904.050 ;
        RECT 650.400 883.350 651.600 884.100 ;
        RECT 656.400 883.350 657.600 885.600 ;
        RECT 661.950 884.100 664.050 886.200 ;
        RECT 662.400 883.350 663.600 884.100 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 652.950 880.950 655.050 883.050 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 646.950 877.950 649.050 880.050 ;
        RECT 653.400 879.900 654.600 880.650 ;
        RECT 659.400 879.900 660.600 880.650 ;
        RECT 668.400 879.900 669.450 901.950 ;
        RECT 671.400 886.200 672.450 910.800 ;
        RECT 677.400 904.050 678.450 916.800 ;
        RECT 683.400 916.350 684.600 917.100 ;
        RECT 689.400 916.350 690.600 917.100 ;
        RECT 695.400 916.350 696.600 917.100 ;
        RECT 682.950 913.950 685.050 916.050 ;
        RECT 685.950 913.950 688.050 916.050 ;
        RECT 688.950 913.950 691.050 916.050 ;
        RECT 691.950 913.950 694.050 916.050 ;
        RECT 694.950 913.950 697.050 916.050 ;
        RECT 686.400 912.900 687.600 913.650 ;
        RECT 685.950 910.800 688.050 912.900 ;
        RECT 692.400 912.000 693.600 913.650 ;
        RECT 691.950 907.950 694.050 912.000 ;
        RECT 701.400 910.050 702.450 934.950 ;
        RECT 704.400 919.200 705.450 961.950 ;
        RECT 713.400 961.350 714.600 962.100 ;
        RECT 737.400 961.350 738.600 963.600 ;
        RECT 743.400 961.350 744.600 963.600 ;
        RECT 748.950 962.100 751.050 964.200 ;
        RECT 760.950 962.100 763.050 964.200 ;
        RECT 766.950 962.100 769.050 964.200 ;
        RECT 772.950 962.100 775.050 964.200 ;
        RECT 778.950 962.100 781.050 964.200 ;
        RECT 787.950 962.100 790.050 964.200 ;
        RECT 793.950 962.100 796.050 964.200 ;
        RECT 817.950 962.100 820.050 964.200 ;
        RECT 712.950 958.950 715.050 961.050 ;
        RECT 715.950 958.950 718.050 961.050 ;
        RECT 733.950 958.950 736.050 961.050 ;
        RECT 736.950 958.950 739.050 961.050 ;
        RECT 739.950 958.950 742.050 961.050 ;
        RECT 742.950 958.950 745.050 961.050 ;
        RECT 716.400 956.400 717.600 958.650 ;
        RECT 734.400 957.450 735.600 958.650 ;
        RECT 731.400 956.400 735.600 957.450 ;
        RECT 740.400 957.000 741.600 958.650 ;
        RECT 716.400 943.050 717.450 956.400 ;
        RECT 715.950 940.950 718.050 943.050 ;
        RECT 716.400 928.050 717.450 940.950 ;
        RECT 721.950 931.950 724.050 934.050 ;
        RECT 727.950 931.950 730.050 934.050 ;
        RECT 706.950 925.950 709.050 928.050 ;
        RECT 715.950 925.950 718.050 928.050 ;
        RECT 703.950 917.100 706.050 919.200 ;
        RECT 700.950 907.950 703.050 910.050 ;
        RECT 676.950 901.950 679.050 904.050 ;
        RECT 704.400 903.450 705.450 917.100 ;
        RECT 701.400 902.400 705.450 903.450 ;
        RECT 701.400 898.050 702.450 902.400 ;
        RECT 703.950 898.950 706.050 901.050 ;
        RECT 673.950 895.950 676.050 898.050 ;
        RECT 679.950 895.950 682.050 898.050 ;
        RECT 700.950 897.450 703.050 898.050 ;
        RECT 698.400 896.400 703.050 897.450 ;
        RECT 670.950 884.100 673.050 886.200 ;
        RECT 647.400 874.050 648.450 877.950 ;
        RECT 652.950 877.800 655.050 879.900 ;
        RECT 658.950 877.800 661.050 879.900 ;
        RECT 667.950 877.800 670.050 879.900 ;
        RECT 646.800 871.950 648.900 874.050 ;
        RECT 649.950 871.950 652.050 877.050 ;
        RECT 671.400 862.050 672.450 884.100 ;
        RECT 674.400 880.050 675.450 895.950 ;
        RECT 680.400 885.600 681.450 895.950 ;
        RECT 680.400 883.350 681.600 885.600 ;
        RECT 685.950 885.000 688.050 889.050 ;
        RECT 691.950 886.950 694.050 892.050 ;
        RECT 694.950 889.950 697.050 892.050 ;
        RECT 686.400 883.350 687.600 885.000 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 673.950 877.950 676.050 880.050 ;
        RECT 683.400 879.900 684.600 880.650 ;
        RECT 682.950 877.800 685.050 879.900 ;
        RECT 685.950 874.950 688.050 877.050 ;
        RECT 679.950 865.950 682.050 868.050 ;
        RECT 670.950 859.950 673.050 862.050 ;
        RECT 643.950 856.950 646.050 859.050 ;
        RECT 628.950 853.950 631.050 856.050 ;
        RECT 629.400 847.050 630.450 853.950 ;
        RECT 661.950 850.950 664.050 853.050 ;
        RECT 646.950 847.950 649.050 850.050 ;
        RECT 628.950 844.950 631.050 847.050 ;
        RECT 625.950 841.950 628.050 844.050 ;
        RECT 626.400 832.050 627.450 841.950 ;
        RECT 628.950 838.950 631.050 841.050 ;
        RECT 637.950 839.100 640.050 841.200 ;
        RECT 629.400 834.900 630.450 838.950 ;
        RECT 638.400 838.350 639.600 839.100 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 635.400 834.900 636.600 835.650 ;
        RECT 641.400 834.900 642.600 835.650 ;
        RECT 647.400 834.900 648.450 847.950 ;
        RECT 662.400 844.200 663.450 850.950 ;
        RECT 661.950 842.100 664.050 844.200 ;
        RECT 661.950 838.950 664.050 841.050 ;
        RECT 667.950 839.100 670.050 841.200 ;
        RECT 673.950 839.100 676.050 841.200 ;
        RECT 662.400 838.350 663.600 838.950 ;
        RECT 668.400 838.350 669.600 839.100 ;
        RECT 658.950 835.950 661.050 838.050 ;
        RECT 661.950 835.950 664.050 838.050 ;
        RECT 664.950 835.950 667.050 838.050 ;
        RECT 667.950 835.950 670.050 838.050 ;
        RECT 628.950 832.800 631.050 834.900 ;
        RECT 634.950 832.800 637.050 834.900 ;
        RECT 640.950 832.800 643.050 834.900 ;
        RECT 646.950 832.800 649.050 834.900 ;
        RECT 659.400 833.400 660.600 835.650 ;
        RECT 665.400 834.900 666.600 835.650 ;
        RECT 625.950 829.950 628.050 832.050 ;
        RECT 659.400 826.050 660.450 833.400 ;
        RECT 664.950 832.800 667.050 834.900 ;
        RECT 669.000 828.450 673.050 829.050 ;
        RECT 668.400 826.950 673.050 828.450 ;
        RECT 658.950 823.950 661.050 826.050 ;
        RECT 622.950 820.950 625.050 823.050 ;
        RECT 637.950 820.950 640.050 823.050 ;
        RECT 622.950 814.950 625.050 817.050 ;
        RECT 628.950 814.950 631.050 817.050 ;
        RECT 617.400 806.400 621.450 807.450 ;
        RECT 623.400 807.600 624.450 814.950 ;
        RECT 629.400 807.600 630.450 814.950 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 599.400 801.900 600.600 802.650 ;
        RECT 605.400 801.900 606.600 802.650 ;
        RECT 617.400 801.900 618.450 806.400 ;
        RECT 623.400 805.350 624.600 807.600 ;
        RECT 629.400 805.350 630.600 807.600 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 598.950 799.800 601.050 801.900 ;
        RECT 604.950 799.800 607.050 801.900 ;
        RECT 616.950 799.800 619.050 801.900 ;
        RECT 626.400 800.400 627.600 802.650 ;
        RECT 632.400 800.400 633.600 802.650 ;
        RECT 592.950 787.950 595.050 790.050 ;
        RECT 601.950 781.950 604.050 784.050 ;
        RECT 595.950 775.950 598.050 778.050 ;
        RECT 589.950 769.950 592.050 772.050 ;
        RECT 589.950 760.950 592.050 766.050 ;
        RECT 596.400 763.200 597.450 775.950 ;
        RECT 595.950 761.100 598.050 763.200 ;
        RECT 602.400 762.600 603.450 781.950 ;
        RECT 626.400 778.050 627.450 800.400 ;
        RECT 632.400 796.050 633.450 800.400 ;
        RECT 631.950 793.950 634.050 796.050 ;
        RECT 634.950 781.950 637.050 784.050 ;
        RECT 625.950 775.950 628.050 778.050 ;
        RECT 631.950 775.950 634.050 778.050 ;
        RECT 607.950 772.950 610.050 775.050 ;
        RECT 596.400 760.350 597.600 761.100 ;
        RECT 602.400 760.350 603.600 762.600 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 593.400 756.000 594.600 757.650 ;
        RECT 592.950 751.950 595.050 756.000 ;
        RECT 599.400 755.400 600.600 757.650 ;
        RECT 599.400 751.050 600.450 755.400 ;
        RECT 604.950 754.950 607.050 757.050 ;
        RECT 601.950 751.950 604.050 754.050 ;
        RECT 592.950 748.800 595.050 750.900 ;
        RECT 598.950 748.950 601.050 751.050 ;
        RECT 586.950 733.950 589.050 736.050 ;
        RECT 593.400 729.600 594.450 748.800 ;
        RECT 602.400 748.050 603.450 751.950 ;
        RECT 601.950 745.950 604.050 748.050 ;
        RECT 601.950 739.950 604.050 742.050 ;
        RECT 602.400 730.050 603.450 739.950 ;
        RECT 593.400 727.350 594.600 729.600 ;
        RECT 601.950 727.950 604.050 730.050 ;
        RECT 589.950 724.950 592.050 727.050 ;
        RECT 592.950 724.950 595.050 727.050 ;
        RECT 595.950 724.950 598.050 727.050 ;
        RECT 583.950 721.800 586.050 723.900 ;
        RECT 586.950 721.950 589.050 724.050 ;
        RECT 590.400 723.900 591.600 724.650 ;
        RECT 596.400 723.900 597.600 724.650 ;
        RECT 605.400 723.900 606.450 754.950 ;
        RECT 608.400 742.050 609.450 772.950 ;
        RECT 610.950 769.950 613.050 772.050 ;
        RECT 607.950 739.950 610.050 742.050 ;
        RECT 587.400 709.050 588.450 721.950 ;
        RECT 589.950 721.800 592.050 723.900 ;
        RECT 595.950 721.800 598.050 723.900 ;
        RECT 604.950 721.800 607.050 723.900 ;
        RECT 604.950 712.950 607.050 715.050 ;
        RECT 583.800 706.950 585.900 709.050 ;
        RECT 586.950 706.950 589.050 709.050 ;
        RECT 580.950 694.950 583.050 697.050 ;
        RECT 568.950 691.950 571.050 694.050 ;
        RECT 569.400 684.600 570.450 691.950 ;
        RECT 580.950 685.950 583.050 688.050 ;
        RECT 569.400 682.350 570.600 684.600 ;
        RECT 574.950 683.100 577.050 685.200 ;
        RECT 575.400 682.350 576.600 683.100 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 571.950 679.950 574.050 682.050 ;
        RECT 574.950 679.950 577.050 682.050 ;
        RECT 566.400 678.900 567.600 679.650 ;
        RECT 572.400 678.900 573.600 679.650 ;
        RECT 559.950 678.450 562.050 678.900 ;
        RECT 559.950 677.400 564.450 678.450 ;
        RECT 559.950 676.800 562.050 677.400 ;
        RECT 550.950 673.950 553.050 676.050 ;
        RECT 556.950 673.950 559.050 676.050 ;
        RECT 541.950 670.950 544.050 673.050 ;
        RECT 530.400 649.350 531.600 650.100 ;
        RECT 536.400 649.350 537.600 651.000 ;
        RECT 538.950 649.950 541.050 652.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 532.950 646.950 535.050 649.050 ;
        RECT 535.950 646.950 538.050 649.050 ;
        RECT 523.950 643.950 526.050 646.050 ;
        RECT 533.400 645.900 534.600 646.650 ;
        RECT 532.950 643.800 535.050 645.900 ;
        RECT 538.950 643.950 541.050 646.050 ;
        RECT 521.400 642.000 525.450 642.450 ;
        RECT 521.400 641.400 526.050 642.000 ;
        RECT 520.800 637.950 522.900 640.050 ;
        RECT 523.950 637.950 526.050 641.400 ;
        RECT 521.400 631.050 522.450 637.950 ;
        RECT 520.950 628.950 523.050 631.050 ;
        RECT 511.950 625.950 514.050 628.050 ;
        RECT 517.950 625.950 520.050 628.050 ;
        RECT 493.950 610.950 496.050 613.050 ;
        RECT 488.400 605.400 492.450 606.450 ;
        RECT 494.400 606.600 495.450 610.950 ;
        RECT 476.400 599.400 483.450 600.450 ;
        RECT 469.950 592.950 472.050 595.050 ;
        RECT 454.950 573.000 457.050 577.050 ;
        RECT 457.950 574.950 460.050 577.050 ;
        RECT 455.400 571.350 456.600 573.000 ;
        RECT 460.950 572.100 463.050 574.200 ;
        RECT 461.400 571.350 462.600 572.100 ;
        RECT 454.950 568.950 457.050 571.050 ;
        RECT 457.950 568.950 460.050 571.050 ;
        RECT 460.950 568.950 463.050 571.050 ;
        RECT 463.950 568.950 466.050 571.050 ;
        RECT 458.400 566.400 459.600 568.650 ;
        RECT 464.400 567.900 465.600 568.650 ;
        RECT 458.400 565.050 459.450 566.400 ;
        RECT 463.950 565.800 466.050 567.900 ;
        RECT 466.950 565.950 469.050 568.050 ;
        RECT 470.400 567.900 471.450 592.950 ;
        RECT 472.950 574.950 475.050 577.050 ;
        RECT 473.400 568.050 474.450 574.950 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 448.950 562.950 451.050 565.050 ;
        RECT 457.950 562.950 460.050 565.050 ;
        RECT 458.400 559.050 459.450 562.950 ;
        RECT 460.950 559.950 463.050 562.050 ;
        RECT 436.950 556.950 439.050 559.050 ;
        RECT 442.950 556.950 445.050 559.050 ;
        RECT 457.950 556.950 460.050 559.050 ;
        RECT 461.400 556.050 462.450 559.950 ;
        RECT 460.950 553.950 463.050 556.050 ;
        RECT 436.950 547.950 439.050 550.050 ;
        RECT 427.950 541.950 430.050 544.050 ;
        RECT 412.950 532.950 415.050 535.050 ;
        RECT 418.950 532.950 421.050 535.050 ;
        RECT 421.950 532.950 424.050 535.050 ;
        RECT 433.950 532.950 436.050 535.050 ;
        RECT 409.950 529.950 412.050 532.050 ;
        RECT 385.950 494.100 388.050 496.200 ;
        RECT 392.400 495.600 393.450 521.400 ;
        RECT 397.950 517.950 400.050 522.000 ;
        RECT 406.950 520.950 409.050 523.050 ;
        RECT 410.400 514.050 411.450 529.950 ;
        RECT 413.400 520.050 414.450 532.950 ;
        RECT 418.950 528.000 421.050 531.900 ;
        RECT 419.400 526.350 420.600 528.000 ;
        RECT 424.950 527.100 427.050 529.200 ;
        RECT 425.400 526.350 426.600 527.100 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 422.400 522.900 423.600 523.650 ;
        RECT 428.400 522.900 429.600 523.650 ;
        RECT 434.400 522.900 435.450 532.950 ;
        RECT 421.950 520.800 424.050 522.900 ;
        RECT 427.950 520.800 430.050 522.900 ;
        RECT 433.950 520.800 436.050 522.900 ;
        RECT 412.950 517.950 415.050 520.050 ;
        RECT 409.950 511.950 412.050 514.050 ;
        RECT 427.950 505.950 430.050 508.050 ;
        RECT 397.950 499.950 400.050 502.050 ;
        RECT 398.400 495.600 399.450 499.950 ;
        RECT 392.400 493.350 393.600 495.600 ;
        RECT 398.400 493.350 399.600 495.600 ;
        RECT 409.950 494.100 412.050 496.200 ;
        RECT 415.950 494.100 418.050 496.200 ;
        RECT 421.950 494.100 424.050 496.200 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 380.400 473.400 384.450 474.450 ;
        RECT 395.400 488.400 396.600 490.650 ;
        RECT 380.400 457.050 381.450 473.400 ;
        RECT 382.950 469.950 385.050 472.050 ;
        RECT 379.950 454.950 382.050 457.050 ;
        RECT 383.400 450.600 384.450 469.950 ;
        RECT 395.400 469.050 396.450 488.400 ;
        RECT 410.400 487.050 411.450 494.100 ;
        RECT 416.400 493.350 417.600 494.100 ;
        RECT 422.400 493.350 423.600 494.100 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 419.400 489.900 420.600 490.650 ;
        RECT 418.950 487.800 421.050 489.900 ;
        RECT 409.950 484.950 412.050 487.050 ;
        RECT 403.950 478.950 406.050 481.050 ;
        RECT 394.950 466.950 397.050 469.050 ;
        RECT 397.950 460.950 400.050 463.050 ;
        RECT 383.400 448.350 384.600 450.600 ;
        RECT 388.950 449.100 391.050 451.200 ;
        RECT 389.400 448.350 390.600 449.100 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 386.400 444.900 387.600 445.650 ;
        RECT 377.400 443.400 381.450 444.450 ;
        RECT 373.950 416.100 376.050 418.200 ;
        RECT 380.400 417.600 381.450 443.400 ;
        RECT 385.950 442.800 388.050 444.900 ;
        RECT 392.400 443.400 393.600 445.650 ;
        RECT 388.950 424.950 391.050 427.050 ;
        RECT 374.400 415.350 375.600 416.100 ;
        RECT 380.400 415.350 381.600 417.600 ;
        RECT 370.950 412.950 373.050 415.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 376.950 412.950 379.050 415.050 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 353.400 401.400 357.450 402.450 ;
        RECT 371.400 410.400 372.600 412.650 ;
        RECT 377.400 410.400 378.600 412.650 ;
        RECT 349.950 397.950 352.050 400.050 ;
        RECT 329.400 367.050 330.450 371.100 ;
        RECT 335.400 370.350 336.600 372.600 ;
        RECT 340.950 371.100 343.050 373.200 ;
        RECT 341.400 370.350 342.600 371.100 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 328.950 364.950 331.050 367.050 ;
        RECT 338.400 365.400 339.600 367.650 ;
        RECT 344.400 366.900 345.600 367.650 ;
        RECT 313.950 358.950 316.050 361.050 ;
        RECT 322.950 358.950 325.050 361.050 ;
        RECT 310.950 346.950 313.050 349.050 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 293.400 337.350 294.600 339.600 ;
        RECT 299.400 337.350 300.600 339.600 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 292.950 334.950 295.050 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 283.950 328.950 286.050 333.900 ;
        RECT 286.950 331.950 289.050 334.050 ;
        RECT 296.400 333.900 297.600 334.650 ;
        RECT 295.950 331.800 298.050 333.900 ;
        RECT 302.400 332.400 303.600 334.650 ;
        RECT 308.400 333.900 309.450 337.950 ;
        RECT 311.400 333.900 312.450 346.950 ;
        RECT 295.950 328.650 298.050 330.750 ;
        RECT 289.950 322.950 292.050 325.050 ;
        RECT 281.400 292.350 282.600 294.600 ;
        RECT 277.950 289.950 280.050 292.050 ;
        RECT 280.950 289.950 283.050 292.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 271.950 286.950 274.050 289.050 ;
        RECT 278.400 287.400 279.600 289.650 ;
        RECT 284.400 288.000 285.600 289.650 ;
        RECT 278.400 283.050 279.450 287.400 ;
        RECT 283.950 283.950 286.050 288.000 ;
        RECT 262.950 281.400 267.450 282.450 ;
        RECT 262.950 280.950 265.050 281.400 ;
        RECT 277.950 280.950 280.050 283.050 ;
        RECT 244.950 259.950 247.050 262.050 ;
        RECT 250.950 260.100 253.050 262.200 ;
        RECT 251.400 259.350 252.600 260.100 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 248.400 254.400 249.600 256.650 ;
        RECT 248.400 250.050 249.450 254.400 ;
        RECT 253.950 253.800 256.050 255.900 ;
        RECT 247.950 247.950 250.050 250.050 ;
        RECT 241.950 223.950 244.050 226.050 ;
        RECT 239.400 214.350 240.600 216.600 ;
        RECT 244.950 216.000 247.050 220.050 ;
        RECT 245.400 214.350 246.600 216.000 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 242.400 210.900 243.600 211.650 ;
        RECT 254.400 211.050 255.450 253.800 ;
        RECT 257.400 241.050 258.450 280.950 ;
        RECT 263.400 250.050 264.450 280.950 ;
        RECT 284.400 262.200 285.450 283.950 ;
        RECT 286.950 277.950 289.050 280.050 ;
        RECT 268.950 260.100 271.050 262.200 ;
        RECT 275.400 261.450 276.600 261.600 ;
        RECT 275.400 260.400 282.450 261.450 ;
        RECT 269.400 259.350 270.600 260.100 ;
        RECT 275.400 259.350 276.600 260.400 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 272.400 255.900 273.600 256.650 ;
        RECT 271.950 253.800 274.050 255.900 ;
        RECT 281.400 253.050 282.450 260.400 ;
        RECT 283.950 260.100 286.050 262.200 ;
        RECT 280.950 250.950 283.050 253.050 ;
        RECT 262.950 247.950 265.050 250.050 ;
        RECT 256.950 238.950 259.050 241.050 ;
        RECT 256.950 232.950 259.050 235.050 ;
        RECT 241.950 208.800 244.050 210.900 ;
        RECT 253.950 208.950 256.050 211.050 ;
        RECT 241.950 202.950 244.050 205.050 ;
        RECT 242.400 183.600 243.450 202.950 ;
        RECT 253.950 190.950 256.050 193.050 ;
        RECT 254.400 186.450 255.450 190.950 ;
        RECT 257.400 190.050 258.450 232.950 ;
        RECT 284.400 226.050 285.450 260.100 ;
        RECT 287.400 256.050 288.450 277.950 ;
        RECT 290.400 268.050 291.450 322.950 ;
        RECT 292.950 298.950 295.050 301.050 ;
        RECT 293.400 277.050 294.450 298.950 ;
        RECT 296.400 280.050 297.450 328.650 ;
        RECT 302.400 328.050 303.450 332.400 ;
        RECT 307.800 331.800 309.900 333.900 ;
        RECT 310.950 331.800 313.050 333.900 ;
        RECT 301.950 325.950 304.050 328.050 ;
        RECT 314.400 316.050 315.450 358.950 ;
        RECT 322.950 338.100 325.050 340.200 ;
        RECT 323.400 337.350 324.600 338.100 ;
        RECT 334.950 337.950 337.050 340.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 320.400 333.900 321.600 334.650 ;
        RECT 326.400 333.900 327.600 334.650 ;
        RECT 335.400 333.900 336.450 337.950 ;
        RECT 319.950 331.800 322.050 333.900 ;
        RECT 325.950 331.800 328.050 333.900 ;
        RECT 334.950 331.800 337.050 333.900 ;
        RECT 326.400 328.050 327.450 331.800 ;
        RECT 325.950 325.950 328.050 328.050 ;
        RECT 338.400 322.050 339.450 365.400 ;
        RECT 343.950 364.800 346.050 366.900 ;
        RECT 350.400 343.050 351.450 397.950 ;
        RECT 353.400 367.050 354.450 401.400 ;
        RECT 371.400 400.050 372.450 410.400 ;
        RECT 370.950 397.950 373.050 400.050 ;
        RECT 377.400 391.050 378.450 410.400 ;
        RECT 385.950 409.800 388.050 411.900 ;
        RECT 382.950 397.950 385.050 400.050 ;
        RECT 376.950 388.950 379.050 391.050 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 355.950 376.950 358.050 379.050 ;
        RECT 352.950 364.950 355.050 367.050 ;
        RECT 356.400 364.050 357.450 376.950 ;
        RECT 359.400 376.050 360.450 382.950 ;
        RECT 379.950 376.950 382.050 379.050 ;
        RECT 358.950 373.950 361.050 376.050 ;
        RECT 355.950 361.950 358.050 364.050 ;
        RECT 359.400 352.050 360.450 373.950 ;
        RECT 370.950 372.000 373.050 376.050 ;
        RECT 380.400 372.600 381.450 376.950 ;
        RECT 371.400 370.350 372.600 372.000 ;
        RECT 380.400 370.350 381.600 372.600 ;
        RECT 364.800 367.950 366.900 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 373.950 367.950 376.050 370.050 ;
        RECT 379.500 367.950 381.600 370.050 ;
        RECT 365.400 365.400 366.600 367.650 ;
        RECT 374.400 366.000 375.600 367.650 ;
        RECT 358.950 349.950 361.050 352.050 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 349.950 340.950 352.050 343.050 ;
        RECT 346.950 338.100 349.050 340.200 ;
        RECT 347.400 337.350 348.600 338.100 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 344.400 332.400 345.600 334.650 ;
        RECT 350.400 333.900 351.600 334.650 ;
        RECT 340.950 325.950 343.050 328.050 ;
        RECT 322.950 319.950 325.050 322.050 ;
        RECT 337.950 319.950 340.050 322.050 ;
        RECT 313.950 313.950 316.050 316.050 ;
        RECT 301.950 293.100 304.050 295.200 ;
        RECT 307.950 294.000 310.050 298.050 ;
        RECT 302.400 292.350 303.600 293.100 ;
        RECT 308.400 292.350 309.600 294.000 ;
        RECT 316.950 293.100 319.050 295.200 ;
        RECT 301.950 289.950 304.050 292.050 ;
        RECT 304.950 289.950 307.050 292.050 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 305.400 287.400 306.600 289.650 ;
        RECT 311.400 288.000 312.600 289.650 ;
        RECT 317.400 289.050 318.450 293.100 ;
        RECT 295.950 277.950 298.050 280.050 ;
        RECT 292.950 274.950 295.050 277.050 ;
        RECT 305.400 274.050 306.450 287.400 ;
        RECT 310.950 283.950 313.050 288.000 ;
        RECT 316.950 286.950 319.050 289.050 ;
        RECT 323.400 286.050 324.450 319.950 ;
        RECT 328.950 313.950 331.050 316.050 ;
        RECT 329.400 294.600 330.450 313.950 ;
        RECT 329.400 292.350 330.600 294.600 ;
        RECT 334.950 293.100 337.050 295.200 ;
        RECT 335.400 292.350 336.600 293.100 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 332.400 288.900 333.600 289.650 ;
        RECT 331.950 286.800 334.050 288.900 ;
        RECT 322.950 283.950 325.050 286.050 ;
        RECT 325.950 277.950 328.050 280.050 ;
        RECT 307.950 274.950 310.050 277.050 ;
        RECT 304.950 271.950 307.050 274.050 ;
        RECT 289.950 265.950 292.050 268.050 ;
        RECT 304.950 265.950 307.050 268.050 ;
        RECT 295.950 260.100 298.050 262.200 ;
        RECT 296.400 259.350 297.600 260.100 ;
        RECT 301.950 259.950 304.050 262.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 286.950 253.950 289.050 256.050 ;
        RECT 293.400 254.400 294.600 256.650 ;
        RECT 293.400 253.050 294.450 254.400 ;
        RECT 292.950 250.950 295.050 253.050 ;
        RECT 265.950 223.950 268.050 226.050 ;
        RECT 283.950 223.950 286.050 226.050 ;
        RECT 266.400 216.600 267.450 223.950 ;
        RECT 293.400 223.050 294.450 250.950 ;
        RECT 302.400 247.050 303.450 259.950 ;
        RECT 301.950 244.950 304.050 247.050 ;
        RECT 305.400 229.050 306.450 265.950 ;
        RECT 308.400 255.900 309.450 274.950 ;
        RECT 316.950 260.100 319.050 262.200 ;
        RECT 317.400 259.350 318.600 260.100 ;
        RECT 326.400 259.200 327.450 277.950 ;
        RECT 331.950 274.950 334.050 277.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 325.950 257.100 328.050 259.200 ;
        RECT 314.400 255.900 315.600 256.650 ;
        RECT 307.950 253.800 310.050 255.900 ;
        RECT 313.950 253.800 316.050 255.900 ;
        RECT 320.400 254.400 321.600 256.650 ;
        RECT 326.400 256.350 327.600 257.100 ;
        RECT 310.950 244.950 313.050 247.050 ;
        RECT 295.950 226.950 298.050 229.050 ;
        RECT 304.950 226.950 307.050 229.050 ;
        RECT 292.950 220.950 295.050 223.050 ;
        RECT 266.400 214.350 267.600 216.600 ;
        RECT 271.950 215.100 274.050 217.200 ;
        RECT 277.950 215.100 280.050 217.200 ;
        RECT 283.950 215.100 286.050 217.200 ;
        RECT 289.950 215.100 292.050 217.200 ;
        RECT 296.400 216.600 297.450 226.950 ;
        RECT 304.950 220.950 307.050 223.050 ;
        RECT 272.400 214.350 273.600 215.100 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 263.400 209.400 264.600 211.650 ;
        RECT 269.400 210.900 270.600 211.650 ;
        RECT 256.950 187.950 259.050 190.050 ;
        RECT 263.400 187.050 264.450 209.400 ;
        RECT 268.950 208.800 271.050 210.900 ;
        RECT 278.400 205.050 279.450 215.100 ;
        RECT 277.950 202.950 280.050 205.050 ;
        RECT 251.400 185.400 255.450 186.450 ;
        RECT 242.400 181.350 243.600 183.600 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 239.400 177.000 240.600 178.650 ;
        RECT 245.400 177.900 246.600 178.650 ;
        RECT 232.950 172.950 235.050 175.050 ;
        RECT 238.950 172.950 241.050 177.000 ;
        RECT 244.950 175.800 247.050 177.900 ;
        RECT 244.950 151.950 247.050 154.050 ;
        RECT 235.950 142.950 238.050 145.050 ;
        RECT 229.950 136.950 232.050 139.050 ;
        RECT 236.400 138.600 237.450 142.950 ;
        RECT 236.400 136.350 237.600 138.600 ;
        RECT 232.950 133.950 235.050 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 233.400 132.900 234.600 133.650 ;
        RECT 232.950 130.800 235.050 132.900 ;
        RECT 239.400 132.000 240.600 133.650 ;
        RECT 238.950 127.950 241.050 132.000 ;
        RECT 245.400 127.050 246.450 151.950 ;
        RECT 247.950 142.950 250.050 145.050 ;
        RECT 244.950 124.950 247.050 127.050 ;
        RECT 245.400 108.450 246.450 124.950 ;
        RECT 242.400 107.400 246.450 108.450 ;
        RECT 235.950 104.100 238.050 106.200 ;
        RECT 242.400 105.600 243.450 107.400 ;
        RECT 236.400 103.350 237.600 104.100 ;
        RECT 242.400 103.350 243.600 105.600 ;
        RECT 248.400 105.450 249.450 142.950 ;
        RECT 251.400 130.050 252.450 185.400 ;
        RECT 262.950 184.950 265.050 187.050 ;
        RECT 253.950 182.100 256.050 184.200 ;
        RECT 265.950 182.100 268.050 184.200 ;
        RECT 271.950 183.000 274.050 187.050 ;
        RECT 280.950 184.950 283.050 187.050 ;
        RECT 254.400 166.050 255.450 182.100 ;
        RECT 266.400 181.350 267.600 182.100 ;
        RECT 272.400 181.350 273.600 183.000 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 263.400 177.900 264.600 178.650 ;
        RECT 256.950 175.800 259.050 177.900 ;
        RECT 262.950 175.800 265.050 177.900 ;
        RECT 269.400 176.400 270.600 178.650 ;
        RECT 275.400 176.400 276.600 178.650 ;
        RECT 281.400 177.450 282.450 184.950 ;
        RECT 278.400 176.400 282.450 177.450 ;
        RECT 253.950 163.950 256.050 166.050 ;
        RECT 257.400 139.200 258.450 175.800 ;
        RECT 269.400 166.050 270.450 176.400 ;
        RECT 275.400 172.050 276.450 176.400 ;
        RECT 274.950 169.950 277.050 172.050 ;
        RECT 268.950 163.950 271.050 166.050 ;
        RECT 271.950 145.950 274.050 148.050 ;
        RECT 262.950 142.950 265.050 145.050 ;
        RECT 256.950 137.100 259.050 139.200 ;
        RECT 263.400 138.600 264.450 142.950 ;
        RECT 257.400 136.350 258.600 137.100 ;
        RECT 263.400 136.350 264.600 138.600 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 260.400 131.400 261.600 133.650 ;
        RECT 266.400 132.900 267.600 133.650 ;
        RECT 250.950 127.950 253.050 130.050 ;
        RECT 260.400 127.050 261.450 131.400 ;
        RECT 265.950 130.800 268.050 132.900 ;
        RECT 259.950 124.950 262.050 127.050 ;
        RECT 268.950 124.950 271.050 127.050 ;
        RECT 256.950 123.450 259.050 124.050 ;
        RECT 262.950 123.450 265.050 124.050 ;
        RECT 256.950 122.400 265.050 123.450 ;
        RECT 256.950 121.950 259.050 122.400 ;
        RECT 262.950 121.950 265.050 122.400 ;
        RECT 269.400 118.050 270.450 124.950 ;
        RECT 268.950 115.950 271.050 118.050 ;
        RECT 256.950 109.950 259.050 112.050 ;
        RECT 265.950 109.950 268.050 112.050 ;
        RECT 248.400 104.400 252.450 105.450 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 239.400 99.900 240.600 100.650 ;
        RECT 245.400 99.900 246.600 100.650 ;
        RECT 251.400 99.900 252.450 104.400 ;
        RECT 238.950 97.800 241.050 99.900 ;
        RECT 244.950 97.800 247.050 99.900 ;
        RECT 250.950 97.800 253.050 99.900 ;
        RECT 250.950 79.950 253.050 82.050 ;
        RECT 229.950 76.950 232.050 79.050 ;
        RECT 230.400 70.050 231.450 76.950 ;
        RECT 229.950 67.950 232.050 70.050 ;
        RECT 230.400 55.050 231.450 67.950 ;
        RECT 238.950 59.100 241.050 61.200 ;
        RECT 251.400 61.050 252.450 79.950 ;
        RECT 257.400 67.050 258.450 109.950 ;
        RECT 266.400 105.600 267.450 109.950 ;
        RECT 272.400 105.600 273.450 145.950 ;
        RECT 274.950 137.100 277.050 139.200 ;
        RECT 275.400 118.050 276.450 137.100 ;
        RECT 278.400 133.050 279.450 176.400 ;
        RECT 284.400 154.050 285.450 215.100 ;
        RECT 290.400 214.350 291.600 215.100 ;
        RECT 296.400 214.350 297.600 216.600 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 293.400 209.400 294.600 211.650 ;
        RECT 299.400 210.900 300.600 211.650 ;
        RECT 305.400 210.900 306.450 220.950 ;
        RECT 293.400 202.050 294.450 209.400 ;
        RECT 298.950 208.800 301.050 210.900 ;
        RECT 304.950 208.800 307.050 210.900 ;
        RECT 292.950 199.950 295.050 202.050 ;
        RECT 298.950 187.950 301.050 190.050 ;
        RECT 292.950 182.100 295.050 184.200 ;
        RECT 299.400 183.600 300.450 187.950 ;
        RECT 293.400 181.350 294.600 182.100 ;
        RECT 299.400 181.350 300.600 183.600 ;
        RECT 307.950 181.950 310.050 184.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 296.400 177.000 297.600 178.650 ;
        RECT 295.950 172.950 298.050 177.000 ;
        RECT 302.400 176.400 303.600 178.650 ;
        RECT 302.400 172.050 303.450 176.400 ;
        RECT 308.400 175.050 309.450 181.950 ;
        RECT 311.400 177.900 312.450 244.950 ;
        RECT 320.400 244.050 321.450 254.400 ;
        RECT 322.950 253.950 325.050 256.050 ;
        RECT 326.100 253.950 328.200 256.050 ;
        RECT 323.400 250.050 324.450 253.950 ;
        RECT 322.950 247.950 325.050 250.050 ;
        RECT 319.950 241.950 322.050 244.050 ;
        RECT 316.950 220.950 319.050 223.050 ;
        RECT 317.400 216.600 318.450 220.950 ;
        RECT 320.400 220.050 321.450 241.950 ;
        RECT 322.950 226.950 325.050 229.050 ;
        RECT 328.950 226.950 331.050 229.050 ;
        RECT 319.950 217.950 322.050 220.050 ;
        RECT 323.400 217.200 324.450 226.950 ;
        RECT 317.400 214.350 318.600 216.600 ;
        RECT 322.950 215.100 325.050 217.200 ;
        RECT 323.400 214.350 324.600 215.100 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 320.400 209.400 321.600 211.650 ;
        RECT 329.400 210.450 330.450 226.950 ;
        RECT 326.400 209.400 330.450 210.450 ;
        RECT 320.400 205.050 321.450 209.400 ;
        RECT 319.950 202.950 322.050 205.050 ;
        RECT 313.950 196.950 316.050 199.050 ;
        RECT 310.950 175.800 313.050 177.900 ;
        RECT 307.950 172.950 310.050 175.050 ;
        RECT 314.400 174.450 315.450 196.950 ;
        RECT 316.950 190.950 319.050 193.050 ;
        RECT 317.400 187.050 318.450 190.950 ;
        RECT 320.400 190.050 321.450 202.950 ;
        RECT 326.400 199.050 327.450 209.400 ;
        RECT 328.950 205.950 331.050 208.050 ;
        RECT 325.950 196.950 328.050 199.050 ;
        RECT 329.400 193.050 330.450 205.950 ;
        RECT 328.950 190.950 331.050 193.050 ;
        RECT 319.950 187.950 322.050 190.050 ;
        RECT 316.950 184.950 319.050 187.050 ;
        RECT 322.950 182.100 325.050 184.200 ;
        RECT 329.400 183.600 330.450 190.950 ;
        RECT 332.400 187.050 333.450 274.950 ;
        RECT 334.950 258.000 337.050 262.050 ;
        RECT 335.400 256.350 336.600 258.000 ;
        RECT 335.100 253.950 337.200 256.050 ;
        RECT 334.950 247.950 337.050 250.050 ;
        RECT 335.400 208.050 336.450 247.950 ;
        RECT 341.400 238.050 342.450 325.950 ;
        RECT 344.400 316.050 345.450 332.400 ;
        RECT 349.950 331.800 352.050 333.900 ;
        RECT 356.400 328.050 357.450 343.950 ;
        RECT 365.400 340.200 366.450 365.400 ;
        RECT 373.950 361.950 376.050 366.000 ;
        RECT 373.950 352.950 376.050 355.050 ;
        RECT 358.950 338.100 361.050 340.200 ;
        RECT 364.950 338.100 367.050 340.200 ;
        RECT 359.400 328.050 360.450 338.100 ;
        RECT 365.400 337.350 366.600 338.100 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 374.400 336.600 375.450 352.950 ;
        RECT 376.800 349.950 378.900 352.050 ;
        RECT 379.950 349.950 382.050 352.050 ;
        RECT 377.400 337.050 378.450 349.950 ;
        RECT 368.400 333.900 369.600 334.650 ;
        RECT 374.400 334.350 375.600 336.600 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 367.950 331.800 370.050 333.900 ;
        RECT 374.100 331.950 376.200 334.050 ;
        RECT 355.950 325.950 358.050 328.050 ;
        RECT 358.950 325.950 361.050 328.050 ;
        RECT 361.950 325.950 364.050 328.050 ;
        RECT 343.950 313.950 346.050 316.050 ;
        RECT 344.400 277.050 345.450 313.950 ;
        RECT 362.400 301.050 363.450 325.950 ;
        RECT 380.400 322.050 381.450 349.950 ;
        RECT 383.400 336.600 384.450 397.950 ;
        RECT 386.400 346.050 387.450 409.800 ;
        RECT 389.400 400.050 390.450 424.950 ;
        RECT 388.950 397.950 391.050 400.050 ;
        RECT 392.400 352.050 393.450 443.400 ;
        RECT 398.400 433.050 399.450 460.950 ;
        RECT 400.950 454.950 403.050 457.050 ;
        RECT 401.400 436.050 402.450 454.950 ;
        RECT 400.950 433.950 403.050 436.050 ;
        RECT 397.950 430.950 400.050 433.050 ;
        RECT 401.400 427.050 402.450 433.950 ;
        RECT 404.400 432.450 405.450 478.950 ;
        RECT 424.950 469.950 427.050 472.050 ;
        RECT 415.950 466.950 418.050 469.050 ;
        RECT 409.950 449.100 412.050 451.200 ;
        RECT 416.400 450.600 417.450 466.950 ;
        RECT 421.950 451.950 424.050 454.050 ;
        RECT 410.400 448.350 411.600 449.100 ;
        RECT 416.400 448.350 417.600 450.600 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 413.400 444.900 414.600 445.650 ;
        RECT 412.950 442.800 415.050 444.900 ;
        RECT 418.950 439.950 421.050 442.050 ;
        RECT 404.400 431.400 408.450 432.450 ;
        RECT 403.950 427.950 406.050 430.050 ;
        RECT 400.950 424.950 403.050 427.050 ;
        RECT 404.400 420.450 405.450 427.950 ;
        RECT 401.400 419.400 405.450 420.450 ;
        RECT 401.400 417.600 402.450 419.400 ;
        RECT 407.400 417.600 408.450 431.400 ;
        RECT 415.950 424.950 418.050 427.050 ;
        RECT 401.400 415.350 402.600 417.600 ;
        RECT 407.400 415.350 408.600 417.600 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 398.400 411.900 399.600 412.650 ;
        RECT 397.950 409.800 400.050 411.900 ;
        RECT 404.400 410.400 405.600 412.650 ;
        RECT 410.400 411.000 411.600 412.650 ;
        RECT 404.400 406.050 405.450 410.400 ;
        RECT 409.950 406.950 412.050 411.000 ;
        RECT 416.400 409.050 417.450 424.950 ;
        RECT 419.400 411.900 420.450 439.950 ;
        RECT 422.400 427.050 423.450 451.950 ;
        RECT 425.400 430.050 426.450 469.950 ;
        RECT 428.400 454.050 429.450 505.950 ;
        RECT 437.400 496.200 438.450 547.950 ;
        RECT 439.950 541.950 442.050 544.050 ;
        RECT 440.400 522.900 441.450 541.950 ;
        RECT 457.950 538.950 460.050 541.050 ;
        RECT 454.950 529.950 457.050 532.050 ;
        RECT 448.950 527.100 451.050 529.200 ;
        RECT 449.400 526.350 450.600 527.100 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 448.950 523.950 451.050 526.050 ;
        RECT 446.400 522.900 447.600 523.650 ;
        RECT 455.400 523.050 456.450 529.950 ;
        RECT 439.950 520.800 442.050 522.900 ;
        RECT 445.950 520.800 448.050 522.900 ;
        RECT 454.950 520.950 457.050 523.050 ;
        RECT 448.950 511.950 451.050 514.050 ;
        RECT 436.950 494.100 439.050 496.200 ;
        RECT 442.950 494.100 445.050 496.200 ;
        RECT 449.400 495.600 450.450 511.950 ;
        RECT 458.400 508.050 459.450 538.950 ;
        RECT 467.400 532.050 468.450 565.950 ;
        RECT 469.950 565.800 472.050 567.900 ;
        RECT 472.950 565.950 475.050 568.050 ;
        RECT 476.400 565.050 477.450 568.950 ;
        RECT 479.400 565.050 480.450 599.400 ;
        RECT 484.950 598.800 487.050 600.900 ;
        RECT 485.400 574.200 486.450 598.800 ;
        RECT 488.400 577.050 489.450 605.400 ;
        RECT 494.400 604.350 495.600 606.600 ;
        RECT 499.950 606.000 502.050 610.050 ;
        RECT 505.800 607.950 507.900 610.050 ;
        RECT 508.950 607.950 511.050 610.050 ;
        RECT 500.400 604.350 501.600 606.000 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 496.950 601.950 499.050 604.050 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 497.400 600.900 498.600 601.650 ;
        RECT 496.950 598.800 499.050 600.900 ;
        RECT 493.950 592.950 496.050 595.050 ;
        RECT 487.950 574.950 490.050 577.050 ;
        RECT 484.950 572.100 487.050 574.200 ;
        RECT 485.400 571.350 486.600 572.100 ;
        RECT 482.100 568.950 484.200 571.050 ;
        RECT 485.400 568.950 487.500 571.050 ;
        RECT 490.800 568.950 492.900 571.050 ;
        RECT 482.400 566.400 483.600 568.650 ;
        RECT 491.400 567.450 492.600 568.650 ;
        RECT 494.400 567.450 495.450 592.950 ;
        RECT 506.400 589.050 507.450 607.950 ;
        RECT 505.950 586.950 508.050 589.050 ;
        RECT 509.400 577.200 510.450 607.950 ;
        RECT 496.950 574.950 499.050 577.050 ;
        RECT 502.950 574.950 505.050 577.050 ;
        RECT 508.950 575.100 511.050 577.200 ;
        RECT 512.400 577.050 513.450 625.950 ;
        RECT 529.950 616.950 532.050 619.050 ;
        RECT 522.000 609.450 526.050 610.050 ;
        RECT 521.400 607.950 526.050 609.450 ;
        RECT 521.400 606.600 522.450 607.950 ;
        RECT 521.400 604.350 522.600 606.600 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 520.950 601.950 523.050 604.050 ;
        RECT 523.950 601.950 526.050 604.050 ;
        RECT 518.400 600.900 519.600 601.650 ;
        RECT 524.400 600.900 525.600 601.650 ;
        RECT 530.400 600.900 531.450 616.950 ;
        RECT 539.400 610.050 540.450 643.950 ;
        RECT 542.400 613.050 543.450 670.950 ;
        RECT 544.950 661.950 547.050 664.050 ;
        RECT 545.400 622.050 546.450 661.950 ;
        RECT 547.950 652.950 550.050 655.050 ;
        RECT 548.400 637.050 549.450 652.950 ;
        RECT 551.400 652.050 552.450 673.950 ;
        RECT 553.950 661.950 556.050 664.050 ;
        RECT 554.400 652.200 555.450 661.950 ;
        RECT 550.800 649.950 552.900 652.050 ;
        RECT 553.950 650.100 556.050 652.200 ;
        RECT 554.400 649.350 555.600 650.100 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 556.950 646.950 559.050 649.050 ;
        RECT 550.950 643.950 553.050 646.050 ;
        RECT 557.400 644.400 558.600 646.650 ;
        RECT 547.950 634.950 550.050 637.050 ;
        RECT 544.950 619.950 547.050 622.050 ;
        RECT 541.950 610.950 544.050 613.050 ;
        RECT 538.950 607.950 541.050 610.050 ;
        RECT 541.950 606.000 544.050 609.900 ;
        RECT 548.400 606.450 549.600 606.600 ;
        RECT 551.400 606.450 552.450 643.950 ;
        RECT 557.400 637.050 558.450 644.400 ;
        RECT 556.950 634.950 559.050 637.050 ;
        RECT 553.950 613.950 556.050 616.050 ;
        RECT 542.400 604.350 543.600 606.000 ;
        RECT 548.400 605.400 552.450 606.450 ;
        RECT 548.400 604.350 549.600 605.400 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 517.950 598.800 520.050 600.900 ;
        RECT 523.950 598.800 526.050 600.900 ;
        RECT 529.950 598.800 532.050 600.900 ;
        RECT 545.400 599.400 546.600 601.650 ;
        RECT 514.950 580.950 517.050 583.050 ;
        RECT 545.400 582.450 546.450 599.400 ;
        RECT 554.400 592.050 555.450 613.950 ;
        RECT 563.400 607.050 564.450 677.400 ;
        RECT 565.950 676.800 568.050 678.900 ;
        RECT 571.950 676.800 574.050 678.900 ;
        RECT 581.400 670.050 582.450 685.950 ;
        RECT 584.400 682.050 585.450 706.950 ;
        RECT 586.950 697.950 589.050 700.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 580.950 667.950 583.050 670.050 ;
        RECT 568.950 664.950 571.050 667.050 ;
        RECT 565.950 649.950 568.050 652.050 ;
        RECT 566.400 631.050 567.450 649.950 ;
        RECT 565.950 628.950 568.050 631.050 ;
        RECT 569.400 616.050 570.450 664.950 ;
        RECT 577.950 650.100 580.050 652.200 ;
        RECT 578.400 649.350 579.600 650.100 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 580.950 646.950 583.050 649.050 ;
        RECT 575.400 645.900 576.600 646.650 ;
        RECT 581.400 645.900 582.600 646.650 ;
        RECT 574.950 643.800 577.050 645.900 ;
        RECT 580.950 643.800 583.050 645.900 ;
        RECT 571.950 628.950 574.050 631.050 ;
        RECT 568.950 613.950 571.050 616.050 ;
        RECT 565.950 610.950 568.050 613.050 ;
        RECT 562.950 604.950 565.050 607.050 ;
        RECT 566.400 606.600 567.450 610.950 ;
        RECT 572.400 606.600 573.450 628.950 ;
        RECT 587.400 619.050 588.450 697.950 ;
        RECT 592.950 688.950 595.050 691.050 ;
        RECT 598.950 688.950 601.050 691.050 ;
        RECT 593.400 684.600 594.450 688.950 ;
        RECT 599.400 684.600 600.450 688.950 ;
        RECT 593.400 682.350 594.600 684.600 ;
        RECT 599.400 682.350 600.600 684.600 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 596.400 677.400 597.600 679.650 ;
        RECT 592.950 673.950 595.050 676.050 ;
        RECT 589.950 658.950 592.050 661.050 ;
        RECT 590.400 645.900 591.450 658.950 ;
        RECT 589.950 643.800 592.050 645.900 ;
        RECT 589.950 631.950 592.050 634.050 ;
        RECT 586.950 616.950 589.050 619.050 ;
        RECT 580.950 607.950 583.050 610.050 ;
        RECT 566.400 604.350 567.600 606.600 ;
        RECT 572.400 604.350 573.600 606.600 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 571.950 601.950 574.050 604.050 ;
        RECT 569.400 599.400 570.600 601.650 ;
        RECT 569.400 595.050 570.450 599.400 ;
        RECT 568.950 592.950 571.050 595.050 ;
        RECT 553.950 589.950 556.050 592.050 ;
        RECT 574.950 583.950 577.050 586.050 ;
        RECT 545.400 581.400 549.450 582.450 ;
        RECT 515.400 577.050 516.450 580.950 ;
        RECT 511.950 574.950 514.050 577.050 ;
        RECT 491.400 566.400 495.450 567.450 ;
        RECT 475.950 562.950 478.050 565.050 ;
        RECT 478.950 562.950 481.050 565.050 ;
        RECT 482.400 556.050 483.450 566.400 ;
        RECT 484.950 556.950 487.050 559.050 ;
        RECT 481.950 553.950 484.050 556.050 ;
        RECT 481.950 547.950 484.050 550.050 ;
        RECT 460.950 529.950 463.050 532.050 ;
        RECT 466.950 529.950 469.050 532.050 ;
        RECT 457.950 505.950 460.050 508.050 ;
        RECT 454.950 499.950 457.050 502.050 ;
        RECT 443.400 493.350 444.600 494.100 ;
        RECT 449.400 493.350 450.600 495.600 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 440.400 489.900 441.600 490.650 ;
        RECT 439.950 487.800 442.050 489.900 ;
        RECT 446.400 488.400 447.600 490.650 ;
        RECT 440.400 472.050 441.450 487.800 ;
        RECT 439.950 469.950 442.050 472.050 ;
        RECT 440.400 454.050 441.450 469.950 ;
        RECT 446.400 469.050 447.450 488.400 ;
        RECT 445.950 466.950 448.050 469.050 ;
        RECT 427.950 451.950 430.050 454.050 ;
        RECT 439.950 451.950 442.050 454.050 ;
        RECT 445.950 451.950 448.050 454.050 ;
        RECT 451.950 451.950 454.050 454.050 ;
        RECT 427.950 448.800 430.050 450.900 ;
        RECT 436.950 449.100 439.050 451.200 ;
        RECT 424.950 427.950 427.050 430.050 ;
        RECT 421.950 424.950 424.050 427.050 ;
        RECT 428.400 424.050 429.450 448.800 ;
        RECT 437.400 448.350 438.600 449.100 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 434.400 444.900 435.600 445.650 ;
        RECT 433.950 442.800 436.050 444.900 ;
        RECT 440.400 443.400 441.600 445.650 ;
        RECT 440.400 433.050 441.450 443.400 ;
        RECT 439.950 430.950 442.050 433.050 ;
        RECT 436.950 424.950 439.050 427.050 ;
        RECT 427.950 421.950 430.050 424.050 ;
        RECT 421.950 416.100 424.050 418.200 ;
        RECT 430.950 416.100 433.050 418.200 ;
        RECT 437.400 417.600 438.450 424.950 ;
        RECT 418.950 409.800 421.050 411.900 ;
        RECT 415.950 406.950 418.050 409.050 ;
        RECT 403.950 403.950 406.050 406.050 ;
        RECT 422.400 385.050 423.450 416.100 ;
        RECT 431.400 415.350 432.600 416.100 ;
        RECT 437.400 415.350 438.600 417.600 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 433.950 412.950 436.050 415.050 ;
        RECT 436.950 412.950 439.050 415.050 ;
        RECT 428.400 411.000 429.600 412.650 ;
        RECT 434.400 411.900 435.600 412.650 ;
        RECT 427.950 406.950 430.050 411.000 ;
        RECT 433.950 409.800 436.050 411.900 ;
        RECT 442.950 409.950 445.050 412.050 ;
        RECT 433.950 408.300 436.050 408.750 ;
        RECT 439.950 408.300 442.050 408.750 ;
        RECT 433.950 407.250 442.050 408.300 ;
        RECT 433.950 406.650 436.050 407.250 ;
        RECT 439.950 406.650 442.050 407.250 ;
        RECT 430.950 397.950 433.050 400.050 ;
        RECT 421.950 382.950 424.050 385.050 ;
        RECT 431.400 373.200 432.450 397.950 ;
        RECT 439.950 385.950 442.050 388.050 ;
        RECT 440.400 379.050 441.450 385.950 ;
        RECT 439.950 376.950 442.050 379.050 ;
        RECT 400.950 371.100 403.050 373.200 ;
        RECT 410.400 372.450 411.600 372.600 ;
        RECT 410.400 371.400 414.450 372.450 ;
        RECT 401.400 370.350 402.600 371.100 ;
        RECT 410.400 370.350 411.600 371.400 ;
        RECT 401.100 367.950 403.200 370.050 ;
        RECT 406.500 367.950 408.600 370.050 ;
        RECT 409.800 367.950 411.900 370.050 ;
        RECT 407.400 366.900 408.600 367.650 ;
        RECT 406.950 364.800 409.050 366.900 ;
        RECT 413.400 352.050 414.450 371.400 ;
        RECT 430.950 371.100 433.050 373.200 ;
        RECT 436.950 371.100 439.050 373.200 ;
        RECT 431.400 370.350 432.600 371.100 ;
        RECT 437.400 370.350 438.600 371.100 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 428.400 366.900 429.600 367.650 ;
        RECT 427.950 364.800 430.050 366.900 ;
        RECT 434.400 365.400 435.600 367.650 ;
        RECT 443.400 366.900 444.450 409.950 ;
        RECT 446.400 373.200 447.450 451.950 ;
        RECT 448.950 448.950 451.050 451.050 ;
        RECT 449.400 418.200 450.450 448.950 ;
        RECT 452.400 439.050 453.450 451.950 ;
        RECT 455.400 451.050 456.450 499.950 ;
        RECT 457.950 493.950 460.050 496.050 ;
        RECT 458.400 489.900 459.450 493.950 ;
        RECT 457.950 487.800 460.050 489.900 ;
        RECT 461.400 478.050 462.450 529.950 ;
        RECT 469.950 527.100 472.050 529.200 ;
        RECT 475.950 528.000 478.050 532.050 ;
        RECT 470.400 526.350 471.600 527.100 ;
        RECT 476.400 526.350 477.600 528.000 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 475.950 523.950 478.050 526.050 ;
        RECT 467.400 522.900 468.600 523.650 ;
        RECT 473.400 522.900 474.600 523.650 ;
        RECT 482.400 523.050 483.450 547.950 ;
        RECT 485.400 523.050 486.450 556.950 ;
        RECT 493.950 544.950 496.050 547.050 ;
        RECT 487.950 532.950 490.050 535.050 ;
        RECT 478.950 522.900 481.050 523.050 ;
        RECT 466.950 520.800 469.050 522.900 ;
        RECT 472.950 520.800 475.050 522.900 ;
        RECT 478.800 520.950 481.050 522.900 ;
        RECT 481.950 520.950 484.050 523.050 ;
        RECT 484.950 520.950 487.050 523.050 ;
        RECT 478.800 520.800 480.900 520.950 ;
        RECT 469.950 517.950 472.050 520.050 ;
        RECT 481.950 517.800 484.050 519.900 ;
        RECT 488.400 502.050 489.450 532.950 ;
        RECT 494.400 528.600 495.450 544.950 ;
        RECT 497.400 532.050 498.450 574.950 ;
        RECT 499.950 568.950 502.050 571.050 ;
        RECT 500.400 562.050 501.450 568.950 ;
        RECT 499.950 559.950 502.050 562.050 ;
        RECT 503.400 535.050 504.450 574.950 ;
        RECT 508.950 571.950 511.050 574.050 ;
        RECT 514.950 573.000 517.050 577.050 ;
        RECT 523.950 574.950 526.050 577.050 ;
        RECT 532.950 574.950 535.050 580.050 ;
        RECT 544.950 577.950 547.050 580.050 ;
        RECT 509.400 571.350 510.600 571.950 ;
        RECT 515.400 571.350 516.600 573.000 ;
        RECT 520.950 571.950 523.050 574.050 ;
        RECT 508.950 568.950 511.050 571.050 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 512.400 567.900 513.600 568.650 ;
        RECT 511.950 565.800 514.050 567.900 ;
        RECT 508.950 562.950 511.050 565.050 ;
        RECT 502.950 532.950 505.050 535.050 ;
        RECT 496.950 529.950 499.050 532.050 ;
        RECT 494.400 526.350 495.600 528.600 ;
        RECT 499.950 528.000 502.050 532.050 ;
        RECT 500.400 526.350 501.600 528.000 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 490.950 520.950 493.050 523.050 ;
        RECT 497.400 522.000 498.600 523.650 ;
        RECT 503.400 522.900 504.600 523.650 ;
        RECT 491.400 514.050 492.450 520.950 ;
        RECT 496.950 517.950 499.050 522.000 ;
        RECT 502.950 520.800 505.050 522.900 ;
        RECT 490.950 511.950 493.050 514.050 ;
        RECT 502.950 508.950 505.050 511.050 ;
        RECT 487.950 499.950 490.050 502.050 ;
        RECT 496.950 499.950 499.050 502.050 ;
        RECT 468.000 498.450 472.050 499.050 ;
        RECT 467.400 496.950 472.050 498.450 ;
        RECT 467.400 495.600 468.450 496.950 ;
        RECT 487.950 496.800 490.050 498.900 ;
        RECT 467.400 493.350 468.600 495.600 ;
        RECT 472.950 494.100 475.050 496.200 ;
        RECT 473.400 493.350 474.600 494.100 ;
        RECT 466.950 490.950 469.050 493.050 ;
        RECT 469.950 490.950 472.050 493.050 ;
        RECT 472.950 490.950 475.050 493.050 ;
        RECT 475.950 490.950 478.050 493.050 ;
        RECT 484.950 490.950 487.050 493.050 ;
        RECT 470.400 489.900 471.600 490.650 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 476.400 489.450 477.600 490.650 ;
        RECT 476.400 488.400 480.450 489.450 ;
        RECT 479.400 487.050 480.450 488.400 ;
        RECT 478.950 484.950 481.050 487.050 ;
        RECT 460.950 475.950 463.050 478.050 ;
        RECT 475.950 466.950 478.050 469.050 ;
        RECT 454.950 448.950 457.050 451.050 ;
        RECT 460.950 450.000 463.050 454.050 ;
        RECT 476.400 451.200 477.450 466.950 ;
        RECT 467.400 450.450 468.600 450.600 ;
        RECT 461.400 448.350 462.600 450.000 ;
        RECT 467.400 449.400 474.450 450.450 ;
        RECT 467.400 448.350 468.600 449.400 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 458.400 443.400 459.600 445.650 ;
        RECT 464.400 444.900 465.600 445.650 ;
        RECT 451.950 436.950 454.050 439.050 ;
        RECT 458.400 433.050 459.450 443.400 ;
        RECT 463.950 442.800 466.050 444.900 ;
        RECT 473.400 442.050 474.450 449.400 ;
        RECT 475.950 449.100 478.050 451.200 ;
        RECT 472.950 439.950 475.050 442.050 ;
        RECT 463.950 436.950 466.050 439.050 ;
        RECT 457.950 430.950 460.050 433.050 ;
        RECT 460.950 424.950 463.050 427.050 ;
        RECT 448.950 416.100 451.050 418.200 ;
        RECT 457.950 416.100 460.050 418.200 ;
        RECT 449.400 376.050 450.450 416.100 ;
        RECT 458.400 415.350 459.600 416.100 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 455.400 410.400 456.600 412.650 ;
        RECT 455.400 409.050 456.450 410.400 ;
        RECT 451.950 407.400 456.450 409.050 ;
        RECT 451.950 406.950 456.000 407.400 ;
        RECT 464.400 400.050 465.450 436.950 ;
        RECT 472.950 436.800 475.050 438.900 ;
        RECT 466.950 430.950 469.050 433.050 ;
        RECT 467.400 412.050 468.450 430.950 ;
        RECT 473.400 427.050 474.450 436.800 ;
        RECT 476.400 427.050 477.450 449.100 ;
        RECT 479.400 445.050 480.450 484.950 ;
        RECT 485.400 451.200 486.450 490.950 ;
        RECT 488.400 489.900 489.450 496.800 ;
        RECT 497.400 495.600 498.450 499.950 ;
        RECT 503.400 496.200 504.450 508.950 ;
        RECT 497.400 493.350 498.600 495.600 ;
        RECT 502.950 494.100 505.050 496.200 ;
        RECT 503.400 493.350 504.600 494.100 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 499.950 490.950 502.050 493.050 ;
        RECT 502.950 490.950 505.050 493.050 ;
        RECT 494.400 489.900 495.600 490.650 ;
        RECT 487.950 487.800 490.050 489.900 ;
        RECT 493.950 487.800 496.050 489.900 ;
        RECT 500.400 489.000 501.600 490.650 ;
        RECT 499.950 486.450 502.050 489.000 ;
        RECT 497.400 485.400 502.050 486.450 ;
        RECT 497.400 454.050 498.450 485.400 ;
        RECT 499.950 484.950 502.050 485.400 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 503.400 481.050 504.450 484.950 ;
        RECT 509.400 484.050 510.450 562.950 ;
        RECT 514.950 559.950 517.050 562.050 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 512.400 520.050 513.450 529.950 ;
        RECT 511.950 517.950 514.050 520.050 ;
        RECT 515.400 511.050 516.450 559.950 ;
        RECT 521.400 550.050 522.450 571.950 ;
        RECT 524.400 568.050 525.450 574.950 ;
        RECT 533.400 573.600 534.450 574.950 ;
        RECT 533.400 571.350 534.600 573.600 ;
        RECT 538.950 572.100 541.050 574.200 ;
        RECT 539.400 571.350 540.600 572.100 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 523.950 565.950 526.050 568.050 ;
        RECT 520.950 547.950 523.050 550.050 ;
        RECT 520.950 541.950 523.050 544.050 ;
        RECT 521.400 528.600 522.450 541.950 ;
        RECT 527.400 541.050 528.450 568.950 ;
        RECT 536.400 567.000 537.600 568.650 ;
        RECT 545.400 568.050 546.450 577.950 ;
        RECT 535.950 562.950 538.050 567.000 ;
        RECT 544.950 565.950 547.050 568.050 ;
        RECT 548.400 555.450 549.450 581.400 ;
        RECT 550.950 571.950 553.050 574.050 ;
        RECT 559.950 572.100 562.050 574.200 ;
        RECT 565.950 572.100 568.050 574.200 ;
        RECT 551.400 556.050 552.450 571.950 ;
        RECT 560.400 571.350 561.600 572.100 ;
        RECT 566.400 571.350 567.600 572.100 ;
        RECT 556.950 568.950 559.050 571.050 ;
        RECT 559.950 568.950 562.050 571.050 ;
        RECT 562.950 568.950 565.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 557.400 567.900 558.600 568.650 ;
        RECT 556.950 565.800 559.050 567.900 ;
        RECT 563.400 566.400 564.600 568.650 ;
        RECT 569.400 567.900 570.600 568.650 ;
        RECT 545.400 554.400 549.450 555.450 ;
        RECT 541.950 547.950 544.050 550.050 ;
        RECT 526.950 538.950 529.050 541.050 ;
        RECT 527.400 528.600 528.450 538.950 ;
        RECT 521.400 526.350 522.600 528.600 ;
        RECT 527.400 526.350 528.600 528.600 ;
        RECT 536.100 526.950 538.200 529.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 536.400 525.900 537.600 526.650 ;
        RECT 535.950 523.800 538.050 525.900 ;
        RECT 517.950 520.950 520.050 523.050 ;
        RECT 524.400 522.000 525.600 523.650 ;
        RECT 514.950 508.950 517.050 511.050 ;
        RECT 514.950 499.950 517.050 502.050 ;
        RECT 508.950 481.950 511.050 484.050 ;
        RECT 515.400 481.050 516.450 499.950 ;
        RECT 518.400 487.050 519.450 520.950 ;
        RECT 523.950 517.950 526.050 522.000 ;
        RECT 530.400 521.400 531.600 523.650 ;
        RECT 530.400 514.050 531.450 521.400 ;
        RECT 538.950 514.950 541.050 517.050 ;
        RECT 529.950 511.950 532.050 514.050 ;
        RECT 523.800 498.300 525.900 500.400 ;
        RECT 526.950 499.950 529.050 502.050 ;
        RECT 527.400 499.200 528.600 499.950 ;
        RECT 520.950 494.100 523.050 496.200 ;
        RECT 521.400 493.350 522.600 494.100 ;
        RECT 521.100 490.950 523.200 493.050 ;
        RECT 524.100 492.900 525.000 498.300 ;
        RECT 527.100 496.800 529.200 498.900 ;
        RECT 531.000 495.900 533.100 497.700 ;
        RECT 525.900 494.700 534.600 495.900 ;
        RECT 525.900 493.800 528.000 494.700 ;
        RECT 524.100 491.700 531.000 492.900 ;
        RECT 517.950 484.950 520.050 487.050 ;
        RECT 524.100 484.500 525.300 491.700 ;
        RECT 527.100 487.950 529.200 490.050 ;
        RECT 530.100 489.300 531.000 491.700 ;
        RECT 527.400 485.400 528.600 487.650 ;
        RECT 530.100 487.200 532.200 489.300 ;
        RECT 533.700 485.700 534.600 494.700 ;
        RECT 535.800 490.950 537.900 493.050 ;
        RECT 536.400 489.900 537.600 490.650 ;
        RECT 535.950 487.800 538.050 489.900 ;
        RECT 523.800 482.400 525.900 484.500 ;
        RECT 533.400 483.600 535.500 485.700 ;
        RECT 502.950 478.950 505.050 481.050 ;
        RECT 514.950 478.950 517.050 481.050 ;
        RECT 511.950 469.950 514.050 472.050 ;
        RECT 526.950 469.950 529.050 472.050 ;
        RECT 512.400 460.050 513.450 469.950 ;
        RECT 511.950 457.950 514.050 460.050 ;
        RECT 496.950 451.950 499.050 454.050 ;
        RECT 484.950 449.100 487.050 451.200 ;
        RECT 490.950 449.100 493.050 451.200 ;
        RECT 485.400 448.350 486.600 449.100 ;
        RECT 491.400 448.350 492.600 449.100 ;
        RECT 502.950 448.950 505.050 451.050 ;
        RECT 508.950 450.000 511.050 454.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 478.950 442.950 481.050 445.050 ;
        RECT 488.400 444.000 489.600 445.650 ;
        RECT 481.950 439.950 484.050 442.050 ;
        RECT 487.950 439.950 490.050 444.000 ;
        RECT 493.950 442.950 496.050 445.050 ;
        RECT 494.400 436.050 495.450 442.950 ;
        RECT 493.950 433.950 496.050 436.050 ;
        RECT 503.400 430.050 504.450 448.950 ;
        RECT 509.400 448.350 510.600 450.000 ;
        RECT 514.950 449.100 517.050 451.200 ;
        RECT 520.800 449.100 522.900 451.200 ;
        RECT 523.950 449.100 526.050 451.200 ;
        RECT 515.400 448.350 516.600 449.100 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 512.400 443.400 513.600 445.650 ;
        RECT 512.400 439.050 513.450 443.400 ;
        RECT 517.950 439.950 520.050 442.050 ;
        RECT 511.950 436.950 514.050 439.050 ;
        RECT 518.400 433.050 519.450 439.950 ;
        RECT 517.950 430.950 520.050 433.050 ;
        RECT 502.950 427.950 505.050 430.050 ;
        RECT 514.950 427.950 517.050 430.050 ;
        RECT 472.950 424.950 475.050 427.050 ;
        RECT 475.950 424.950 478.050 427.050 ;
        RECT 469.950 421.950 472.050 424.050 ;
        RECT 478.950 421.950 481.050 424.050 ;
        RECT 466.950 409.950 469.050 412.050 ;
        RECT 463.950 397.950 466.050 400.050 ;
        RECT 463.950 376.950 466.050 379.050 ;
        RECT 448.950 373.950 451.050 376.050 ;
        RECT 445.950 371.100 448.050 373.200 ;
        RECT 454.950 371.100 457.050 373.200 ;
        RECT 391.950 349.950 394.050 352.050 ;
        RECT 412.950 349.950 415.050 352.050 ;
        RECT 385.950 343.950 388.050 346.050 ;
        RECT 392.700 345.300 394.800 347.400 ;
        RECT 383.400 334.350 384.600 336.600 ;
        RECT 383.100 331.950 385.200 334.050 ;
        RECT 393.300 327.600 394.800 345.300 ;
        RECT 392.700 325.500 394.800 327.600 ;
        RECT 379.950 319.950 382.050 322.050 ;
        RECT 393.300 320.700 394.800 325.500 ;
        RECT 380.400 307.050 381.450 319.950 ;
        RECT 392.700 318.600 394.800 320.700 ;
        RECT 395.700 345.300 397.800 347.400 ;
        RECT 398.700 345.300 400.800 347.400 ;
        RECT 401.700 345.300 403.800 347.400 ;
        RECT 395.700 323.700 396.900 345.300 ;
        RECT 398.700 327.600 400.200 345.300 ;
        RECT 401.700 333.000 402.900 345.300 ;
        RECT 407.100 344.400 409.200 346.500 ;
        RECT 415.200 345.300 417.300 347.400 ;
        RECT 418.200 345.300 420.300 347.400 ;
        RECT 421.200 345.300 423.300 347.400 ;
        RECT 403.800 338.400 405.900 340.500 ;
        RECT 407.700 333.900 408.600 344.400 ;
        RECT 410.100 337.950 412.200 340.050 ;
        RECT 410.400 336.000 411.600 337.650 ;
        RECT 401.100 330.900 403.200 333.000 ;
        RECT 406.500 331.800 408.600 333.900 ;
        RECT 409.950 331.950 412.050 336.000 ;
        RECT 398.100 325.500 400.200 327.600 ;
        RECT 395.700 318.600 397.800 323.700 ;
        RECT 398.700 320.700 400.200 325.500 ;
        RECT 401.700 323.700 402.900 330.900 ;
        RECT 407.700 325.200 408.600 331.800 ;
        RECT 401.100 321.600 403.200 323.700 ;
        RECT 406.500 323.100 408.600 325.200 ;
        RECT 416.100 323.700 417.300 345.300 ;
        RECT 415.200 321.600 417.300 323.700 ;
        RECT 418.500 328.800 419.700 345.300 ;
        RECT 421.500 341.700 422.700 345.300 ;
        RECT 421.500 339.600 423.600 341.700 ;
        RECT 434.400 340.200 435.450 365.400 ;
        RECT 442.950 364.800 445.050 366.900 ;
        RECT 446.400 358.050 447.450 371.100 ;
        RECT 455.400 370.350 456.600 371.100 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 458.400 366.450 459.600 367.650 ;
        RECT 464.400 366.450 465.450 376.950 ;
        RECT 458.400 365.400 465.450 366.450 ;
        RECT 445.950 355.950 448.050 358.050 ;
        RECT 445.950 349.950 448.050 352.050 ;
        RECT 439.950 343.950 442.050 346.050 ;
        RECT 418.500 326.700 420.600 328.800 ;
        RECT 418.500 320.700 419.700 326.700 ;
        RECT 422.100 320.700 423.600 339.600 ;
        RECT 433.950 338.100 436.050 340.200 ;
        RECT 440.400 334.050 441.450 343.950 ;
        RECT 428.100 331.950 430.200 334.050 ;
        RECT 434.100 331.950 436.200 334.050 ;
        RECT 439.950 331.950 442.050 334.050 ;
        RECT 446.400 333.900 447.450 349.950 ;
        RECT 466.950 346.950 469.050 349.050 ;
        RECT 460.950 343.950 463.050 346.050 ;
        RECT 454.950 338.100 457.050 340.200 ;
        RECT 461.400 339.600 462.450 343.950 ;
        RECT 467.400 339.600 468.450 346.950 ;
        RECT 455.400 337.350 456.600 338.100 ;
        RECT 461.400 337.350 462.600 339.600 ;
        RECT 467.400 337.350 468.600 339.600 ;
        RECT 470.400 339.450 471.450 421.950 ;
        RECT 479.400 417.600 480.450 421.950 ;
        RECT 499.800 420.300 501.900 422.400 ;
        RECT 502.950 421.950 505.050 424.050 ;
        RECT 503.400 421.200 504.600 421.950 ;
        RECT 479.400 415.350 480.600 417.600 ;
        RECT 496.950 416.100 499.050 418.200 ;
        RECT 497.400 415.350 498.600 416.100 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 497.100 412.950 499.200 415.050 ;
        RECT 500.100 414.900 501.000 420.300 ;
        RECT 503.100 418.800 505.200 420.900 ;
        RECT 507.000 417.900 509.100 419.700 ;
        RECT 501.900 416.700 510.600 417.900 ;
        RECT 501.900 415.800 504.000 416.700 ;
        RECT 500.100 413.700 507.000 414.900 ;
        RECT 476.400 411.900 477.600 412.650 ;
        RECT 475.950 409.800 478.050 411.900 ;
        RECT 500.100 406.500 501.300 413.700 ;
        RECT 503.100 409.950 505.200 412.050 ;
        RECT 506.100 411.300 507.000 413.700 ;
        RECT 503.400 407.400 504.600 409.650 ;
        RECT 506.100 409.200 508.200 411.300 ;
        RECT 509.700 407.700 510.600 416.700 ;
        RECT 511.800 412.950 513.900 415.050 ;
        RECT 512.400 411.450 513.600 412.650 ;
        RECT 515.400 411.450 516.450 427.950 ;
        RECT 521.400 427.050 522.450 449.100 ;
        RECT 524.400 439.050 525.450 449.100 ;
        RECT 527.400 445.050 528.450 469.950 ;
        RECT 532.950 457.950 535.050 460.050 ;
        RECT 533.400 450.600 534.450 457.950 ;
        RECT 539.400 457.050 540.450 514.950 ;
        RECT 542.400 492.600 543.450 547.950 ;
        RECT 545.400 544.050 546.450 554.400 ;
        RECT 550.950 553.950 553.050 556.050 ;
        RECT 547.950 550.950 550.050 553.050 ;
        RECT 544.950 541.950 547.050 544.050 ;
        RECT 548.400 532.050 549.450 550.950 ;
        RECT 563.400 547.050 564.450 566.400 ;
        RECT 568.950 565.800 571.050 567.900 ;
        RECT 562.950 544.950 565.050 547.050 ;
        RECT 575.400 544.050 576.450 583.950 ;
        RECT 577.950 580.950 580.050 583.050 ;
        RECT 578.400 562.050 579.450 580.950 ;
        RECT 577.950 559.950 580.050 562.050 ;
        RECT 581.400 553.050 582.450 607.950 ;
        RECT 590.400 606.600 591.450 631.950 ;
        RECT 593.400 628.050 594.450 673.950 ;
        RECT 596.400 652.050 597.450 677.400 ;
        RECT 601.950 673.950 604.050 679.050 ;
        RECT 605.400 667.050 606.450 712.950 ;
        RECT 607.950 700.950 610.050 703.050 ;
        RECT 604.950 664.950 607.050 667.050 ;
        RECT 601.950 661.950 604.050 664.050 ;
        RECT 595.950 649.950 598.050 652.050 ;
        RECT 602.400 651.600 603.450 661.950 ;
        RECT 608.400 652.050 609.450 700.950 ;
        RECT 602.400 649.350 603.600 651.600 ;
        RECT 607.950 649.950 610.050 652.050 ;
        RECT 598.950 646.950 601.050 649.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 599.400 645.900 600.600 646.650 ;
        RECT 598.950 643.800 601.050 645.900 ;
        RECT 605.400 645.450 606.600 646.650 ;
        RECT 605.400 644.400 609.450 645.450 ;
        RECT 592.950 625.950 595.050 628.050 ;
        RECT 595.950 610.950 598.050 613.050 ;
        RECT 596.400 606.600 597.450 610.950 ;
        RECT 590.400 604.350 591.600 606.600 ;
        RECT 596.400 604.350 597.600 606.600 ;
        RECT 601.950 605.100 604.050 607.200 ;
        RECT 602.400 604.350 603.600 605.100 ;
        RECT 608.400 604.050 609.450 644.400 ;
        RECT 611.400 634.050 612.450 769.950 ;
        RECT 613.950 760.950 616.050 763.050 ;
        RECT 622.950 761.100 625.050 763.200 ;
        RECT 614.400 756.900 615.450 760.950 ;
        RECT 623.400 760.350 624.600 761.100 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 620.400 756.900 621.600 757.650 ;
        RECT 626.400 756.900 627.600 757.650 ;
        RECT 613.950 754.800 616.050 756.900 ;
        RECT 619.950 754.800 622.050 756.900 ;
        RECT 625.950 754.800 628.050 756.900 ;
        RECT 616.950 732.450 619.050 733.050 ;
        RECT 622.950 732.450 625.050 733.050 ;
        RECT 616.950 731.400 625.050 732.450 ;
        RECT 616.950 730.950 619.050 731.400 ;
        RECT 622.950 730.950 625.050 731.400 ;
        RECT 619.950 728.100 622.050 730.200 ;
        RECT 620.400 727.350 621.600 728.100 ;
        RECT 625.950 727.950 628.050 730.050 ;
        RECT 614.100 724.950 616.200 727.050 ;
        RECT 619.500 724.950 621.600 727.050 ;
        RECT 622.800 724.950 624.900 727.050 ;
        RECT 614.400 722.400 615.600 724.650 ;
        RECT 623.400 722.400 624.600 724.650 ;
        RECT 614.400 712.050 615.450 722.400 ;
        RECT 623.400 712.050 624.450 722.400 ;
        RECT 613.950 709.950 616.050 712.050 ;
        RECT 622.950 709.950 625.050 712.050 ;
        RECT 619.950 691.950 622.050 694.050 ;
        RECT 613.950 682.950 616.050 688.050 ;
        RECT 620.400 684.600 621.450 691.950 ;
        RECT 626.400 688.050 627.450 727.950 ;
        RECT 632.400 715.050 633.450 775.950 ;
        RECT 635.400 756.900 636.450 781.950 ;
        RECT 638.400 769.050 639.450 820.950 ;
        RECT 643.950 814.950 646.050 817.050 ;
        RECT 644.400 801.900 645.450 814.950 ;
        RECT 652.950 807.000 655.050 811.050 ;
        RECT 653.400 805.350 654.600 807.000 ;
        RECT 668.400 805.050 669.450 826.950 ;
        RECT 670.950 817.950 673.050 820.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 655.950 802.950 658.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 643.950 799.800 646.050 801.900 ;
        RECT 650.400 800.400 651.600 802.650 ;
        RECT 656.400 801.900 657.600 802.650 ;
        RECT 650.400 796.050 651.450 800.400 ;
        RECT 655.950 799.800 658.050 801.900 ;
        RECT 649.950 793.950 652.050 796.050 ;
        RECT 671.400 778.050 672.450 817.950 ;
        RECT 674.400 814.050 675.450 839.100 ;
        RECT 680.400 834.450 681.450 865.950 ;
        RECT 686.400 841.200 687.450 874.950 ;
        RECT 688.950 871.950 691.050 874.050 ;
        RECT 689.400 844.050 690.450 871.950 ;
        RECT 692.400 862.050 693.450 886.950 ;
        RECT 691.950 859.950 694.050 862.050 ;
        RECT 688.950 841.950 691.050 844.050 ;
        RECT 685.950 839.100 688.050 841.200 ;
        RECT 691.950 840.000 694.050 844.050 ;
        RECT 695.400 840.450 696.450 889.950 ;
        RECT 698.400 877.050 699.450 896.400 ;
        RECT 700.950 895.950 703.050 896.400 ;
        RECT 704.400 892.050 705.450 898.950 ;
        RECT 707.400 892.050 708.450 925.950 ;
        RECT 722.400 925.050 723.450 931.950 ;
        RECT 715.950 922.800 718.050 924.900 ;
        RECT 721.950 922.950 724.050 925.050 ;
        RECT 716.400 918.600 717.450 922.800 ;
        RECT 724.950 919.950 727.050 922.050 ;
        RECT 716.400 916.350 717.600 918.600 ;
        RECT 712.950 913.950 715.050 916.050 ;
        RECT 715.950 913.950 718.050 916.050 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 713.400 911.400 714.600 913.650 ;
        RECT 719.400 912.900 720.600 913.650 ;
        RECT 725.400 912.900 726.450 919.950 ;
        RECT 713.400 909.450 714.450 911.400 ;
        RECT 718.950 910.800 721.050 912.900 ;
        RECT 724.950 910.800 727.050 912.900 ;
        RECT 713.400 908.400 717.450 909.450 ;
        RECT 703.950 889.950 706.050 892.050 ;
        RECT 706.950 889.950 709.050 892.050 ;
        RECT 707.400 888.450 708.450 889.950 ;
        RECT 707.400 887.400 711.450 888.450 ;
        RECT 703.950 884.100 706.050 886.200 ;
        RECT 710.400 885.600 711.450 887.400 ;
        RECT 704.400 883.350 705.600 884.100 ;
        RECT 710.400 883.350 711.600 885.600 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 700.950 877.950 703.050 880.050 ;
        RECT 707.400 879.900 708.600 880.650 ;
        RECT 716.400 880.050 717.450 908.400 ;
        RECT 721.950 904.950 724.050 907.050 ;
        RECT 697.950 874.950 700.050 877.050 ;
        RECT 701.400 868.050 702.450 877.950 ;
        RECT 706.950 877.800 709.050 879.900 ;
        RECT 712.950 877.950 715.050 880.050 ;
        RECT 715.950 877.950 718.050 880.050 ;
        RECT 703.950 874.950 706.050 877.050 ;
        RECT 713.400 871.050 714.450 877.950 ;
        RECT 712.950 868.950 715.050 871.050 ;
        RECT 700.950 865.950 703.050 868.050 ;
        RECT 703.950 859.950 706.050 862.050 ;
        RECT 700.950 841.950 703.050 844.050 ;
        RECT 686.400 838.350 687.600 839.100 ;
        RECT 692.400 838.350 693.600 840.000 ;
        RECT 695.400 839.400 699.450 840.450 ;
        RECT 685.950 835.950 688.050 838.050 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 689.400 834.900 690.600 835.650 ;
        RECT 680.400 833.400 684.450 834.450 ;
        RECT 673.950 811.950 676.050 814.050 ;
        RECT 683.400 811.050 684.450 833.400 ;
        RECT 688.950 832.800 691.050 834.900 ;
        RECT 691.950 829.950 694.050 832.050 ;
        RECT 685.950 820.950 688.050 823.050 ;
        RECT 682.950 808.950 685.050 811.050 ;
        RECT 679.950 806.100 682.050 808.200 ;
        RECT 680.400 805.350 681.600 806.100 ;
        RECT 674.100 802.950 676.200 805.050 ;
        RECT 679.500 802.950 681.600 805.050 ;
        RECT 682.800 802.950 684.900 805.050 ;
        RECT 674.400 800.400 675.600 802.650 ;
        RECT 683.400 801.450 684.600 802.650 ;
        RECT 686.400 801.450 687.450 820.950 ;
        RECT 688.950 806.100 691.050 808.200 ;
        RECT 689.400 802.050 690.450 806.100 ;
        RECT 683.400 800.400 687.450 801.450 ;
        RECT 674.400 796.050 675.450 800.400 ;
        RECT 688.950 799.950 691.050 802.050 ;
        RECT 673.950 793.950 676.050 796.050 ;
        RECT 670.950 775.950 673.050 778.050 ;
        RECT 637.950 766.950 640.050 769.050 ;
        RECT 646.950 761.100 649.050 763.200 ;
        RECT 652.950 761.100 655.050 763.200 ;
        RECT 671.400 762.600 672.450 775.950 ;
        RECT 688.950 772.950 691.050 775.050 ;
        RECT 676.950 769.950 679.050 772.050 ;
        RECT 685.950 769.950 688.050 772.050 ;
        RECT 677.400 762.600 678.450 769.950 ;
        RECT 682.950 763.950 685.050 766.050 ;
        RECT 647.400 760.350 648.600 761.100 ;
        RECT 653.400 760.350 654.600 761.100 ;
        RECT 671.400 760.350 672.600 762.600 ;
        RECT 677.400 760.350 678.600 762.600 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 646.950 757.950 649.050 760.050 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 652.950 757.950 655.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 634.950 754.800 637.050 756.900 ;
        RECT 638.400 751.050 639.450 757.950 ;
        RECT 644.400 755.400 645.600 757.650 ;
        RECT 650.400 756.900 651.600 757.650 ;
        RECT 674.400 756.900 675.600 757.650 ;
        RECT 637.950 748.950 640.050 751.050 ;
        RECT 644.400 739.050 645.450 755.400 ;
        RECT 649.950 754.800 652.050 756.900 ;
        RECT 673.950 754.800 676.050 756.900 ;
        RECT 670.950 751.950 673.050 754.050 ;
        RECT 667.950 748.950 670.050 751.050 ;
        RECT 661.950 745.950 664.050 748.050 ;
        RECT 662.400 742.050 663.450 745.950 ;
        RECT 661.950 739.950 664.050 742.050 ;
        RECT 643.950 736.950 646.050 739.050 ;
        RECT 640.950 733.050 643.050 733.200 ;
        RECT 643.950 733.050 646.050 733.200 ;
        RECT 640.950 731.100 646.050 733.050 ;
        RECT 642.000 730.950 645.000 731.100 ;
        RECT 640.950 727.950 643.050 730.050 ;
        RECT 646.950 728.100 649.050 730.200 ;
        RECT 653.400 729.450 654.600 729.600 ;
        RECT 653.400 728.400 660.450 729.450 ;
        RECT 641.400 727.350 642.600 727.950 ;
        RECT 647.400 727.350 648.600 728.100 ;
        RECT 653.400 727.350 654.600 728.400 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 649.950 724.950 652.050 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 634.950 721.950 637.050 724.050 ;
        RECT 644.400 722.400 645.600 724.650 ;
        RECT 650.400 723.900 651.600 724.650 ;
        RECT 631.950 712.950 634.050 715.050 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 620.400 682.350 621.600 684.600 ;
        RECT 625.950 684.000 628.050 688.050 ;
        RECT 629.400 685.050 630.450 697.950 ;
        RECT 631.950 688.950 634.050 691.050 ;
        RECT 626.400 682.350 627.600 684.000 ;
        RECT 628.950 682.950 631.050 685.050 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 619.950 679.950 622.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 617.400 678.900 618.600 679.650 ;
        RECT 623.400 678.900 624.600 679.650 ;
        RECT 616.950 676.800 619.050 678.900 ;
        RECT 622.950 676.800 625.050 678.900 ;
        RECT 628.950 667.950 631.050 670.050 ;
        RECT 622.950 664.950 625.050 667.050 ;
        RECT 616.950 658.950 619.050 661.050 ;
        RECT 613.950 655.950 616.050 658.050 ;
        RECT 610.950 631.950 613.050 634.050 ;
        RECT 610.950 625.950 613.050 628.050 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 593.400 599.400 594.600 601.650 ;
        RECT 599.400 600.000 600.600 601.650 ;
        RECT 593.400 592.050 594.450 599.400 ;
        RECT 598.950 595.950 601.050 600.000 ;
        RECT 592.950 589.950 595.050 592.050 ;
        RECT 601.950 586.950 604.050 589.050 ;
        RECT 586.950 580.950 589.050 583.050 ;
        RECT 587.400 573.600 588.450 580.950 ;
        RECT 587.400 571.350 588.600 573.600 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 590.400 566.400 591.600 568.650 ;
        RECT 580.950 550.950 583.050 553.050 ;
        RECT 590.400 550.050 591.450 566.400 ;
        RECT 589.950 547.950 592.050 550.050 ;
        RECT 554.700 540.300 556.800 542.400 ;
        RECT 555.300 535.500 556.800 540.300 ;
        RECT 554.700 533.400 556.800 535.500 ;
        RECT 547.950 529.950 550.050 532.050 ;
        RECT 545.100 526.950 547.200 529.050 ;
        RECT 545.400 525.450 546.600 526.650 ;
        RECT 545.400 524.400 549.450 525.450 ;
        RECT 544.950 499.950 547.050 502.050 ;
        RECT 545.400 496.050 546.450 499.950 ;
        RECT 544.950 493.950 547.050 496.050 ;
        RECT 542.400 490.350 543.600 492.600 ;
        RECT 548.400 492.450 549.450 524.400 ;
        RECT 550.950 524.100 553.050 526.200 ;
        RECT 551.400 502.050 552.450 524.100 ;
        RECT 555.300 515.700 556.800 533.400 ;
        RECT 554.700 513.600 556.800 515.700 ;
        RECT 557.700 537.300 559.800 542.400 ;
        RECT 560.700 540.300 562.800 542.400 ;
        RECT 574.950 541.950 577.050 544.050 ;
        RECT 579.600 540.300 581.700 542.400 ;
        RECT 582.600 540.300 585.600 542.400 ;
        RECT 586.950 541.950 589.050 544.050 ;
        RECT 557.700 515.700 558.900 537.300 ;
        RECT 560.700 535.500 562.200 540.300 ;
        RECT 563.100 537.300 565.200 539.400 ;
        RECT 560.100 533.400 562.200 535.500 ;
        RECT 560.700 515.700 562.200 533.400 ;
        RECT 563.700 530.100 564.900 537.300 ;
        RECT 568.500 535.800 570.600 537.900 ;
        RECT 577.200 537.300 579.300 539.400 ;
        RECT 563.100 528.000 565.200 530.100 ;
        RECT 569.700 529.200 570.600 535.800 ;
        RECT 563.700 515.700 564.900 528.000 ;
        RECT 568.500 527.100 570.600 529.200 ;
        RECT 565.800 520.500 567.900 522.600 ;
        RECT 569.700 516.600 570.600 527.100 ;
        RECT 571.950 524.100 574.050 526.200 ;
        RECT 572.400 523.350 573.600 524.100 ;
        RECT 572.100 520.950 574.200 523.050 ;
        RECT 557.700 513.600 559.800 515.700 ;
        RECT 560.700 513.600 562.800 515.700 ;
        RECT 563.700 513.600 565.800 515.700 ;
        RECT 569.100 514.500 571.200 516.600 ;
        RECT 578.100 515.700 579.300 537.300 ;
        RECT 580.500 534.300 581.700 540.300 ;
        RECT 580.500 532.200 582.600 534.300 ;
        RECT 580.500 515.700 581.700 532.200 ;
        RECT 584.100 521.400 585.600 540.300 ;
        RECT 583.500 519.300 585.600 521.400 ;
        RECT 583.500 515.700 584.700 519.300 ;
        RECT 577.200 513.600 579.300 515.700 ;
        RECT 580.200 513.600 582.300 515.700 ;
        RECT 583.200 513.600 585.300 515.700 ;
        RECT 587.400 508.050 588.450 541.950 ;
        RECT 602.400 534.450 603.450 586.950 ;
        RECT 607.950 580.950 610.050 583.050 ;
        RECT 608.400 573.600 609.450 580.950 ;
        RECT 611.400 577.050 612.450 625.950 ;
        RECT 614.400 625.050 615.450 655.950 ;
        RECT 617.400 637.050 618.450 658.950 ;
        RECT 623.400 651.600 624.450 664.950 ;
        RECT 629.400 651.600 630.450 667.950 ;
        RECT 632.400 664.050 633.450 688.950 ;
        RECT 635.400 685.200 636.450 721.950 ;
        RECT 644.400 720.450 645.450 722.400 ;
        RECT 649.950 721.800 652.050 723.900 ;
        RECT 655.950 721.950 658.050 724.050 ;
        RECT 641.400 719.400 645.450 720.450 ;
        RECT 641.400 700.050 642.450 719.400 ;
        RECT 649.950 718.650 652.050 720.750 ;
        RECT 643.950 715.950 646.050 718.050 ;
        RECT 640.950 697.950 643.050 700.050 ;
        RECT 637.950 694.950 640.050 697.050 ;
        RECT 634.950 683.100 637.050 685.200 ;
        RECT 631.950 661.950 634.050 664.050 ;
        RECT 635.400 652.050 636.450 683.100 ;
        RECT 623.400 649.350 624.600 651.600 ;
        RECT 629.400 649.350 630.600 651.600 ;
        RECT 634.950 649.950 637.050 652.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 626.400 645.900 627.600 646.650 ;
        RECT 616.950 634.950 619.050 637.050 ;
        RECT 613.950 622.950 616.050 625.050 ;
        RECT 613.950 616.950 616.050 619.050 ;
        RECT 614.400 601.050 615.450 616.950 ;
        RECT 620.400 616.050 621.450 643.950 ;
        RECT 625.950 643.800 628.050 645.900 ;
        RECT 632.400 644.400 633.600 646.650 ;
        RECT 632.400 637.050 633.450 644.400 ;
        RECT 631.950 634.950 634.050 637.050 ;
        RECT 628.950 622.950 631.050 625.050 ;
        RECT 619.950 613.950 622.050 616.050 ;
        RECT 619.950 606.000 622.050 610.050 ;
        RECT 620.400 604.350 621.600 606.000 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 613.950 598.950 616.050 601.050 ;
        RECT 623.400 600.900 624.600 601.650 ;
        RECT 622.950 598.800 625.050 600.900 ;
        RECT 610.950 574.950 613.050 577.050 ;
        RECT 608.400 571.350 609.600 573.600 ;
        RECT 613.950 572.100 616.050 574.200 ;
        RECT 620.400 573.450 621.600 573.600 ;
        RECT 623.400 573.450 624.450 598.800 ;
        RECT 620.400 572.400 627.450 573.450 ;
        RECT 614.400 571.350 615.600 572.100 ;
        RECT 620.400 571.350 621.600 572.400 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 619.950 568.950 622.050 571.050 ;
        RECT 611.400 566.400 612.600 568.650 ;
        RECT 617.400 567.900 618.600 568.650 ;
        RECT 611.400 556.050 612.450 566.400 ;
        RECT 616.950 565.800 619.050 567.900 ;
        RECT 617.400 564.450 618.450 565.800 ;
        RECT 614.400 563.400 618.450 564.450 ;
        RECT 610.950 553.950 613.050 556.050 ;
        RECT 610.950 541.950 613.050 544.050 ;
        RECT 602.400 533.400 606.450 534.450 ;
        RECT 595.950 530.100 598.050 532.200 ;
        RECT 601.950 530.100 604.050 532.200 ;
        RECT 596.400 529.350 597.600 530.100 ;
        RECT 590.100 526.950 592.200 529.050 ;
        RECT 596.100 526.950 598.200 529.050 ;
        RECT 586.950 505.950 589.050 508.050 ;
        RECT 598.950 505.950 601.050 508.050 ;
        RECT 550.950 499.950 553.050 502.050 ;
        RECT 560.700 501.300 562.800 503.400 ;
        RECT 556.950 493.950 559.050 496.050 ;
        RECT 551.400 492.450 552.600 492.600 ;
        RECT 548.400 491.400 552.600 492.450 ;
        RECT 542.100 487.950 544.200 490.050 ;
        RECT 544.950 484.950 547.050 487.050 ;
        RECT 541.950 481.950 544.050 484.050 ;
        RECT 542.400 460.050 543.450 481.950 ;
        RECT 545.400 468.450 546.450 484.950 ;
        RECT 548.400 472.050 549.450 491.400 ;
        RECT 551.400 490.350 552.600 491.400 ;
        RECT 557.400 490.050 558.450 493.950 ;
        RECT 551.100 487.950 553.200 490.050 ;
        RECT 556.950 487.950 559.050 490.050 ;
        RECT 561.300 483.600 562.800 501.300 ;
        RECT 560.700 481.500 562.800 483.600 ;
        RECT 561.300 476.700 562.800 481.500 ;
        RECT 560.700 474.600 562.800 476.700 ;
        RECT 563.700 501.300 565.800 503.400 ;
        RECT 566.700 501.300 568.800 503.400 ;
        RECT 569.700 501.300 571.800 503.400 ;
        RECT 563.700 479.700 564.900 501.300 ;
        RECT 566.700 483.600 568.200 501.300 ;
        RECT 569.700 489.000 570.900 501.300 ;
        RECT 575.100 500.400 577.200 502.500 ;
        RECT 583.200 501.300 585.300 503.400 ;
        RECT 586.200 501.300 588.300 503.400 ;
        RECT 589.200 501.300 591.300 503.400 ;
        RECT 571.800 494.400 573.900 496.500 ;
        RECT 575.700 489.900 576.600 500.400 ;
        RECT 578.100 493.950 580.200 496.050 ;
        RECT 578.400 492.000 579.600 493.650 ;
        RECT 569.100 486.900 571.200 489.000 ;
        RECT 574.500 487.800 576.600 489.900 ;
        RECT 577.950 487.950 580.050 492.000 ;
        RECT 580.950 490.950 583.050 493.050 ;
        RECT 566.100 481.500 568.200 483.600 ;
        RECT 563.700 474.600 565.800 479.700 ;
        RECT 566.700 476.700 568.200 481.500 ;
        RECT 569.700 479.700 570.900 486.900 ;
        RECT 575.700 481.200 576.600 487.800 ;
        RECT 581.400 483.450 582.450 490.950 ;
        RECT 569.100 477.600 571.200 479.700 ;
        RECT 574.500 479.100 576.600 481.200 ;
        RECT 578.400 482.400 582.450 483.450 ;
        RECT 566.700 474.600 568.800 476.700 ;
        RECT 547.950 469.950 550.050 472.050 ;
        RECT 545.400 467.400 549.450 468.450 ;
        RECT 541.950 457.950 544.050 460.050 ;
        RECT 538.950 454.950 541.050 457.050 ;
        RECT 533.400 448.350 534.600 450.600 ;
        RECT 538.950 449.100 541.050 451.200 ;
        RECT 539.400 448.350 540.600 449.100 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 535.950 445.950 538.050 448.050 ;
        RECT 538.950 445.950 541.050 448.050 ;
        RECT 541.950 445.950 544.050 448.050 ;
        RECT 526.950 442.950 529.050 445.050 ;
        RECT 536.400 443.400 537.600 445.650 ;
        RECT 542.400 444.900 543.600 445.650 ;
        RECT 548.400 445.050 549.450 467.400 ;
        RECT 553.950 454.950 556.050 457.050 ;
        RECT 536.400 439.050 537.450 443.400 ;
        RECT 541.950 442.800 544.050 444.900 ;
        RECT 547.950 442.950 550.050 445.050 ;
        RECT 554.400 441.450 555.450 454.950 ;
        RECT 559.950 449.100 562.050 451.200 ;
        RECT 565.950 449.100 568.050 451.200 ;
        RECT 574.950 449.100 577.050 451.200 ;
        RECT 560.400 448.350 561.600 449.100 ;
        RECT 566.400 448.350 567.600 449.100 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 562.950 445.950 565.050 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 563.400 443.400 564.600 445.650 ;
        RECT 569.400 444.450 570.600 445.650 ;
        RECT 569.400 443.400 573.450 444.450 ;
        RECT 551.400 440.400 555.450 441.450 ;
        RECT 523.950 436.950 526.050 439.050 ;
        RECT 535.950 436.950 538.050 439.050 ;
        RECT 544.950 427.950 547.050 430.050 ;
        RECT 520.950 424.950 523.050 427.050 ;
        RECT 535.950 424.950 538.050 427.050 ;
        RECT 521.400 418.200 522.450 424.950 ;
        RECT 520.950 416.100 523.050 418.200 ;
        RECT 529.950 416.100 532.050 418.200 ;
        RECT 536.400 417.600 537.450 424.950 ;
        RECT 530.400 415.350 531.600 416.100 ;
        RECT 536.400 415.350 537.600 417.600 ;
        RECT 541.950 416.100 544.050 418.200 ;
        RECT 529.950 412.950 532.050 415.050 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 512.400 410.400 516.450 411.450 ;
        RECT 499.800 404.400 501.900 406.500 ;
        RECT 509.400 405.600 511.500 407.700 ;
        RECT 508.950 388.950 511.050 391.050 ;
        RECT 475.950 371.100 478.050 373.200 ;
        RECT 481.950 371.100 484.050 373.200 ;
        RECT 499.950 371.100 502.050 373.200 ;
        RECT 476.400 370.350 477.600 371.100 ;
        RECT 482.400 370.350 483.600 371.100 ;
        RECT 500.400 370.350 501.600 371.100 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 479.400 365.400 480.600 367.650 ;
        RECT 503.400 366.900 504.600 367.650 ;
        RECT 509.400 366.900 510.450 388.950 ;
        RECT 475.950 355.950 478.050 358.050 ;
        RECT 470.400 338.400 474.450 339.450 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 463.950 334.950 466.050 337.050 ;
        RECT 466.950 334.950 469.050 337.050 ;
        RECT 458.400 333.900 459.600 334.650 ;
        RECT 445.950 331.800 448.050 333.900 ;
        RECT 457.950 331.800 460.050 333.900 ;
        RECT 464.400 332.400 465.600 334.650 ;
        RECT 434.400 330.000 435.600 331.650 ;
        RECT 433.950 325.950 436.050 330.000 ;
        RECT 451.950 325.950 454.050 328.050 ;
        RECT 442.950 322.950 445.050 325.050 ;
        RECT 398.700 318.600 400.800 320.700 ;
        RECT 417.600 318.600 419.700 320.700 ;
        RECT 420.600 318.600 423.600 320.700 ;
        RECT 379.950 304.950 382.050 307.050 ;
        RECT 427.950 304.950 430.050 307.050 ;
        RECT 361.950 298.950 364.050 301.050 ;
        RECT 409.950 298.950 412.050 301.050 ;
        RECT 424.950 298.950 427.050 301.050 ;
        RECT 346.950 292.950 349.050 295.050 ;
        RECT 352.950 293.100 355.050 295.200 ;
        RECT 347.400 286.050 348.450 292.950 ;
        RECT 353.400 292.350 354.600 293.100 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 356.400 287.400 357.600 289.650 ;
        RECT 346.950 283.950 349.050 286.050 ;
        RECT 356.400 280.050 357.450 287.400 ;
        RECT 362.400 280.050 363.450 298.950 ;
        RECT 367.950 292.950 370.050 295.050 ;
        RECT 376.950 293.100 379.050 295.200 ;
        RECT 368.400 280.050 369.450 292.950 ;
        RECT 377.400 292.350 378.600 293.100 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 376.950 289.950 379.050 292.050 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 374.400 288.000 375.600 289.650 ;
        RECT 380.400 289.050 381.600 289.650 ;
        RECT 373.950 285.450 376.050 288.000 ;
        RECT 380.400 287.400 385.050 289.050 ;
        RECT 394.950 288.450 397.050 292.050 ;
        RECT 400.800 289.950 402.900 292.050 ;
        RECT 381.000 286.950 385.050 287.400 ;
        RECT 392.400 287.400 397.050 288.450 ;
        RECT 373.950 284.400 378.450 285.450 ;
        RECT 373.950 283.950 376.050 284.400 ;
        RECT 355.950 277.950 358.050 280.050 ;
        RECT 361.950 277.950 364.050 280.050 ;
        RECT 367.950 277.950 370.050 280.050 ;
        RECT 343.950 274.950 346.050 277.050 ;
        RECT 344.700 267.300 346.800 269.400 ;
        RECT 345.300 249.600 346.800 267.300 ;
        RECT 344.700 247.500 346.800 249.600 ;
        RECT 345.300 242.700 346.800 247.500 ;
        RECT 344.700 240.600 346.800 242.700 ;
        RECT 347.700 267.300 349.800 269.400 ;
        RECT 350.700 267.300 352.800 269.400 ;
        RECT 353.700 267.300 355.800 269.400 ;
        RECT 347.700 245.700 348.900 267.300 ;
        RECT 350.700 249.600 352.200 267.300 ;
        RECT 353.700 255.000 354.900 267.300 ;
        RECT 359.100 266.400 361.200 268.500 ;
        RECT 367.200 267.300 369.300 269.400 ;
        RECT 370.200 267.300 372.300 269.400 ;
        RECT 373.200 267.300 375.300 269.400 ;
        RECT 355.800 260.400 357.900 262.500 ;
        RECT 359.700 255.900 360.600 266.400 ;
        RECT 362.100 259.950 364.200 262.050 ;
        RECT 362.400 258.900 363.600 259.650 ;
        RECT 361.950 256.800 364.050 258.900 ;
        RECT 353.100 252.900 355.200 255.000 ;
        RECT 358.500 253.800 360.600 255.900 ;
        RECT 350.100 247.500 352.200 249.600 ;
        RECT 347.700 240.600 349.800 245.700 ;
        RECT 350.700 242.700 352.200 247.500 ;
        RECT 353.700 245.700 354.900 252.900 ;
        RECT 359.700 247.200 360.600 253.800 ;
        RECT 353.100 243.600 355.200 245.700 ;
        RECT 358.500 245.100 360.600 247.200 ;
        RECT 368.100 245.700 369.300 267.300 ;
        RECT 367.200 243.600 369.300 245.700 ;
        RECT 370.500 250.800 371.700 267.300 ;
        RECT 373.500 263.700 374.700 267.300 ;
        RECT 373.500 261.600 375.600 263.700 ;
        RECT 370.500 248.700 372.600 250.800 ;
        RECT 370.500 242.700 371.700 248.700 ;
        RECT 374.100 242.700 375.600 261.600 ;
        RECT 350.700 240.600 352.800 242.700 ;
        RECT 369.600 240.600 371.700 242.700 ;
        RECT 372.600 240.600 375.600 242.700 ;
        RECT 340.950 235.950 343.050 238.050 ;
        RECT 352.950 235.950 355.050 238.050 ;
        RECT 340.950 215.100 343.050 217.200 ;
        RECT 348.000 216.600 352.050 217.050 ;
        RECT 341.400 214.350 342.600 215.100 ;
        RECT 347.400 214.950 352.050 216.600 ;
        RECT 347.400 214.350 348.600 214.950 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 346.950 211.950 349.050 214.050 ;
        RECT 337.950 208.950 340.050 211.050 ;
        RECT 344.400 210.900 345.600 211.650 ;
        RECT 353.400 211.050 354.450 235.950 ;
        RECT 377.400 229.050 378.450 284.400 ;
        RECT 382.950 277.950 385.050 280.050 ;
        RECT 383.400 258.900 384.450 277.950 ;
        RECT 382.950 256.800 385.050 258.900 ;
        RECT 380.100 253.950 382.200 256.050 ;
        RECT 386.100 253.950 388.200 256.050 ;
        RECT 382.950 250.950 385.050 253.050 ;
        RECT 386.400 251.400 387.600 253.650 ;
        RECT 364.950 226.950 367.050 229.050 ;
        RECT 376.950 226.950 379.050 229.050 ;
        RECT 358.950 220.950 361.050 223.050 ;
        RECT 355.950 215.100 358.050 217.200 ;
        RECT 334.950 205.950 337.050 208.050 ;
        RECT 338.400 202.050 339.450 208.950 ;
        RECT 343.950 208.800 346.050 210.900 ;
        RECT 352.950 208.950 355.050 211.050 ;
        RECT 340.950 205.950 343.050 208.050 ;
        RECT 337.950 199.950 340.050 202.050 ;
        RECT 334.950 187.950 337.050 190.050 ;
        RECT 331.950 184.950 334.050 187.050 ;
        RECT 323.400 181.350 324.600 182.100 ;
        RECT 329.400 181.350 330.600 183.600 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 320.400 177.900 321.600 178.650 ;
        RECT 326.400 177.900 327.600 178.650 ;
        RECT 335.400 177.900 336.450 187.950 ;
        RECT 337.950 181.950 340.050 184.050 ;
        RECT 319.950 175.800 322.050 177.900 ;
        RECT 325.950 175.800 328.050 177.900 ;
        RECT 334.950 175.800 337.050 177.900 ;
        RECT 311.400 173.400 315.450 174.450 ;
        RECT 301.950 169.950 304.050 172.050 ;
        RECT 289.950 166.950 292.050 169.050 ;
        RECT 283.950 151.950 286.050 154.050 ;
        RECT 283.950 137.100 286.050 139.200 ;
        RECT 290.400 138.600 291.450 166.950 ;
        RECT 301.950 163.800 304.050 165.900 ;
        RECT 298.950 154.950 301.050 157.050 ;
        RECT 284.400 136.350 285.600 137.100 ;
        RECT 290.400 136.350 291.600 138.600 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 277.950 130.950 280.050 133.050 ;
        RECT 287.400 132.900 288.600 133.650 ;
        RECT 286.950 130.800 289.050 132.900 ;
        RECT 283.950 124.950 286.050 127.050 ;
        RECT 277.950 118.950 280.050 121.050 ;
        RECT 274.950 115.950 277.050 118.050 ;
        RECT 275.400 106.050 276.450 115.950 ;
        RECT 266.400 103.350 267.600 105.600 ;
        RECT 272.400 103.350 273.600 105.600 ;
        RECT 274.950 103.950 277.050 106.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 263.400 99.900 264.600 100.650 ;
        RECT 262.950 97.800 265.050 99.900 ;
        RECT 269.400 99.000 270.600 100.650 ;
        RECT 278.400 99.900 279.450 118.950 ;
        RECT 284.400 100.050 285.450 124.950 ;
        RECT 299.400 118.050 300.450 154.950 ;
        RECT 302.400 127.050 303.450 163.800 ;
        RECT 311.400 138.600 312.450 173.400 ;
        RECT 338.400 172.050 339.450 181.950 ;
        RECT 337.950 169.950 340.050 172.050 ;
        RECT 319.950 142.950 322.050 145.050 ;
        RECT 311.400 136.350 312.600 138.600 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 308.400 132.000 309.600 133.650 ;
        RECT 307.950 127.950 310.050 132.000 ;
        RECT 314.400 131.400 315.600 133.650 ;
        RECT 301.950 124.950 304.050 127.050 ;
        RECT 308.400 121.050 309.450 127.950 ;
        RECT 314.400 124.050 315.450 131.400 ;
        RECT 313.950 121.950 316.050 124.050 ;
        RECT 307.950 118.950 310.050 121.050 ;
        RECT 320.400 118.050 321.450 142.950 ;
        RECT 325.950 137.100 328.050 139.200 ;
        RECT 334.950 137.100 337.050 139.200 ;
        RECT 341.400 138.600 342.450 205.950 ;
        RECT 356.400 195.450 357.450 215.100 ;
        RECT 359.400 199.050 360.450 220.950 ;
        RECT 365.400 216.600 366.450 226.950 ;
        RECT 377.400 223.050 378.450 226.950 ;
        RECT 370.950 220.950 373.050 223.050 ;
        RECT 376.950 220.950 379.050 223.050 ;
        RECT 371.400 216.600 372.450 220.950 ;
        RECT 365.400 214.350 366.600 216.600 ;
        RECT 371.400 214.350 372.600 216.600 ;
        RECT 377.100 214.950 379.200 217.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 377.400 212.400 378.600 214.650 ;
        RECT 383.400 213.450 384.450 250.950 ;
        RECT 386.400 223.050 387.450 251.400 ;
        RECT 385.950 220.950 388.050 223.050 ;
        RECT 386.100 214.950 388.200 217.050 ;
        RECT 386.400 213.450 387.600 214.650 ;
        RECT 383.400 212.400 387.600 213.450 ;
        RECT 361.950 208.950 364.050 211.050 ;
        RECT 368.400 210.900 369.600 211.650 ;
        RECT 367.950 208.800 370.050 210.900 ;
        RECT 377.400 210.450 378.450 212.400 ;
        RECT 374.400 209.400 378.450 210.450 ;
        RECT 358.950 196.950 361.050 199.050 ;
        RECT 374.400 196.050 375.450 209.400 ;
        RECT 382.950 199.950 385.050 202.050 ;
        RECT 356.400 194.400 360.450 195.450 ;
        RECT 355.950 190.950 358.050 193.050 ;
        RECT 356.400 184.200 357.450 190.950 ;
        RECT 349.950 182.100 352.050 184.200 ;
        RECT 355.950 182.100 358.050 184.200 ;
        RECT 359.400 184.050 360.450 194.400 ;
        RECT 367.950 193.950 370.050 196.050 ;
        RECT 373.950 193.950 376.050 196.050 ;
        RECT 350.400 181.350 351.600 182.100 ;
        RECT 356.400 181.350 357.600 182.100 ;
        RECT 358.950 181.950 361.050 184.050 ;
        RECT 361.950 182.100 364.050 184.200 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 347.400 176.400 348.600 178.650 ;
        RECT 353.400 177.900 354.600 178.650 ;
        RECT 347.400 166.050 348.450 176.400 ;
        RECT 352.950 175.800 355.050 177.900 ;
        RECT 358.950 175.950 361.050 178.050 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 359.400 160.050 360.450 175.950 ;
        RECT 346.950 157.950 349.050 160.050 ;
        RECT 358.950 157.950 361.050 160.050 ;
        RECT 326.400 124.050 327.450 137.100 ;
        RECT 335.400 136.350 336.600 137.100 ;
        RECT 341.400 136.350 342.600 138.600 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 332.400 131.400 333.600 133.650 ;
        RECT 338.400 132.900 339.600 133.650 ;
        RECT 347.400 133.050 348.450 157.950 ;
        RECT 362.400 154.050 363.450 182.100 ;
        RECT 368.400 166.050 369.450 193.950 ;
        RECT 376.950 190.950 379.050 193.050 ;
        RECT 377.400 187.050 378.450 190.950 ;
        RECT 376.950 183.000 379.050 187.050 ;
        RECT 377.400 181.350 378.600 183.000 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 374.400 176.400 375.600 178.650 ;
        RECT 374.400 175.050 375.450 176.400 ;
        RECT 383.400 175.050 384.450 199.950 ;
        RECT 374.400 173.400 379.050 175.050 ;
        RECT 375.000 172.950 379.050 173.400 ;
        RECT 382.950 172.950 385.050 175.050 ;
        RECT 386.400 172.050 387.450 212.400 ;
        RECT 392.400 183.450 393.450 287.400 ;
        RECT 394.950 286.950 397.050 287.400 ;
        RECT 410.400 268.050 411.450 298.950 ;
        RECT 419.400 294.450 420.600 294.600 ;
        RECT 419.400 293.400 423.450 294.450 ;
        RECT 419.400 292.350 420.600 293.400 ;
        RECT 418.800 289.950 420.900 292.050 ;
        RECT 422.400 277.050 423.450 293.400 ;
        RECT 425.400 292.050 426.450 298.950 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 428.400 286.050 429.450 304.950 ;
        RECT 443.400 301.050 444.450 322.950 ;
        RECT 442.950 298.950 445.050 301.050 ;
        RECT 443.400 294.600 444.450 298.950 ;
        RECT 452.400 298.200 453.450 325.950 ;
        RECT 464.400 325.050 465.450 332.400 ;
        RECT 463.950 322.950 466.050 325.050 ;
        RECT 464.400 319.050 465.450 322.950 ;
        RECT 463.950 316.950 466.050 319.050 ;
        RECT 473.400 316.050 474.450 338.400 ;
        RECT 476.400 333.900 477.450 355.950 ;
        RECT 479.400 340.200 480.450 365.400 ;
        RECT 502.950 364.800 505.050 366.900 ;
        RECT 508.950 364.800 511.050 366.900 ;
        RECT 515.400 355.050 516.450 410.400 ;
        RECT 533.400 410.400 534.600 412.650 ;
        RECT 533.400 379.050 534.450 410.400 ;
        RECT 542.400 406.050 543.450 416.100 ;
        RECT 541.950 403.950 544.050 406.050 ;
        RECT 532.950 376.950 535.050 379.050 ;
        RECT 520.950 371.100 523.050 373.200 ;
        RECT 526.950 371.100 529.050 373.200 ;
        RECT 533.400 373.050 534.450 376.950 ;
        RECT 521.400 370.350 522.600 371.100 ;
        RECT 527.400 370.350 528.600 371.100 ;
        RECT 532.950 370.950 535.050 373.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 524.400 366.900 525.600 367.650 ;
        RECT 530.400 366.900 531.600 367.650 ;
        RECT 523.950 364.800 526.050 366.900 ;
        RECT 529.950 364.800 532.050 366.900 ;
        RECT 526.950 361.950 529.050 364.050 ;
        RECT 514.950 352.950 517.050 355.050 ;
        RECT 520.950 352.950 523.050 355.050 ;
        RECT 478.950 338.100 481.050 340.200 ;
        RECT 484.950 338.100 487.050 343.050 ;
        RECT 490.950 338.100 493.050 340.200 ;
        RECT 485.400 337.350 486.600 338.100 ;
        RECT 491.400 337.350 492.600 338.100 ;
        RECT 505.950 337.950 508.050 340.050 ;
        RECT 514.950 339.000 517.050 343.050 ;
        RECT 521.400 339.600 522.450 352.950 ;
        RECT 527.400 343.050 528.450 361.950 ;
        RECT 545.400 349.050 546.450 427.950 ;
        RECT 551.400 420.450 552.450 440.400 ;
        RECT 559.950 439.950 562.050 442.050 ;
        RECT 548.400 419.400 552.450 420.450 ;
        RECT 548.400 388.050 549.450 419.400 ;
        RECT 553.950 417.000 556.050 421.050 ;
        RECT 560.400 418.200 561.450 439.950 ;
        RECT 563.400 439.050 564.450 443.400 ;
        RECT 562.950 436.950 565.050 439.050 ;
        RECT 572.400 433.050 573.450 443.400 ;
        RECT 575.400 442.050 576.450 449.100 ;
        RECT 574.950 439.950 577.050 442.050 ;
        RECT 571.950 430.950 574.050 433.050 ;
        RECT 568.950 424.950 571.050 427.050 ;
        RECT 565.950 418.950 568.050 421.050 ;
        RECT 554.400 415.350 555.600 417.000 ;
        RECT 559.950 416.100 562.050 418.200 ;
        RECT 560.400 415.350 561.600 416.100 ;
        RECT 553.950 412.950 556.050 415.050 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 557.400 410.400 558.600 412.650 ;
        RECT 557.400 391.050 558.450 410.400 ;
        RECT 566.400 403.050 567.450 418.950 ;
        RECT 569.400 409.050 570.450 424.950 ;
        RECT 572.400 424.050 573.450 430.950 ;
        RECT 578.400 430.050 579.450 482.400 ;
        RECT 584.100 479.700 585.300 501.300 ;
        RECT 583.200 477.600 585.300 479.700 ;
        RECT 586.500 484.800 587.700 501.300 ;
        RECT 589.500 497.700 590.700 501.300 ;
        RECT 589.500 495.600 591.600 497.700 ;
        RECT 586.500 482.700 588.600 484.800 ;
        RECT 586.500 476.700 587.700 482.700 ;
        RECT 590.100 476.700 591.600 495.600 ;
        RECT 599.400 493.050 600.450 505.950 ;
        RECT 602.400 495.450 603.450 530.100 ;
        RECT 605.400 499.050 606.450 533.400 ;
        RECT 611.400 529.050 612.450 541.950 ;
        RECT 610.950 526.950 613.050 529.050 ;
        RECT 610.950 520.950 613.050 523.050 ;
        RECT 607.950 517.950 610.050 520.050 ;
        RECT 608.400 499.050 609.450 517.950 ;
        RECT 611.400 514.050 612.450 520.950 ;
        RECT 614.400 514.050 615.450 563.400 ;
        RECT 616.950 556.950 619.050 559.050 ;
        RECT 617.400 541.050 618.450 556.950 ;
        RECT 626.400 547.050 627.450 572.400 ;
        RECT 625.950 544.950 628.050 547.050 ;
        RECT 616.950 538.950 619.050 541.050 ;
        RECT 629.400 538.050 630.450 622.950 ;
        RECT 638.400 621.450 639.450 694.950 ;
        RECT 644.400 691.050 645.450 715.950 ;
        RECT 650.400 700.050 651.450 718.650 ;
        RECT 656.400 718.050 657.450 721.950 ;
        RECT 655.950 715.950 658.050 718.050 ;
        RECT 652.950 706.950 658.050 709.050 ;
        RECT 655.950 703.800 658.050 705.900 ;
        RECT 649.950 697.950 652.050 700.050 ;
        RECT 643.950 688.950 646.050 691.050 ;
        RECT 643.950 683.100 646.050 685.200 ;
        RECT 649.950 684.000 652.050 688.050 ;
        RECT 644.400 682.350 645.600 683.100 ;
        RECT 650.400 682.350 651.600 684.000 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 647.400 678.900 648.600 679.650 ;
        RECT 646.950 676.800 649.050 678.900 ;
        RECT 656.400 673.050 657.450 703.800 ;
        RECT 659.400 700.050 660.450 728.400 ;
        RECT 662.400 718.050 663.450 739.950 ;
        RECT 664.950 736.950 667.050 739.050 ;
        RECT 661.950 715.950 664.050 718.050 ;
        RECT 661.950 712.800 664.050 714.900 ;
        RECT 662.400 703.050 663.450 712.800 ;
        RECT 665.400 706.050 666.450 736.950 ;
        RECT 668.400 730.050 669.450 748.950 ;
        RECT 671.400 742.050 672.450 751.950 ;
        RECT 670.950 739.950 673.050 742.050 ;
        RECT 667.950 727.950 670.050 730.050 ;
        RECT 673.950 728.100 676.050 730.200 ;
        RECT 674.400 727.350 675.600 728.100 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 671.400 723.900 672.600 724.650 ;
        RECT 670.950 718.950 673.050 723.900 ;
        RECT 677.400 722.400 678.600 724.650 ;
        RECT 677.400 718.050 678.450 722.400 ;
        RECT 676.950 715.950 679.050 718.050 ;
        RECT 670.950 712.950 673.050 715.050 ;
        RECT 671.400 709.050 672.450 712.950 ;
        RECT 667.950 706.950 670.050 709.050 ;
        RECT 670.950 706.950 673.050 709.050 ;
        RECT 664.950 703.950 667.050 706.050 ;
        RECT 668.400 703.050 669.450 706.950 ;
        RECT 661.950 700.950 664.050 703.050 ;
        RECT 667.950 700.950 670.050 703.050 ;
        RECT 658.950 697.950 661.050 700.050 ;
        RECT 661.950 697.800 664.050 699.900 ;
        RECT 664.950 697.950 667.050 700.050 ;
        RECT 658.950 685.950 661.050 688.050 ;
        RECT 659.400 678.900 660.450 685.950 ;
        RECT 658.950 676.800 661.050 678.900 ;
        RECT 655.950 670.950 658.050 673.050 ;
        RECT 643.950 664.950 646.050 667.050 ;
        RECT 640.950 649.950 643.050 652.050 ;
        RECT 641.400 622.050 642.450 649.950 ;
        RECT 644.400 646.050 645.450 664.950 ;
        RECT 652.950 650.100 655.050 652.200 ;
        RECT 659.400 651.450 660.600 651.600 ;
        RECT 662.400 651.450 663.450 697.800 ;
        RECT 665.400 691.050 666.450 697.950 ;
        RECT 677.400 697.050 678.450 715.950 ;
        RECT 679.950 709.950 682.050 712.050 ;
        RECT 676.950 694.950 679.050 697.050 ;
        RECT 664.950 685.950 667.050 691.050 ;
        RECT 667.950 684.000 670.050 688.050 ;
        RECT 673.950 684.000 676.050 688.050 ;
        RECT 680.400 685.050 681.450 709.950 ;
        RECT 668.400 682.350 669.600 684.000 ;
        RECT 674.400 682.350 675.600 684.000 ;
        RECT 679.950 682.950 682.050 685.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 671.400 677.400 672.600 679.650 ;
        RECT 677.400 678.900 678.600 679.650 ;
        RECT 667.950 670.950 670.050 673.050 ;
        RECT 659.400 650.400 663.450 651.450 ;
        RECT 653.400 649.350 654.600 650.100 ;
        RECT 659.400 649.350 660.600 650.400 ;
        RECT 664.950 650.100 667.050 652.200 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 658.950 646.950 661.050 649.050 ;
        RECT 643.950 643.950 646.050 646.050 ;
        RECT 650.400 645.900 651.600 646.650 ;
        RECT 649.950 643.800 652.050 645.900 ;
        RECT 656.400 645.000 657.600 646.650 ;
        RECT 665.400 646.050 666.450 650.100 ;
        RECT 643.950 640.800 646.050 642.900 ;
        RECT 655.950 640.950 658.050 645.000 ;
        RECT 664.950 643.950 667.050 646.050 ;
        RECT 635.400 620.400 639.450 621.450 ;
        RECT 631.950 613.950 634.050 616.050 ;
        RECT 628.950 535.950 631.050 538.050 ;
        RECT 632.400 537.450 633.450 613.950 ;
        RECT 635.400 583.050 636.450 620.400 ;
        RECT 640.950 619.950 643.050 622.050 ;
        RECT 641.400 610.050 642.450 619.950 ;
        RECT 640.950 607.950 643.050 610.050 ;
        RECT 644.400 606.600 645.450 640.800 ;
        RECT 646.950 637.950 649.050 640.050 ;
        RECT 647.400 619.050 648.450 637.950 ;
        RECT 658.950 622.950 661.050 625.050 ;
        RECT 646.950 616.950 649.050 619.050 ;
        RECT 652.950 607.950 655.050 610.050 ;
        RECT 644.400 604.350 645.600 606.600 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 641.400 600.900 642.600 601.650 ;
        RECT 640.950 598.800 643.050 600.900 ;
        RECT 647.400 600.000 648.600 601.650 ;
        RECT 653.400 601.050 654.450 607.950 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 646.950 595.950 649.050 600.000 ;
        RECT 652.950 598.950 655.050 601.050 ;
        RECT 652.950 595.800 655.050 597.900 ;
        RECT 637.950 586.950 640.050 589.050 ;
        RECT 634.950 580.950 637.050 583.050 ;
        RECT 638.400 573.600 639.450 586.950 ;
        RECT 638.400 571.350 639.600 573.600 ;
        RECT 643.950 572.100 646.050 574.200 ;
        RECT 644.400 571.350 645.600 572.100 ;
        RECT 637.950 568.950 640.050 571.050 ;
        RECT 640.950 568.950 643.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 641.400 567.900 642.600 568.650 ;
        RECT 640.950 565.800 643.050 567.900 ;
        RECT 647.400 566.400 648.600 568.650 ;
        RECT 647.400 559.050 648.450 566.400 ;
        RECT 653.400 565.050 654.450 595.800 ;
        RECT 656.400 589.050 657.450 601.950 ;
        RECT 655.950 586.950 658.050 589.050 ;
        RECT 655.950 572.100 658.050 574.200 ;
        RECT 656.400 568.050 657.450 572.100 ;
        RECT 659.400 571.050 660.450 622.950 ;
        RECT 664.950 613.950 667.050 616.050 ;
        RECT 665.400 607.200 666.450 613.950 ;
        RECT 668.400 610.050 669.450 670.950 ;
        RECT 671.400 670.050 672.450 677.400 ;
        RECT 676.950 676.800 679.050 678.900 ;
        RECT 679.950 676.950 682.050 679.050 ;
        RECT 680.400 670.050 681.450 676.950 ;
        RECT 670.950 667.950 673.050 670.050 ;
        RECT 679.950 667.950 682.050 670.050 ;
        RECT 683.400 667.050 684.450 763.950 ;
        RECT 686.400 756.900 687.450 769.950 ;
        RECT 685.950 754.800 688.050 756.900 ;
        RECT 685.950 730.950 688.050 733.050 ;
        RECT 686.400 688.050 687.450 730.950 ;
        RECT 689.400 696.450 690.450 772.950 ;
        RECT 692.400 763.050 693.450 829.950 ;
        RECT 698.400 807.450 699.450 839.400 ;
        RECT 701.400 826.050 702.450 841.950 ;
        RECT 704.400 832.050 705.450 859.950 ;
        RECT 712.950 847.950 715.050 850.050 ;
        RECT 713.400 840.600 714.450 847.950 ;
        RECT 718.950 844.950 721.050 847.050 ;
        RECT 715.950 841.950 718.050 844.050 ;
        RECT 719.400 841.050 720.450 844.950 ;
        RECT 713.400 838.350 714.600 840.600 ;
        RECT 718.950 838.950 721.050 841.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 710.400 834.900 711.600 835.650 ;
        RECT 716.400 834.900 717.600 835.650 ;
        RECT 722.400 834.900 723.450 904.950 ;
        RECT 725.400 886.050 726.450 910.800 ;
        RECT 728.400 901.050 729.450 931.950 ;
        RECT 731.400 912.900 732.450 956.400 ;
        RECT 739.950 952.950 742.050 957.000 ;
        RECT 749.400 955.050 750.450 962.100 ;
        RECT 761.400 961.350 762.600 962.100 ;
        RECT 767.400 961.350 768.600 962.100 ;
        RECT 760.950 958.950 763.050 961.050 ;
        RECT 763.950 958.950 766.050 961.050 ;
        RECT 766.950 958.950 769.050 961.050 ;
        RECT 764.400 957.900 765.600 958.650 ;
        RECT 763.950 955.800 766.050 957.900 ;
        RECT 748.950 952.950 751.050 955.050 ;
        RECT 739.950 946.950 742.050 949.050 ;
        RECT 740.400 922.050 741.450 946.950 ;
        RECT 739.950 918.000 742.050 922.050 ;
        RECT 749.400 919.200 750.450 952.950 ;
        RECT 766.950 925.950 769.050 928.050 ;
        RECT 740.400 916.350 741.600 918.000 ;
        RECT 748.950 917.100 751.050 919.200 ;
        RECT 760.950 917.100 763.050 919.200 ;
        RECT 767.400 918.600 768.450 925.950 ;
        RECT 736.950 913.950 739.050 916.050 ;
        RECT 739.950 913.950 742.050 916.050 ;
        RECT 737.400 912.900 738.600 913.650 ;
        RECT 730.950 910.800 733.050 912.900 ;
        RECT 736.950 910.800 739.050 912.900 ;
        RECT 731.400 907.050 732.450 910.800 ;
        RECT 730.950 904.950 733.050 907.050 ;
        RECT 730.950 901.800 733.050 903.900 ;
        RECT 727.800 898.950 729.900 901.050 ;
        RECT 724.950 883.950 727.050 886.050 ;
        RECT 731.400 885.600 732.450 901.800 ;
        RECT 749.400 895.050 750.450 917.100 ;
        RECT 761.400 916.350 762.600 917.100 ;
        RECT 767.400 916.350 768.600 918.600 ;
        RECT 757.950 913.950 760.050 916.050 ;
        RECT 760.950 913.950 763.050 916.050 ;
        RECT 763.950 913.950 766.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 758.400 912.000 759.600 913.650 ;
        RECT 757.950 907.950 760.050 912.000 ;
        RECT 764.400 911.400 765.600 913.650 ;
        RECT 764.400 907.050 765.450 911.400 ;
        RECT 773.400 910.050 774.450 962.100 ;
        RECT 775.950 958.950 778.050 961.050 ;
        RECT 776.400 943.050 777.450 958.950 ;
        RECT 779.400 958.050 780.450 962.100 ;
        RECT 788.400 961.350 789.600 962.100 ;
        RECT 794.400 961.350 795.600 962.100 ;
        RECT 818.400 961.350 819.600 962.100 ;
        RECT 826.950 961.950 829.050 964.050 ;
        RECT 784.950 958.950 787.050 961.050 ;
        RECT 787.950 958.950 790.050 961.050 ;
        RECT 790.950 958.950 793.050 961.050 ;
        RECT 793.950 958.950 796.050 961.050 ;
        RECT 796.950 958.950 799.050 961.050 ;
        RECT 815.100 958.950 817.200 961.050 ;
        RECT 818.400 958.950 820.500 961.050 ;
        RECT 823.800 958.950 825.900 961.050 ;
        RECT 778.950 955.950 781.050 958.050 ;
        RECT 785.400 956.400 786.600 958.650 ;
        RECT 791.400 956.400 792.600 958.650 ;
        RECT 797.400 957.900 798.600 958.650 ;
        RECT 815.400 957.900 816.600 958.650 ;
        RECT 824.400 957.900 825.600 958.650 ;
        RECT 785.400 949.050 786.450 956.400 ;
        RECT 784.950 946.950 787.050 949.050 ;
        RECT 791.400 946.050 792.450 956.400 ;
        RECT 796.950 955.800 799.050 957.900 ;
        RECT 814.950 955.800 817.050 957.900 ;
        RECT 823.950 955.800 826.050 957.900 ;
        RECT 815.400 952.050 816.450 955.800 ;
        RECT 814.950 949.950 817.050 952.050 ;
        RECT 790.950 943.950 793.050 946.050 ;
        RECT 824.400 943.050 825.450 955.800 ;
        RECT 775.950 940.950 778.050 943.050 ;
        RECT 796.950 940.950 799.050 943.050 ;
        RECT 823.950 940.950 826.050 943.050 ;
        RECT 778.950 931.950 781.050 934.050 ;
        RECT 784.950 931.950 787.050 934.050 ;
        RECT 775.950 922.950 778.050 925.050 ;
        RECT 772.950 907.950 775.050 910.050 ;
        RECT 763.950 904.950 766.050 907.050 ;
        RECT 739.950 892.950 742.050 895.050 ;
        RECT 748.950 892.950 751.050 895.050 ;
        RECT 731.400 883.350 732.600 885.600 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 724.950 877.950 727.050 880.050 ;
        RECT 728.400 878.400 729.600 880.650 ;
        RECT 734.400 878.400 735.600 880.650 ;
        RECT 725.400 835.050 726.450 877.950 ;
        RECT 728.400 871.050 729.450 878.400 ;
        RECT 727.950 868.950 730.050 871.050 ;
        RECT 734.400 862.050 735.450 878.400 ;
        RECT 740.400 868.050 741.450 892.950 ;
        RECT 751.950 891.450 754.050 895.050 ;
        RECT 749.400 891.000 754.050 891.450 ;
        RECT 749.400 890.400 753.450 891.000 ;
        RECT 742.950 883.950 745.050 886.050 ;
        RECT 749.400 885.450 750.450 890.400 ;
        RECT 769.950 889.950 772.050 892.050 ;
        RECT 746.400 884.400 750.450 885.450 ;
        RECT 751.950 885.000 754.050 889.050 ;
        RECT 739.950 865.950 742.050 868.050 ;
        RECT 733.950 859.950 736.050 862.050 ;
        RECT 743.400 850.050 744.450 883.950 ;
        RECT 746.400 877.050 747.450 884.400 ;
        RECT 752.400 883.350 753.600 885.000 ;
        RECT 757.950 884.100 760.050 886.200 ;
        RECT 766.950 884.100 769.050 886.200 ;
        RECT 758.400 883.350 759.600 884.100 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 755.400 879.900 756.600 880.650 ;
        RECT 754.950 877.800 757.050 879.900 ;
        RECT 761.400 878.400 762.600 880.650 ;
        RECT 745.950 874.950 748.050 877.050 ;
        RECT 755.400 871.050 756.450 877.800 ;
        RECT 761.400 871.050 762.450 878.400 ;
        RECT 754.950 868.950 757.050 871.050 ;
        RECT 760.950 868.950 763.050 871.050 ;
        RECT 751.950 865.950 754.050 868.050 ;
        RECT 742.950 847.950 745.050 850.050 ;
        RECT 727.950 844.950 730.050 847.050 ;
        RECT 709.950 832.800 712.050 834.900 ;
        RECT 715.950 832.800 718.050 834.900 ;
        RECT 721.950 832.800 724.050 834.900 ;
        RECT 724.950 832.950 727.050 835.050 ;
        RECT 703.950 829.950 706.050 832.050 ;
        RECT 722.400 826.050 723.450 832.800 ;
        RECT 724.950 829.800 727.050 831.900 ;
        RECT 700.950 823.950 703.050 826.050 ;
        RECT 721.950 823.950 724.050 826.050 ;
        RECT 703.950 814.950 706.050 817.050 ;
        RECT 695.400 806.400 699.450 807.450 ;
        RECT 704.400 807.600 705.450 814.950 ;
        RECT 718.950 808.950 721.050 811.050 ;
        RECT 695.400 766.050 696.450 806.400 ;
        RECT 704.400 805.350 705.600 807.600 ;
        RECT 709.950 806.100 712.050 808.200 ;
        RECT 715.950 806.100 718.050 808.200 ;
        RECT 710.400 805.350 711.600 806.100 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 701.400 801.900 702.600 802.650 ;
        RECT 700.950 799.800 703.050 801.900 ;
        RECT 707.400 801.000 708.600 802.650 ;
        RECT 701.400 796.050 702.450 799.800 ;
        RECT 706.950 796.950 709.050 801.000 ;
        RECT 700.950 793.950 703.050 796.050 ;
        RECT 709.950 793.950 712.050 796.050 ;
        RECT 716.400 795.450 717.450 806.100 ;
        RECT 719.400 799.050 720.450 808.950 ;
        RECT 718.950 796.950 721.050 799.050 ;
        RECT 713.400 794.400 717.450 795.450 ;
        RECT 697.950 781.950 700.050 784.050 ;
        RECT 694.950 763.950 697.050 766.050 ;
        RECT 691.950 760.950 694.050 763.050 ;
        RECT 698.400 762.600 699.450 781.950 ;
        RECT 703.950 775.950 706.050 778.050 ;
        RECT 704.400 763.050 705.450 775.950 ;
        RECT 706.950 766.950 709.050 769.050 ;
        RECT 698.400 760.350 699.600 762.600 ;
        RECT 703.950 760.950 706.050 763.050 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 695.400 756.900 696.600 757.650 ;
        RECT 701.400 757.050 702.600 757.650 ;
        RECT 694.950 754.800 697.050 756.900 ;
        RECT 701.400 755.400 706.050 757.050 ;
        RECT 702.000 754.950 706.050 755.400 ;
        RECT 703.950 742.950 706.050 745.050 ;
        RECT 704.400 736.050 705.450 742.950 ;
        RECT 703.950 733.950 706.050 736.050 ;
        RECT 694.950 728.100 697.050 730.200 ;
        RECT 700.950 729.000 703.050 733.050 ;
        RECT 695.400 727.350 696.600 728.100 ;
        RECT 701.400 727.350 702.600 729.000 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 698.400 722.400 699.600 724.650 ;
        RECT 694.950 715.950 697.050 718.050 ;
        RECT 689.400 695.400 693.450 696.450 ;
        RECT 688.950 691.950 691.050 694.050 ;
        RECT 685.950 685.950 688.050 688.050 ;
        RECT 686.400 682.050 687.450 685.950 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 689.400 679.050 690.450 691.950 ;
        RECT 692.400 685.050 693.450 695.400 ;
        RECT 695.400 691.050 696.450 715.950 ;
        RECT 698.400 712.050 699.450 722.400 ;
        RECT 697.950 709.950 700.050 712.050 ;
        RECT 707.400 694.050 708.450 766.950 ;
        RECT 710.400 724.050 711.450 793.950 ;
        RECT 713.400 778.050 714.450 794.400 ;
        RECT 718.950 793.800 721.050 795.900 ;
        RECT 712.950 775.950 715.050 778.050 ;
        RECT 713.400 748.050 714.450 775.950 ;
        RECT 719.400 775.050 720.450 793.800 ;
        RECT 722.400 775.050 723.450 823.950 ;
        RECT 725.400 792.450 726.450 829.800 ;
        RECT 728.400 820.050 729.450 844.950 ;
        RECT 730.950 838.950 733.050 844.050 ;
        RECT 742.950 839.100 745.050 841.200 ;
        RECT 752.400 840.600 753.450 865.950 ;
        RECT 754.950 859.950 757.050 862.050 ;
        RECT 743.400 838.350 744.600 839.100 ;
        RECT 752.400 838.350 753.600 840.600 ;
        RECT 736.800 835.950 738.900 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 751.500 835.950 753.600 838.050 ;
        RECT 733.950 832.950 736.050 835.050 ;
        RECT 737.400 834.900 738.600 835.650 ;
        RECT 734.400 826.050 735.450 832.950 ;
        RECT 736.950 832.800 739.050 834.900 ;
        RECT 746.400 833.400 747.600 835.650 ;
        RECT 746.400 828.450 747.450 833.400 ;
        RECT 748.950 829.950 751.050 832.050 ;
        RECT 746.400 827.400 750.450 828.450 ;
        RECT 733.950 823.950 736.050 826.050 ;
        RECT 742.950 823.950 745.050 826.050 ;
        RECT 727.950 817.950 730.050 820.050 ;
        RECT 734.400 807.600 735.450 823.950 ;
        RECT 739.950 814.950 742.050 817.050 ;
        RECT 734.400 805.350 735.600 807.600 ;
        RECT 728.100 802.950 730.200 805.050 ;
        RECT 733.500 802.950 735.600 805.050 ;
        RECT 736.800 802.950 738.900 805.050 ;
        RECT 728.400 801.900 729.600 802.650 ;
        RECT 737.400 801.900 738.600 802.650 ;
        RECT 727.950 799.800 730.050 801.900 ;
        RECT 736.950 799.800 739.050 801.900 ;
        RECT 728.400 796.050 729.450 799.800 ;
        RECT 727.950 793.950 730.050 796.050 ;
        RECT 725.400 791.400 729.450 792.450 ;
        RECT 718.800 772.950 720.900 775.050 ;
        RECT 721.950 772.950 724.050 775.050 ;
        RECT 719.400 762.600 720.450 772.950 ;
        RECT 719.400 760.350 720.600 762.600 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 722.400 756.900 723.600 757.650 ;
        RECT 721.950 754.800 724.050 756.900 ;
        RECT 715.950 751.950 718.050 754.050 ;
        RECT 712.950 745.950 715.050 748.050 ;
        RECT 716.400 729.450 717.450 751.950 ;
        RECT 722.400 745.050 723.450 754.800 ;
        RECT 721.950 742.950 724.050 745.050 ;
        RECT 728.400 739.050 729.450 791.400 ;
        RECT 736.950 790.950 739.050 793.050 ;
        RECT 730.950 781.950 733.050 784.050 ;
        RECT 727.950 736.950 730.050 739.050 ;
        RECT 713.400 728.400 717.450 729.450 ;
        RECT 721.950 729.000 724.050 733.050 ;
        RECT 709.950 721.950 712.050 724.050 ;
        RECT 706.950 691.950 709.050 694.050 ;
        RECT 694.950 688.950 697.050 691.050 ;
        RECT 703.950 688.950 706.050 691.050 ;
        RECT 709.950 688.950 712.050 691.050 ;
        RECT 691.950 682.950 694.050 685.050 ;
        RECT 697.950 684.000 700.050 688.050 ;
        RECT 704.400 685.200 705.450 688.950 ;
        RECT 698.400 682.350 699.600 684.000 ;
        RECT 703.950 683.100 706.050 685.200 ;
        RECT 704.400 682.350 705.600 683.100 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 688.950 676.950 691.050 679.050 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 695.400 678.900 696.600 679.650 ;
        RECT 701.400 678.900 702.600 679.650 ;
        RECT 685.950 670.950 688.050 673.050 ;
        RECT 682.950 664.950 685.050 667.050 ;
        RECT 679.950 661.050 682.050 664.050 ;
        RECT 676.950 658.950 679.050 661.050 ;
        RECT 679.950 660.000 685.050 661.050 ;
        RECT 680.400 659.400 685.050 660.000 ;
        RECT 681.000 658.950 685.050 659.400 ;
        RECT 677.400 651.600 678.450 658.950 ;
        RECT 679.950 654.450 682.050 655.050 ;
        RECT 686.400 654.450 687.450 670.950 ;
        RECT 679.950 653.400 687.450 654.450 ;
        RECT 679.950 652.950 682.050 653.400 ;
        RECT 677.400 649.350 678.600 651.600 ;
        RECT 682.950 650.100 685.050 652.200 ;
        RECT 688.950 650.100 691.050 652.200 ;
        RECT 683.400 649.350 684.600 650.100 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 680.400 645.900 681.600 646.650 ;
        RECT 679.950 643.800 682.050 645.900 ;
        RECT 689.400 640.050 690.450 650.100 ;
        RECT 688.950 637.950 691.050 640.050 ;
        RECT 679.950 625.950 682.050 628.050 ;
        RECT 676.950 622.950 679.050 625.050 ;
        RECT 667.950 607.950 670.050 610.050 ;
        RECT 664.950 605.100 667.050 607.200 ;
        RECT 670.950 605.100 673.050 607.200 ;
        RECT 677.400 606.600 678.450 622.950 ;
        RECT 680.400 607.050 681.450 625.950 ;
        RECT 692.400 615.450 693.450 676.950 ;
        RECT 694.950 676.800 697.050 678.900 ;
        RECT 700.950 676.800 703.050 678.900 ;
        RECT 694.950 673.650 697.050 675.750 ;
        RECT 695.400 643.050 696.450 673.650 ;
        RECT 710.400 670.050 711.450 688.950 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 703.950 650.100 706.050 652.200 ;
        RECT 704.400 649.350 705.600 650.100 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 706.950 646.950 709.050 649.050 ;
        RECT 697.950 643.950 700.050 646.050 ;
        RECT 701.400 645.000 702.600 646.650 ;
        RECT 707.400 645.000 708.600 646.650 ;
        RECT 694.950 640.950 697.050 643.050 ;
        RECT 698.400 631.050 699.450 643.950 ;
        RECT 700.950 640.950 703.050 645.000 ;
        RECT 706.950 640.950 709.050 645.000 ;
        RECT 713.400 640.050 714.450 728.400 ;
        RECT 722.400 727.350 723.600 729.000 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 719.400 723.900 720.600 724.650 ;
        RECT 725.400 724.050 726.600 724.650 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 725.400 721.950 730.050 724.050 ;
        RECT 718.950 718.650 721.050 720.750 ;
        RECT 719.400 709.050 720.450 718.650 ;
        RECT 718.950 706.950 721.050 709.050 ;
        RECT 715.950 691.950 718.050 694.050 ;
        RECT 718.950 691.950 721.050 694.050 ;
        RECT 709.950 637.950 712.050 640.050 ;
        RECT 712.950 637.950 715.050 640.050 ;
        RECT 706.950 634.950 709.050 637.050 ;
        RECT 697.950 628.950 700.050 631.050 ;
        RECT 689.400 614.400 693.450 615.450 ;
        RECT 685.950 607.950 688.050 610.050 ;
        RECT 665.400 604.350 666.600 605.100 ;
        RECT 671.400 604.350 672.600 605.100 ;
        RECT 677.400 604.350 678.600 606.600 ;
        RECT 679.950 604.950 682.050 607.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 668.400 599.400 669.600 601.650 ;
        RECT 674.400 600.000 675.600 601.650 ;
        RECT 668.400 595.050 669.450 599.400 ;
        RECT 673.950 595.950 676.050 600.000 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 667.950 592.950 670.050 595.050 ;
        RECT 674.400 592.050 675.450 595.950 ;
        RECT 676.950 592.950 679.050 598.050 ;
        RECT 673.950 589.950 676.050 592.050 ;
        RECT 679.950 589.950 682.050 592.050 ;
        RECT 673.950 583.950 676.050 586.050 ;
        RECT 667.950 577.950 670.050 580.050 ;
        RECT 668.400 573.600 669.450 577.950 ;
        RECT 674.400 573.600 675.450 583.950 ;
        RECT 680.400 577.050 681.450 589.950 ;
        RECT 679.950 574.950 682.050 577.050 ;
        RECT 668.400 571.350 669.600 573.600 ;
        RECT 674.400 571.350 675.600 573.600 ;
        RECT 658.950 568.950 661.050 571.050 ;
        RECT 664.950 568.950 667.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 655.950 565.950 658.050 568.050 ;
        RECT 665.400 566.400 666.600 568.650 ;
        RECT 671.400 567.900 672.600 568.650 ;
        RECT 677.400 567.900 678.600 568.650 ;
        RECT 683.400 567.900 684.450 601.950 ;
        RECT 652.950 562.950 655.050 565.050 ;
        RECT 655.950 562.800 658.050 564.900 ;
        RECT 649.950 559.950 652.050 562.050 ;
        RECT 646.950 556.950 649.050 559.050 ;
        RECT 650.400 550.050 651.450 559.950 ;
        RECT 649.950 547.950 652.050 550.050 ;
        RECT 637.950 544.950 640.050 547.050 ;
        RECT 632.400 536.400 636.450 537.450 ;
        RECT 619.800 532.500 621.900 534.600 ;
        RECT 617.100 523.950 619.200 526.050 ;
        RECT 620.100 525.300 621.300 532.500 ;
        RECT 623.400 529.350 624.600 531.600 ;
        RECT 629.400 531.300 631.500 533.400 ;
        RECT 623.100 526.950 625.200 529.050 ;
        RECT 626.100 527.700 628.200 529.800 ;
        RECT 626.100 525.300 627.000 527.700 ;
        RECT 620.100 524.100 627.000 525.300 ;
        RECT 617.400 522.900 618.600 523.650 ;
        RECT 616.950 520.800 619.050 522.900 ;
        RECT 620.100 518.700 621.000 524.100 ;
        RECT 621.900 522.300 624.000 523.200 ;
        RECT 629.700 522.300 630.600 531.300 ;
        RECT 631.950 527.100 634.050 529.200 ;
        RECT 632.400 526.350 633.600 527.100 ;
        RECT 631.800 523.950 633.900 526.050 ;
        RECT 621.900 521.100 630.600 522.300 ;
        RECT 619.800 516.600 621.900 518.700 ;
        RECT 623.100 518.100 625.200 520.200 ;
        RECT 627.000 519.300 629.100 521.100 ;
        RECT 623.400 516.000 624.600 517.800 ;
        RECT 610.800 511.950 612.900 514.050 ;
        RECT 613.950 511.950 616.050 514.050 ;
        RECT 622.950 511.950 625.050 516.000 ;
        RECT 604.950 496.950 607.050 499.050 ;
        RECT 607.950 496.950 610.050 499.050 ;
        RECT 602.400 494.400 609.450 495.450 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 596.100 487.950 598.200 490.050 ;
        RECT 602.100 487.950 604.200 490.050 ;
        RECT 585.600 474.600 587.700 476.700 ;
        RECT 588.600 474.600 591.600 476.700 ;
        RECT 602.400 485.400 603.600 487.650 ;
        RECT 602.400 466.050 603.450 485.400 ;
        RECT 604.950 469.950 607.050 472.050 ;
        RECT 601.950 463.950 604.050 466.050 ;
        RECT 601.950 457.950 604.050 460.050 ;
        RECT 580.950 451.950 583.050 454.050 ;
        RECT 581.400 444.900 582.450 451.950 ;
        RECT 589.950 449.100 592.050 451.200 ;
        RECT 590.400 448.350 591.600 449.100 ;
        RECT 598.950 448.950 601.050 451.050 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 587.400 444.900 588.600 445.650 ;
        RECT 593.400 444.900 594.600 445.650 ;
        RECT 599.400 444.900 600.450 448.950 ;
        RECT 580.950 442.800 583.050 444.900 ;
        RECT 586.950 442.800 589.050 444.900 ;
        RECT 592.950 442.800 595.050 444.900 ;
        RECT 598.950 442.800 601.050 444.900 ;
        RECT 586.950 439.650 589.050 441.750 ;
        RECT 577.950 427.950 580.050 430.050 ;
        RECT 571.950 421.950 574.050 424.050 ;
        RECT 583.950 418.950 586.050 421.050 ;
        RECT 574.950 416.100 577.050 418.200 ;
        RECT 575.400 415.350 576.600 416.100 ;
        RECT 574.950 412.950 577.050 415.050 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 571.950 409.950 574.050 412.050 ;
        RECT 578.400 411.000 579.600 412.650 ;
        RECT 568.950 406.950 571.050 409.050 ;
        RECT 565.950 400.950 568.050 403.050 ;
        RECT 572.400 394.050 573.450 409.950 ;
        RECT 577.950 406.950 580.050 411.000 ;
        RECT 571.950 393.450 574.050 394.050 ;
        RECT 569.400 392.400 574.050 393.450 ;
        RECT 556.950 388.950 559.050 391.050 ;
        RECT 547.950 385.950 550.050 388.050 ;
        RECT 565.950 385.950 568.050 388.050 ;
        RECT 547.950 372.000 550.050 376.050 ;
        RECT 557.400 372.450 558.600 372.600 ;
        RECT 548.400 370.350 549.600 372.000 ;
        RECT 557.400 371.400 561.450 372.450 ;
        RECT 557.400 370.350 558.600 371.400 ;
        RECT 548.100 367.950 550.200 370.050 ;
        RECT 551.400 367.950 553.500 370.050 ;
        RECT 556.800 367.950 558.900 370.050 ;
        RECT 551.400 365.400 552.600 367.650 ;
        RECT 551.400 361.050 552.450 365.400 ;
        RECT 550.950 358.950 553.050 361.050 ;
        RECT 544.950 346.950 547.050 349.050 ;
        RECT 560.400 346.050 561.450 371.400 ;
        RECT 562.950 370.950 565.050 373.050 ;
        RECT 563.400 361.050 564.450 370.950 ;
        RECT 562.950 358.950 565.050 361.050 ;
        RECT 566.400 355.050 567.450 385.950 ;
        RECT 569.400 366.900 570.450 392.400 ;
        RECT 571.950 391.950 574.050 392.400 ;
        RECT 573.000 390.450 577.050 391.050 ;
        RECT 572.400 390.000 577.050 390.450 ;
        RECT 571.950 388.950 577.050 390.000 ;
        RECT 571.950 385.950 574.050 388.950 ;
        RECT 584.400 388.050 585.450 418.950 ;
        RECT 587.400 418.050 588.450 439.650 ;
        RECT 602.400 430.050 603.450 457.950 ;
        RECT 589.950 427.950 592.050 430.050 ;
        RECT 601.950 427.950 604.050 430.050 ;
        RECT 586.950 415.950 589.050 418.050 ;
        RECT 587.400 400.050 588.450 415.950 ;
        RECT 586.950 397.950 589.050 400.050 ;
        RECT 583.950 385.950 586.050 388.050 ;
        RECT 574.950 382.950 577.050 385.050 ;
        RECT 575.400 376.050 576.450 382.950 ;
        RECT 586.950 376.950 589.050 379.050 ;
        RECT 574.950 372.000 577.050 376.050 ;
        RECT 575.400 370.350 576.600 372.000 ;
        RECT 580.950 371.100 583.050 373.200 ;
        RECT 581.400 370.350 582.600 371.100 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 568.950 364.800 571.050 366.900 ;
        RECT 578.400 365.400 579.600 367.650 ;
        RECT 574.950 361.950 577.050 364.050 ;
        RECT 565.950 352.950 568.050 355.050 ;
        RECT 562.950 346.950 565.050 349.050 ;
        RECT 553.950 343.950 556.050 346.050 ;
        RECT 559.950 343.950 562.050 346.050 ;
        RECT 526.950 340.950 529.050 343.050 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 487.950 334.950 490.050 337.050 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 475.950 331.800 478.050 333.900 ;
        RECT 488.400 332.400 489.600 334.650 ;
        RECT 494.400 333.900 495.600 334.650 ;
        RECT 506.400 333.900 507.450 337.950 ;
        RECT 515.400 337.350 516.600 339.000 ;
        RECT 521.400 337.350 522.600 339.600 ;
        RECT 538.950 339.000 541.050 343.050 ;
        RECT 539.400 337.350 540.600 339.000 ;
        RECT 511.950 334.950 514.050 337.050 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 493.950 333.450 496.050 333.900 ;
        RECT 493.950 332.400 498.450 333.450 ;
        RECT 488.400 328.050 489.450 332.400 ;
        RECT 493.950 331.800 496.050 332.400 ;
        RECT 487.950 325.950 490.050 328.050 ;
        RECT 472.950 313.950 475.050 316.050 ;
        RECT 464.400 306.300 467.400 308.400 ;
        RECT 468.300 306.300 470.400 308.400 ;
        RECT 487.200 306.300 489.300 308.400 ;
        RECT 451.950 296.100 454.050 298.200 ;
        RECT 460.950 296.100 463.050 298.200 ;
        RECT 452.400 295.350 453.600 296.100 ;
        RECT 443.400 292.350 444.600 294.600 ;
        RECT 451.800 292.950 453.900 295.050 ;
        RECT 457.800 292.950 459.900 295.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 440.400 288.000 441.600 289.650 ;
        RECT 427.950 283.950 430.050 286.050 ;
        RECT 439.950 283.950 442.050 288.000 ;
        RECT 446.400 287.400 447.600 289.650 ;
        RECT 446.400 283.050 447.450 287.400 ;
        RECT 445.950 280.950 448.050 283.050 ;
        RECT 421.950 274.950 424.050 277.050 ;
        RECT 409.950 265.950 412.050 268.050 ;
        RECT 413.700 267.300 415.800 269.400 ;
        RECT 394.950 257.100 397.050 259.200 ;
        RECT 400.950 257.100 403.050 259.200 ;
        RECT 403.950 258.000 406.050 262.050 ;
        RECT 409.950 259.950 412.050 262.050 ;
        RECT 395.400 256.350 396.600 257.100 ;
        RECT 395.100 253.950 397.200 256.050 ;
        RECT 401.400 244.050 402.450 257.100 ;
        RECT 404.400 256.350 405.600 258.000 ;
        RECT 404.100 253.950 406.200 256.050 ;
        RECT 410.400 253.050 411.450 259.950 ;
        RECT 409.950 250.950 412.050 253.050 ;
        RECT 414.300 249.600 415.800 267.300 ;
        RECT 413.700 247.500 415.800 249.600 ;
        RECT 400.950 241.950 403.050 244.050 ;
        RECT 414.300 242.700 415.800 247.500 ;
        RECT 413.700 240.600 415.800 242.700 ;
        RECT 416.700 267.300 418.800 269.400 ;
        RECT 419.700 267.300 421.800 269.400 ;
        RECT 422.700 267.300 424.800 269.400 ;
        RECT 416.700 245.700 417.900 267.300 ;
        RECT 419.700 249.600 421.200 267.300 ;
        RECT 422.700 255.000 423.900 267.300 ;
        RECT 428.100 266.400 430.200 268.500 ;
        RECT 436.200 267.300 438.300 269.400 ;
        RECT 439.200 267.300 441.300 269.400 ;
        RECT 442.200 267.300 444.300 269.400 ;
        RECT 424.800 260.400 426.900 262.500 ;
        RECT 428.700 255.900 429.600 266.400 ;
        RECT 431.100 259.950 433.200 262.050 ;
        RECT 422.100 252.900 424.200 255.000 ;
        RECT 427.500 253.800 429.600 255.900 ;
        RECT 419.100 247.500 421.200 249.600 ;
        RECT 416.700 240.600 418.800 245.700 ;
        RECT 419.700 242.700 421.200 247.500 ;
        RECT 422.700 245.700 423.900 252.900 ;
        RECT 428.700 247.200 429.600 253.800 ;
        RECT 422.100 243.600 424.200 245.700 ;
        RECT 427.500 245.100 429.600 247.200 ;
        RECT 431.400 257.400 432.600 259.650 ;
        RECT 419.700 240.600 421.800 242.700 ;
        RECT 431.400 238.050 432.450 257.400 ;
        RECT 437.100 245.700 438.300 267.300 ;
        RECT 436.200 243.600 438.300 245.700 ;
        RECT 439.500 250.800 440.700 267.300 ;
        RECT 442.500 263.700 443.700 267.300 ;
        RECT 442.500 261.600 444.600 263.700 ;
        RECT 439.500 248.700 441.600 250.800 ;
        RECT 439.500 242.700 440.700 248.700 ;
        RECT 443.100 242.700 444.600 261.600 ;
        RECT 461.400 259.050 462.450 296.100 ;
        RECT 464.400 287.400 465.900 306.300 ;
        RECT 468.300 300.300 469.500 306.300 ;
        RECT 467.400 298.200 469.500 300.300 ;
        RECT 464.400 285.300 466.500 287.400 ;
        RECT 465.300 281.700 466.500 285.300 ;
        RECT 468.300 281.700 469.500 298.200 ;
        RECT 470.700 303.300 472.800 305.400 ;
        RECT 470.700 281.700 471.900 303.300 ;
        RECT 479.400 301.800 481.500 303.900 ;
        RECT 484.800 303.300 486.900 305.400 ;
        RECT 479.400 295.200 480.300 301.800 ;
        RECT 485.100 296.100 486.300 303.300 ;
        RECT 487.800 301.500 489.300 306.300 ;
        RECT 490.200 303.300 492.300 308.400 ;
        RECT 487.800 299.400 489.900 301.500 ;
        RECT 479.400 293.100 481.500 295.200 ;
        RECT 484.800 294.000 486.900 296.100 ;
        RECT 475.950 290.100 478.050 292.200 ;
        RECT 476.400 289.350 477.600 290.100 ;
        RECT 475.800 286.950 477.900 289.050 ;
        RECT 479.400 282.600 480.300 293.100 ;
        RECT 482.100 286.500 484.200 288.600 ;
        RECT 464.700 279.600 466.800 281.700 ;
        RECT 467.700 279.600 469.800 281.700 ;
        RECT 470.700 279.600 472.800 281.700 ;
        RECT 478.800 280.500 480.900 282.600 ;
        RECT 485.100 281.700 486.300 294.000 ;
        RECT 487.800 281.700 489.300 299.400 ;
        RECT 491.100 281.700 492.300 303.300 ;
        RECT 484.200 279.600 486.300 281.700 ;
        RECT 487.200 279.600 489.300 281.700 ;
        RECT 490.200 279.600 492.300 281.700 ;
        RECT 493.200 306.300 495.300 308.400 ;
        RECT 493.200 301.500 494.700 306.300 ;
        RECT 493.200 299.400 495.300 301.500 ;
        RECT 493.200 281.700 494.700 299.400 ;
        RECT 493.200 279.600 495.300 281.700 ;
        RECT 497.400 274.050 498.450 332.400 ;
        RECT 505.950 331.800 508.050 333.900 ;
        RECT 512.400 332.400 513.600 334.650 ;
        RECT 518.400 333.900 519.600 334.650 ;
        RECT 512.400 328.050 513.450 332.400 ;
        RECT 517.950 331.800 520.050 333.900 ;
        RECT 542.400 332.400 543.600 334.650 ;
        RECT 542.400 328.050 543.450 332.400 ;
        RECT 554.400 331.050 555.450 343.950 ;
        RECT 563.400 339.600 564.450 346.950 ;
        RECT 563.400 337.350 564.600 339.600 ;
        RECT 568.950 338.100 571.050 340.200 ;
        RECT 569.400 337.350 570.600 338.100 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 560.400 332.400 561.600 334.650 ;
        RECT 566.400 333.000 567.600 334.650 ;
        RECT 553.950 328.950 556.050 331.050 ;
        RECT 511.950 325.950 514.050 328.050 ;
        RECT 541.950 325.950 544.050 328.050 ;
        RECT 560.400 319.050 561.450 332.400 ;
        RECT 565.950 328.950 568.050 333.000 ;
        RECT 559.950 316.950 562.050 319.050 ;
        RECT 514.950 313.950 517.050 316.050 ;
        RECT 505.950 307.950 508.050 310.050 ;
        RECT 502.800 292.950 504.900 295.050 ;
        RECT 503.400 290.400 504.600 292.650 ;
        RECT 503.400 277.050 504.450 290.400 ;
        RECT 506.400 283.050 507.450 307.950 ;
        RECT 511.800 292.950 513.900 295.050 ;
        RECT 512.400 291.450 513.600 292.650 ;
        RECT 509.400 290.400 513.600 291.450 ;
        RECT 505.950 280.950 508.050 283.050 ;
        RECT 509.400 279.450 510.450 290.400 ;
        RECT 515.400 286.050 516.450 313.950 ;
        RECT 533.400 306.300 536.400 308.400 ;
        RECT 537.300 306.300 539.400 308.400 ;
        RECT 556.200 306.300 558.300 308.400 ;
        RECT 520.950 296.100 523.050 298.200 ;
        RECT 521.400 295.350 522.600 296.100 ;
        RECT 520.800 292.950 522.900 295.050 ;
        RECT 526.800 292.950 528.900 295.050 ;
        RECT 517.950 290.100 520.050 292.200 ;
        RECT 514.950 283.950 517.050 286.050 ;
        RECT 518.400 283.050 519.450 290.100 ;
        RECT 533.400 287.400 534.900 306.300 ;
        RECT 537.300 300.300 538.500 306.300 ;
        RECT 536.400 298.200 538.500 300.300 ;
        RECT 533.400 285.300 535.500 287.400 ;
        RECT 517.950 280.950 520.050 283.050 ;
        RECT 534.300 281.700 535.500 285.300 ;
        RECT 537.300 281.700 538.500 298.200 ;
        RECT 539.700 303.300 541.800 305.400 ;
        RECT 539.700 281.700 540.900 303.300 ;
        RECT 548.400 301.800 550.500 303.900 ;
        RECT 553.800 303.300 555.900 305.400 ;
        RECT 544.950 298.950 547.050 301.050 ;
        RECT 545.400 291.600 546.450 298.950 ;
        RECT 548.400 295.200 549.300 301.800 ;
        RECT 554.100 296.100 555.300 303.300 ;
        RECT 556.800 301.500 558.300 306.300 ;
        RECT 559.200 303.300 561.300 308.400 ;
        RECT 556.800 299.400 558.900 301.500 ;
        RECT 548.400 293.100 550.500 295.200 ;
        RECT 553.800 294.000 555.900 296.100 ;
        RECT 545.400 289.350 546.600 291.600 ;
        RECT 544.800 286.950 546.900 289.050 ;
        RECT 548.400 282.600 549.300 293.100 ;
        RECT 551.100 286.500 553.200 288.600 ;
        RECT 517.950 279.450 520.050 279.900 ;
        RECT 533.700 279.600 535.800 281.700 ;
        RECT 536.700 279.600 538.800 281.700 ;
        RECT 539.700 279.600 541.800 281.700 ;
        RECT 547.800 280.500 549.900 282.600 ;
        RECT 554.100 281.700 555.300 294.000 ;
        RECT 556.800 281.700 558.300 299.400 ;
        RECT 560.100 281.700 561.300 303.300 ;
        RECT 553.200 279.600 555.300 281.700 ;
        RECT 556.200 279.600 558.300 281.700 ;
        RECT 559.200 279.600 561.300 281.700 ;
        RECT 562.200 306.300 564.300 308.400 ;
        RECT 562.200 301.500 563.700 306.300 ;
        RECT 562.200 299.400 564.300 301.500 ;
        RECT 562.200 281.700 563.700 299.400 ;
        RECT 565.950 295.950 568.050 298.050 ;
        RECT 562.200 279.600 564.300 281.700 ;
        RECT 566.400 280.050 567.450 295.950 ;
        RECT 571.800 292.950 573.900 295.050 ;
        RECT 572.400 290.400 573.600 292.650 ;
        RECT 568.950 283.950 571.050 286.050 ;
        RECT 509.400 278.400 520.050 279.450 ;
        RECT 517.950 277.800 520.050 278.400 ;
        RECT 565.950 277.950 568.050 280.050 ;
        RECT 502.950 274.950 505.050 277.050 ;
        RECT 514.950 274.950 517.050 277.050 ;
        RECT 496.950 271.950 499.050 274.050 ;
        RECT 508.950 271.950 511.050 274.050 ;
        RECT 476.700 267.300 478.800 269.400 ;
        RECT 479.700 267.300 481.800 269.400 ;
        RECT 482.700 267.300 484.800 269.400 ;
        RECT 477.300 263.700 478.500 267.300 ;
        RECT 476.400 261.600 478.500 263.700 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 449.100 253.950 451.200 256.050 ;
        RECT 455.100 253.950 457.200 256.050 ;
        RECT 463.800 253.950 465.900 256.050 ;
        RECT 469.800 253.950 471.900 256.050 ;
        RECT 455.400 252.900 456.600 253.650 ;
        RECT 464.400 252.900 465.600 253.650 ;
        RECT 454.950 250.800 457.050 252.900 ;
        RECT 463.950 250.800 466.050 252.900 ;
        RECT 438.600 240.600 440.700 242.700 ;
        RECT 441.600 240.600 444.600 242.700 ;
        RECT 476.400 242.700 477.900 261.600 ;
        RECT 480.300 250.800 481.500 267.300 ;
        RECT 479.400 248.700 481.500 250.800 ;
        RECT 480.300 242.700 481.500 248.700 ;
        RECT 482.700 245.700 483.900 267.300 ;
        RECT 490.800 266.400 492.900 268.500 ;
        RECT 496.200 267.300 498.300 269.400 ;
        RECT 499.200 267.300 501.300 269.400 ;
        RECT 502.200 267.300 504.300 269.400 ;
        RECT 487.800 259.950 489.900 262.050 ;
        RECT 488.400 258.900 489.600 259.650 ;
        RECT 487.950 256.800 490.050 258.900 ;
        RECT 491.400 255.900 492.300 266.400 ;
        RECT 494.100 260.400 496.200 262.500 ;
        RECT 491.400 253.800 493.500 255.900 ;
        RECT 497.100 255.000 498.300 267.300 ;
        RECT 487.950 250.800 490.050 252.900 ;
        RECT 482.700 243.600 484.800 245.700 ;
        RECT 476.400 240.600 479.400 242.700 ;
        RECT 480.300 240.600 482.400 242.700 ;
        RECT 484.950 238.950 487.050 241.050 ;
        RECT 430.950 235.950 433.050 238.050 ;
        RECT 439.950 235.950 442.050 238.050 ;
        RECT 395.700 228.300 397.800 230.400 ;
        RECT 396.300 223.500 397.800 228.300 ;
        RECT 395.700 221.400 397.800 223.500 ;
        RECT 396.300 203.700 397.800 221.400 ;
        RECT 395.700 201.600 397.800 203.700 ;
        RECT 398.700 225.300 400.800 230.400 ;
        RECT 401.700 228.300 403.800 230.400 ;
        RECT 412.950 229.950 415.050 232.050 ;
        RECT 398.700 203.700 399.900 225.300 ;
        RECT 401.700 223.500 403.200 228.300 ;
        RECT 404.100 225.300 406.200 227.400 ;
        RECT 401.100 221.400 403.200 223.500 ;
        RECT 401.700 203.700 403.200 221.400 ;
        RECT 404.700 218.100 405.900 225.300 ;
        RECT 409.500 223.800 411.600 225.900 ;
        RECT 404.100 216.000 406.200 218.100 ;
        RECT 410.700 217.200 411.600 223.800 ;
        RECT 404.700 203.700 405.900 216.000 ;
        RECT 409.500 215.100 411.600 217.200 ;
        RECT 406.800 208.500 408.900 210.600 ;
        RECT 410.700 204.600 411.600 215.100 ;
        RECT 413.400 213.600 414.450 229.950 ;
        RECT 420.600 228.300 422.700 230.400 ;
        RECT 423.600 228.300 426.600 230.400 ;
        RECT 418.200 225.300 420.300 227.400 ;
        RECT 413.400 211.350 414.600 213.600 ;
        RECT 413.100 208.950 415.200 211.050 ;
        RECT 398.700 201.600 400.800 203.700 ;
        RECT 401.700 201.600 403.800 203.700 ;
        RECT 404.700 201.600 406.800 203.700 ;
        RECT 410.100 202.500 412.200 204.600 ;
        RECT 419.100 203.700 420.300 225.300 ;
        RECT 421.500 222.300 422.700 228.300 ;
        RECT 421.500 220.200 423.600 222.300 ;
        RECT 421.500 203.700 422.700 220.200 ;
        RECT 425.100 209.400 426.600 228.300 ;
        RECT 440.400 223.050 441.450 235.950 ;
        RECT 445.950 229.800 448.050 231.900 ;
        RECT 460.950 229.950 463.050 232.050 ;
        RECT 478.950 229.950 481.050 232.050 ;
        RECT 439.950 220.950 442.050 223.050 ;
        RECT 427.950 218.100 430.050 220.200 ;
        RECT 436.950 218.100 439.050 220.200 ;
        RECT 424.500 207.300 426.600 209.400 ;
        RECT 424.500 203.700 425.700 207.300 ;
        RECT 418.200 201.600 420.300 203.700 ;
        RECT 421.200 201.600 423.300 203.700 ;
        RECT 424.200 201.600 426.300 203.700 ;
        RECT 428.400 199.050 429.450 218.100 ;
        RECT 437.400 217.350 438.600 218.100 ;
        RECT 431.100 214.950 433.200 217.050 ;
        RECT 437.100 214.950 439.200 217.050 ;
        RECT 446.400 211.050 447.450 229.800 ;
        RECT 461.400 216.600 462.450 229.950 ;
        RECT 472.950 220.950 475.050 223.050 ;
        RECT 461.400 214.350 462.600 216.600 ;
        RECT 466.950 215.100 469.050 217.200 ;
        RECT 467.400 214.350 468.600 215.100 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 445.950 208.950 448.050 211.050 ;
        RECT 458.400 209.400 459.600 211.650 ;
        RECT 464.400 210.900 465.600 211.650 ;
        RECT 473.400 211.050 474.450 220.950 ;
        RECT 479.400 220.050 480.450 229.950 ;
        RECT 485.400 223.050 486.450 238.950 ;
        RECT 488.400 229.050 489.450 250.800 ;
        RECT 491.400 247.200 492.300 253.800 ;
        RECT 496.800 252.900 498.900 255.000 ;
        RECT 491.400 245.100 493.500 247.200 ;
        RECT 497.100 245.700 498.300 252.900 ;
        RECT 499.800 249.600 501.300 267.300 ;
        RECT 499.800 247.500 501.900 249.600 ;
        RECT 496.800 243.600 498.900 245.700 ;
        RECT 499.800 242.700 501.300 247.500 ;
        RECT 503.100 245.700 504.300 267.300 ;
        RECT 499.200 240.600 501.300 242.700 ;
        RECT 502.200 240.600 504.300 245.700 ;
        RECT 505.200 267.300 507.300 269.400 ;
        RECT 505.200 249.600 506.700 267.300 ;
        RECT 505.200 247.500 507.300 249.600 ;
        RECT 505.200 242.700 506.700 247.500 ;
        RECT 505.200 240.600 507.300 242.700 ;
        RECT 487.950 226.950 490.050 229.050 ;
        RECT 484.950 220.950 487.050 223.050 ;
        RECT 505.950 220.950 508.050 223.050 ;
        RECT 478.950 217.950 481.050 220.050 ;
        RECT 475.950 215.100 478.050 217.200 ;
        RECT 487.950 216.000 490.050 220.050 ;
        RECT 430.950 202.950 433.050 205.050 ;
        RECT 394.950 196.950 397.050 199.050 ;
        RECT 427.950 196.950 430.050 199.050 ;
        RECT 389.400 182.400 393.450 183.450 ;
        RECT 395.400 183.600 396.450 196.950 ;
        RECT 385.950 169.950 388.050 172.050 ;
        RECT 379.950 166.950 382.050 169.050 ;
        RECT 367.950 163.950 370.050 166.050 ;
        RECT 376.950 163.950 379.050 166.050 ;
        RECT 349.950 151.950 352.050 154.050 ;
        RECT 361.950 151.950 364.050 154.050 ;
        RECT 332.400 130.050 333.450 131.400 ;
        RECT 337.950 130.800 340.050 132.900 ;
        RECT 346.950 130.950 349.050 133.050 ;
        RECT 331.950 127.950 334.050 130.050 ;
        RECT 325.950 121.950 328.050 124.050 ;
        RECT 332.400 118.050 333.450 127.950 ;
        RECT 350.400 127.050 351.450 151.950 ;
        RECT 362.400 138.600 363.450 151.950 ;
        RECT 367.950 142.950 370.050 145.050 ;
        RECT 362.400 136.350 363.600 138.600 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 359.400 131.400 360.600 133.650 ;
        RECT 359.400 127.050 360.450 131.400 ;
        RECT 349.950 124.950 352.050 127.050 ;
        RECT 358.950 124.950 361.050 127.050 ;
        RECT 292.950 115.950 295.050 118.050 ;
        RECT 298.950 115.950 301.050 118.050 ;
        RECT 310.950 115.950 313.050 118.050 ;
        RECT 319.950 115.950 322.050 118.050 ;
        RECT 331.950 115.950 334.050 118.050 ;
        RECT 293.400 105.600 294.450 115.950 ;
        RECT 298.950 106.950 301.050 109.050 ;
        RECT 304.950 106.950 307.050 109.050 ;
        RECT 293.400 103.350 294.600 105.600 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 299.400 102.600 300.450 106.950 ;
        RECT 259.950 94.950 262.050 97.050 ;
        RECT 268.950 94.950 271.050 99.000 ;
        RECT 277.950 97.800 280.050 99.900 ;
        RECT 283.950 97.950 286.050 100.050 ;
        RECT 290.400 99.900 291.600 100.650 ;
        RECT 299.400 100.350 300.600 102.600 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 299.100 97.950 301.200 100.050 ;
        RECT 256.950 64.950 259.050 67.050 ;
        RECT 239.400 58.350 240.600 59.100 ;
        RECT 250.950 58.950 253.050 61.050 ;
        RECT 260.400 60.600 261.450 94.950 ;
        RECT 305.400 82.050 306.450 106.950 ;
        RECT 308.400 102.450 309.600 102.600 ;
        RECT 311.400 102.450 312.450 115.950 ;
        RECT 317.700 111.300 319.800 113.400 ;
        RECT 308.400 101.400 312.450 102.450 ;
        RECT 308.400 100.350 309.600 101.400 ;
        RECT 308.100 97.950 310.200 100.050 ;
        RECT 313.950 97.950 316.050 100.050 ;
        RECT 304.950 79.950 307.050 82.050 ;
        RECT 274.950 73.950 277.050 76.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 226.800 52.800 228.900 54.900 ;
        RECT 229.950 52.950 232.050 55.050 ;
        RECT 236.400 54.900 237.600 55.650 ;
        RECT 251.400 54.900 252.450 58.950 ;
        RECT 260.400 58.350 261.600 60.600 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 235.950 52.800 238.050 54.900 ;
        RECT 250.950 52.800 253.050 54.900 ;
        RECT 257.400 53.400 258.600 55.650 ;
        RECT 263.400 54.900 264.600 55.650 ;
        RECT 275.400 54.900 276.450 73.950 ;
        RECT 304.800 64.950 306.900 67.050 ;
        RECT 283.950 59.100 286.050 61.200 ;
        RECT 289.950 60.000 292.050 64.050 ;
        RECT 284.400 58.350 285.600 59.100 ;
        RECT 290.400 58.350 291.600 60.000 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 281.400 54.900 282.600 55.650 ;
        RECT 257.400 49.050 258.450 53.400 ;
        RECT 262.950 52.800 265.050 54.900 ;
        RECT 274.950 52.800 277.050 54.900 ;
        RECT 280.950 52.800 283.050 54.900 ;
        RECT 287.400 53.400 288.600 55.650 ;
        RECT 293.400 53.400 294.600 55.650 ;
        RECT 305.400 54.900 306.450 64.950 ;
        RECT 307.950 61.950 310.050 67.050 ;
        RECT 314.400 61.200 315.450 97.950 ;
        RECT 318.300 93.600 319.800 111.300 ;
        RECT 317.700 91.500 319.800 93.600 ;
        RECT 318.300 86.700 319.800 91.500 ;
        RECT 317.700 84.600 319.800 86.700 ;
        RECT 320.700 111.300 322.800 113.400 ;
        RECT 323.700 111.300 325.800 113.400 ;
        RECT 326.700 111.300 328.800 113.400 ;
        RECT 320.700 89.700 321.900 111.300 ;
        RECT 323.700 93.600 325.200 111.300 ;
        RECT 326.700 99.000 327.900 111.300 ;
        RECT 332.100 110.400 334.200 112.500 ;
        RECT 340.200 111.300 342.300 113.400 ;
        RECT 343.200 111.300 345.300 113.400 ;
        RECT 346.200 111.300 348.300 113.400 ;
        RECT 328.800 104.400 330.900 106.500 ;
        RECT 332.700 99.900 333.600 110.400 ;
        RECT 335.100 103.950 337.200 106.050 ;
        RECT 335.400 102.900 336.600 103.650 ;
        RECT 334.950 100.800 337.050 102.900 ;
        RECT 326.100 96.900 328.200 99.000 ;
        RECT 331.500 97.800 333.600 99.900 ;
        RECT 323.100 91.500 325.200 93.600 ;
        RECT 320.700 84.600 322.800 89.700 ;
        RECT 323.700 86.700 325.200 91.500 ;
        RECT 326.700 89.700 327.900 96.900 ;
        RECT 332.700 91.200 333.600 97.800 ;
        RECT 326.100 87.600 328.200 89.700 ;
        RECT 331.500 89.100 333.600 91.200 ;
        RECT 341.100 89.700 342.300 111.300 ;
        RECT 340.200 87.600 342.300 89.700 ;
        RECT 343.500 94.800 344.700 111.300 ;
        RECT 346.500 107.700 347.700 111.300 ;
        RECT 349.950 109.950 352.050 112.050 ;
        RECT 346.500 105.600 348.600 107.700 ;
        RECT 343.500 92.700 345.600 94.800 ;
        RECT 343.500 86.700 344.700 92.700 ;
        RECT 347.100 86.700 348.600 105.600 ;
        RECT 350.400 102.900 351.450 109.950 ;
        RECT 349.950 100.800 352.050 102.900 ;
        RECT 353.100 97.950 355.200 100.050 ;
        RECT 359.100 97.950 361.200 100.050 ;
        RECT 359.400 96.900 360.600 97.650 ;
        RECT 358.950 94.800 361.050 96.900 ;
        RECT 323.700 84.600 325.800 86.700 ;
        RECT 342.600 84.600 344.700 86.700 ;
        RECT 345.600 84.600 348.600 86.700 ;
        RECT 340.950 79.950 343.050 82.050 ;
        RECT 355.950 79.950 358.050 82.050 ;
        RECT 319.950 64.950 322.050 67.050 ;
        RECT 313.950 59.100 316.050 61.200 ;
        RECT 320.400 60.600 321.450 64.950 ;
        RECT 341.400 60.600 342.450 79.950 ;
        RECT 314.400 58.350 315.600 59.100 ;
        RECT 320.400 58.350 321.600 60.600 ;
        RECT 341.400 58.350 342.600 60.600 ;
        RECT 346.950 59.100 349.050 61.200 ;
        RECT 347.400 58.350 348.600 59.100 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 311.400 54.900 312.600 55.650 ;
        RECT 247.950 46.950 250.050 49.050 ;
        RECT 256.950 46.950 259.050 49.050 ;
        RECT 223.950 43.950 226.050 46.050 ;
        RECT 218.400 25.350 219.600 27.600 ;
        RECT 232.950 27.450 235.050 28.200 ;
        RECT 236.400 27.450 237.600 27.600 ;
        RECT 232.950 26.400 237.600 27.450 ;
        RECT 232.950 26.100 235.050 26.400 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 215.400 21.900 216.600 22.650 ;
        RECT 233.400 22.050 234.450 26.100 ;
        RECT 236.400 25.350 237.600 26.400 ;
        RECT 236.400 22.950 238.500 25.050 ;
        RECT 241.800 22.950 243.900 25.050 ;
        RECT 248.400 24.600 249.450 46.950 ;
        RECT 287.400 40.050 288.450 53.400 ;
        RECT 293.400 46.050 294.450 53.400 ;
        RECT 304.950 52.800 307.050 54.900 ;
        RECT 310.950 52.800 313.050 54.900 ;
        RECT 317.400 53.400 318.600 55.650 ;
        RECT 323.400 54.900 324.600 55.650 ;
        RECT 292.950 43.950 295.050 46.050 ;
        RECT 286.950 37.950 289.050 40.050 ;
        RECT 298.950 37.950 301.050 40.050 ;
        RECT 266.700 33.300 268.800 35.400 ;
        RECT 248.400 22.350 249.600 24.600 ;
        RECT 256.950 24.000 259.050 28.050 ;
        RECT 257.400 22.350 258.600 24.000 ;
        RECT 214.950 19.800 217.050 21.900 ;
        RECT 232.950 19.950 235.050 22.050 ;
        RECT 248.100 19.950 250.200 22.050 ;
        RECT 257.100 19.950 259.200 22.050 ;
        RECT 267.300 15.600 268.800 33.300 ;
        RECT 266.700 13.500 268.800 15.600 ;
        RECT 205.950 10.950 208.050 13.050 ;
        RECT 267.300 8.700 268.800 13.500 ;
        RECT 266.700 6.600 268.800 8.700 ;
        RECT 269.700 33.300 271.800 35.400 ;
        RECT 272.700 33.300 274.800 35.400 ;
        RECT 275.700 33.300 277.800 35.400 ;
        RECT 269.700 11.700 270.900 33.300 ;
        RECT 272.700 15.600 274.200 33.300 ;
        RECT 275.700 21.000 276.900 33.300 ;
        RECT 281.100 32.400 283.200 34.500 ;
        RECT 289.200 33.300 291.300 35.400 ;
        RECT 292.200 33.300 294.300 35.400 ;
        RECT 295.200 33.300 297.300 35.400 ;
        RECT 277.800 26.400 279.900 28.500 ;
        RECT 281.700 21.900 282.600 32.400 ;
        RECT 284.100 25.950 286.200 28.050 ;
        RECT 284.400 24.900 285.600 25.650 ;
        RECT 283.950 22.800 286.050 24.900 ;
        RECT 275.100 18.900 277.200 21.000 ;
        RECT 280.500 19.800 282.600 21.900 ;
        RECT 272.100 13.500 274.200 15.600 ;
        RECT 269.700 6.600 271.800 11.700 ;
        RECT 272.700 8.700 274.200 13.500 ;
        RECT 275.700 11.700 276.900 18.900 ;
        RECT 281.700 13.200 282.600 19.800 ;
        RECT 275.100 9.600 277.200 11.700 ;
        RECT 280.500 11.100 282.600 13.200 ;
        RECT 290.100 11.700 291.300 33.300 ;
        RECT 289.200 9.600 291.300 11.700 ;
        RECT 292.500 16.800 293.700 33.300 ;
        RECT 295.500 29.700 296.700 33.300 ;
        RECT 295.500 27.600 297.600 29.700 ;
        RECT 292.500 14.700 294.600 16.800 ;
        RECT 292.500 8.700 293.700 14.700 ;
        RECT 296.100 8.700 297.600 27.600 ;
        RECT 299.400 24.900 300.450 37.950 ;
        RECT 317.400 27.450 318.450 53.400 ;
        RECT 322.950 52.800 325.050 54.900 ;
        RECT 344.400 53.400 345.600 55.650 ;
        RECT 344.400 40.050 345.450 53.400 ;
        RECT 349.950 52.800 352.050 54.900 ;
        RECT 350.400 43.050 351.450 52.800 ;
        RECT 356.400 52.050 357.450 79.950 ;
        RECT 355.950 49.950 358.050 52.050 ;
        RECT 349.950 40.950 352.050 43.050 ;
        RECT 343.950 37.950 346.050 40.050 ;
        RECT 359.400 39.450 360.450 94.800 ;
        RECT 368.400 85.050 369.450 142.950 ;
        RECT 370.950 136.950 373.050 139.050 ;
        RECT 371.400 96.900 372.450 136.950 ;
        RECT 377.400 124.050 378.450 163.950 ;
        RECT 380.400 139.200 381.450 166.950 ;
        RECT 382.950 163.950 385.050 166.050 ;
        RECT 383.400 148.050 384.450 163.950 ;
        RECT 382.950 145.950 385.050 148.050 ;
        RECT 386.400 145.050 387.450 169.950 ;
        RECT 385.950 142.950 388.050 145.050 ;
        RECT 379.950 137.100 382.050 139.200 ;
        RECT 380.400 136.350 381.600 137.100 ;
        RECT 380.100 133.950 382.200 136.050 ;
        RECT 385.500 133.950 387.600 136.050 ;
        RECT 386.400 132.900 387.600 133.650 ;
        RECT 385.950 130.800 388.050 132.900 ;
        RECT 389.400 127.050 390.450 182.400 ;
        RECT 395.400 181.350 396.600 183.600 ;
        RECT 400.950 182.100 403.050 184.200 ;
        RECT 401.400 181.350 402.600 182.100 ;
        RECT 409.950 181.950 412.050 184.050 ;
        RECT 415.950 182.100 418.050 184.200 ;
        RECT 424.950 182.100 427.050 184.200 ;
        RECT 431.400 183.600 432.450 202.950 ;
        RECT 433.950 196.950 436.050 199.050 ;
        RECT 442.950 196.950 445.050 199.050 ;
        RECT 454.950 196.950 457.050 199.050 ;
        RECT 434.400 184.050 435.450 196.950 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 397.950 178.950 400.050 181.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 398.400 177.000 399.600 178.650 ;
        RECT 404.400 177.000 405.600 178.650 ;
        RECT 397.950 172.950 400.050 177.000 ;
        RECT 403.950 172.950 406.050 177.000 ;
        RECT 410.400 175.050 411.450 181.950 ;
        RECT 416.400 175.050 417.450 182.100 ;
        RECT 425.400 181.350 426.600 182.100 ;
        RECT 431.400 181.350 432.600 183.600 ;
        RECT 433.950 181.950 436.050 184.050 ;
        RECT 439.950 182.100 442.050 184.200 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 422.400 177.000 423.600 178.650 ;
        RECT 409.950 172.950 412.050 175.050 ;
        RECT 415.950 172.950 418.050 175.050 ;
        RECT 421.950 172.950 424.050 177.000 ;
        RECT 428.400 176.400 429.600 178.650 ;
        RECT 428.400 166.050 429.450 176.400 ;
        RECT 433.950 169.950 436.050 172.050 ;
        RECT 434.400 166.050 435.450 169.950 ;
        RECT 427.950 163.950 430.050 166.050 ;
        RECT 433.950 163.950 436.050 166.050 ;
        RECT 440.400 157.050 441.450 182.100 ;
        RECT 439.950 154.950 442.050 157.050 ;
        RECT 397.950 142.950 400.050 145.050 ;
        RECT 398.400 132.900 399.450 142.950 ;
        RECT 406.950 137.100 409.050 139.200 ;
        RECT 407.400 136.350 408.600 137.100 ;
        RECT 421.950 136.950 424.050 139.050 ;
        RECT 427.950 137.100 430.050 139.200 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 406.950 133.950 409.050 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 397.950 130.800 400.050 132.900 ;
        RECT 404.400 131.400 405.600 133.650 ;
        RECT 410.400 132.900 411.600 133.650 ;
        RECT 422.400 132.900 423.450 136.950 ;
        RECT 428.400 136.350 429.600 137.100 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 430.950 133.950 433.050 136.050 ;
        RECT 431.400 132.900 432.600 133.650 ;
        RECT 388.950 124.950 391.050 127.050 ;
        RECT 397.950 124.950 400.050 127.050 ;
        RECT 376.950 121.950 379.050 124.050 ;
        RECT 385.950 109.950 388.050 112.050 ;
        RECT 373.950 104.100 376.050 106.200 ;
        RECT 379.950 104.100 382.050 106.200 ;
        RECT 386.400 105.600 387.450 109.950 ;
        RECT 370.950 94.800 373.050 96.900 ;
        RECT 367.950 82.950 370.050 85.050 ;
        RECT 374.400 79.050 375.450 104.100 ;
        RECT 380.400 103.350 381.600 104.100 ;
        RECT 386.400 103.350 387.600 105.600 ;
        RECT 391.950 104.100 394.050 106.200 ;
        RECT 392.400 103.350 393.600 104.100 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 383.400 99.900 384.600 100.650 ;
        RECT 382.950 97.800 385.050 99.900 ;
        RECT 389.400 98.400 390.600 100.650 ;
        RECT 398.400 99.900 399.450 124.950 ;
        RECT 404.400 124.050 405.450 131.400 ;
        RECT 409.950 130.800 412.050 132.900 ;
        RECT 418.800 130.800 420.900 132.900 ;
        RECT 421.950 130.800 424.050 132.900 ;
        RECT 430.950 130.800 433.050 132.900 ;
        RECT 403.950 121.950 406.050 124.050 ;
        RECT 406.950 118.950 409.050 121.050 ;
        RECT 407.400 106.200 408.450 118.950 ;
        RECT 409.950 115.950 412.050 118.050 ;
        RECT 406.950 104.100 409.050 106.200 ;
        RECT 410.400 105.600 411.450 115.950 ;
        RECT 410.400 103.350 411.600 105.600 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 389.400 85.050 390.450 98.400 ;
        RECT 397.950 97.800 400.050 99.900 ;
        RECT 413.400 98.400 414.600 100.650 ;
        RECT 391.950 94.950 394.050 97.050 ;
        RECT 376.950 82.950 379.050 85.050 ;
        RECT 388.950 82.950 391.050 85.050 ;
        RECT 373.950 76.950 376.050 79.050 ;
        RECT 370.950 70.950 373.050 73.050 ;
        RECT 364.950 59.100 367.050 61.200 ;
        RECT 365.400 58.350 366.600 59.100 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 368.400 54.000 369.600 55.650 ;
        RECT 364.950 49.950 367.050 52.050 ;
        RECT 367.950 49.950 370.050 54.000 ;
        RECT 359.400 38.400 363.450 39.450 ;
        RECT 329.700 33.300 331.800 35.400 ;
        RECT 332.700 33.300 334.800 35.400 ;
        RECT 335.700 33.300 337.800 35.400 ;
        RECT 330.300 29.700 331.500 33.300 ;
        RECT 329.400 27.600 331.500 29.700 ;
        RECT 317.400 27.000 321.450 27.450 ;
        RECT 317.400 26.400 322.050 27.000 ;
        RECT 298.950 22.800 301.050 24.900 ;
        RECT 319.950 22.800 322.050 26.400 ;
        RECT 302.100 19.950 304.200 22.050 ;
        RECT 308.100 19.950 310.200 22.050 ;
        RECT 316.800 19.950 318.900 22.050 ;
        RECT 322.800 19.950 324.900 22.050 ;
        RECT 308.400 18.900 309.600 19.650 ;
        RECT 317.400 18.900 318.600 19.650 ;
        RECT 307.950 16.800 310.050 18.900 ;
        RECT 316.950 16.800 319.050 18.900 ;
        RECT 272.700 6.600 274.800 8.700 ;
        RECT 291.600 6.600 293.700 8.700 ;
        RECT 294.600 6.600 297.600 8.700 ;
        RECT 329.400 8.700 330.900 27.600 ;
        RECT 333.300 16.800 334.500 33.300 ;
        RECT 332.400 14.700 334.500 16.800 ;
        RECT 333.300 8.700 334.500 14.700 ;
        RECT 335.700 11.700 336.900 33.300 ;
        RECT 343.800 32.400 345.900 34.500 ;
        RECT 349.200 33.300 351.300 35.400 ;
        RECT 352.200 33.300 354.300 35.400 ;
        RECT 355.200 33.300 357.300 35.400 ;
        RECT 340.800 25.950 342.900 28.050 ;
        RECT 341.400 24.900 342.600 25.650 ;
        RECT 340.950 22.800 343.050 24.900 ;
        RECT 344.400 21.900 345.300 32.400 ;
        RECT 347.100 26.400 349.200 28.500 ;
        RECT 344.400 19.800 346.500 21.900 ;
        RECT 350.100 21.000 351.300 33.300 ;
        RECT 344.400 13.200 345.300 19.800 ;
        RECT 349.800 18.900 351.900 21.000 ;
        RECT 335.700 9.600 337.800 11.700 ;
        RECT 344.400 11.100 346.500 13.200 ;
        RECT 350.100 11.700 351.300 18.900 ;
        RECT 352.800 15.600 354.300 33.300 ;
        RECT 352.800 13.500 354.900 15.600 ;
        RECT 349.800 9.600 351.900 11.700 ;
        RECT 352.800 8.700 354.300 13.500 ;
        RECT 356.100 11.700 357.300 33.300 ;
        RECT 329.400 6.600 332.400 8.700 ;
        RECT 333.300 6.600 335.400 8.700 ;
        RECT 352.200 6.600 354.300 8.700 ;
        RECT 355.200 6.600 357.300 11.700 ;
        RECT 358.200 33.300 360.300 35.400 ;
        RECT 358.200 15.600 359.700 33.300 ;
        RECT 362.400 18.900 363.450 38.400 ;
        RECT 365.400 37.050 366.450 49.950 ;
        RECT 364.950 34.950 367.050 37.050 ;
        RECT 377.400 31.050 378.450 82.950 ;
        RECT 385.950 76.950 388.050 79.050 ;
        RECT 379.950 70.950 382.050 76.050 ;
        RECT 379.950 59.100 382.050 61.200 ;
        RECT 386.400 60.600 387.450 76.950 ;
        RECT 389.400 67.050 390.450 82.950 ;
        RECT 388.950 64.950 391.050 67.050 ;
        RECT 392.400 61.200 393.450 94.950 ;
        RECT 398.400 73.050 399.450 97.800 ;
        RECT 413.400 79.050 414.450 98.400 ;
        RECT 412.950 76.950 415.050 79.050 ;
        RECT 397.950 70.950 400.050 73.050 ;
        RECT 419.400 64.050 420.450 130.800 ;
        RECT 440.400 112.050 441.450 154.950 ;
        RECT 443.400 151.050 444.450 196.950 ;
        RECT 448.950 187.950 451.050 190.050 ;
        RECT 449.400 184.200 450.450 187.950 ;
        RECT 448.950 182.100 451.050 184.200 ;
        RECT 455.400 183.600 456.450 196.950 ;
        RECT 458.400 190.050 459.450 209.400 ;
        RECT 463.950 208.800 466.050 210.900 ;
        RECT 472.950 208.950 475.050 211.050 ;
        RECT 476.400 202.050 477.450 215.100 ;
        RECT 488.400 214.350 489.600 216.000 ;
        RECT 493.950 215.100 496.050 217.200 ;
        RECT 499.950 215.100 502.050 217.200 ;
        RECT 494.400 214.350 495.600 215.100 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 485.400 209.400 486.600 211.650 ;
        RECT 491.400 210.900 492.600 211.650 ;
        RECT 475.950 199.950 478.050 202.050 ;
        RECT 485.400 199.050 486.450 209.400 ;
        RECT 490.950 208.800 493.050 210.900 ;
        RECT 484.950 196.950 487.050 199.050 ;
        RECT 500.400 196.050 501.450 215.100 ;
        RECT 499.950 193.950 502.050 196.050 ;
        RECT 457.950 187.950 460.050 190.050 ;
        RECT 473.700 189.300 475.800 191.400 ;
        RECT 476.700 189.300 478.800 191.400 ;
        RECT 479.700 189.300 481.800 191.400 ;
        RECT 474.300 185.700 475.500 189.300 ;
        RECT 473.400 183.600 475.500 185.700 ;
        RECT 449.400 181.350 450.600 182.100 ;
        RECT 455.400 181.350 456.600 183.600 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 445.950 175.950 448.050 178.050 ;
        RECT 452.400 177.900 453.600 178.650 ;
        RECT 446.400 169.050 447.450 175.950 ;
        RECT 451.950 175.800 454.050 177.900 ;
        RECT 460.800 175.950 462.900 178.050 ;
        RECT 466.800 175.950 468.900 178.050 ;
        RECT 461.400 173.400 462.600 175.650 ;
        RECT 461.400 169.050 462.450 173.400 ;
        RECT 445.950 166.950 448.050 169.050 ;
        RECT 460.950 166.950 463.050 169.050 ;
        RECT 473.400 164.700 474.900 183.600 ;
        RECT 477.300 172.800 478.500 189.300 ;
        RECT 476.400 170.700 478.500 172.800 ;
        RECT 477.300 164.700 478.500 170.700 ;
        RECT 479.700 167.700 480.900 189.300 ;
        RECT 487.800 188.400 489.900 190.500 ;
        RECT 493.200 189.300 495.300 191.400 ;
        RECT 496.200 189.300 498.300 191.400 ;
        RECT 499.200 189.300 501.300 191.400 ;
        RECT 484.800 181.950 486.900 184.050 ;
        RECT 485.400 179.400 486.600 181.650 ;
        RECT 479.700 165.600 481.800 167.700 ;
        RECT 473.400 162.600 476.400 164.700 ;
        RECT 477.300 162.600 479.400 164.700 ;
        RECT 442.950 148.950 445.050 151.050 ;
        RECT 451.950 145.950 454.050 148.050 ;
        RECT 452.400 138.600 453.450 145.950 ;
        RECT 452.400 136.350 453.600 138.600 ;
        RECT 463.950 136.950 466.050 139.050 ;
        RECT 472.950 137.100 475.050 139.200 ;
        RECT 478.950 137.100 481.050 139.200 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 449.400 133.050 450.600 133.650 ;
        RECT 445.950 131.400 450.600 133.050 ;
        RECT 455.400 132.900 456.600 133.650 ;
        RECT 445.950 130.950 450.000 131.400 ;
        RECT 448.950 127.950 451.050 130.050 ;
        RECT 454.950 127.950 457.050 132.900 ;
        RECT 460.950 127.950 463.050 130.050 ;
        RECT 430.950 109.950 433.050 112.050 ;
        RECT 439.950 109.950 442.050 112.050 ;
        RECT 424.950 104.100 427.050 106.200 ;
        RECT 431.400 105.600 432.450 109.950 ;
        RECT 425.400 97.050 426.450 104.100 ;
        RECT 431.400 103.350 432.600 105.600 ;
        RECT 436.950 104.100 439.050 106.200 ;
        RECT 437.400 103.350 438.600 104.100 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 434.400 99.900 435.600 100.650 ;
        RECT 449.400 100.050 450.450 127.950 ;
        RECT 457.950 109.950 460.050 112.050 ;
        RECT 458.400 105.600 459.450 109.950 ;
        RECT 461.400 109.050 462.450 127.950 ;
        RECT 464.400 126.450 465.450 136.950 ;
        RECT 473.400 136.350 474.600 137.100 ;
        RECT 479.400 136.350 480.600 137.100 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 470.400 132.000 471.600 133.650 ;
        RECT 469.950 127.950 472.050 132.000 ;
        RECT 476.400 131.400 477.600 133.650 ;
        RECT 476.400 129.450 477.450 131.400 ;
        RECT 473.400 128.400 477.450 129.450 ;
        RECT 473.400 126.450 474.450 128.400 ;
        RECT 464.400 125.400 474.450 126.450 ;
        RECT 478.950 115.950 481.050 118.050 ;
        RECT 460.950 106.950 463.050 109.050 ;
        RECT 466.950 106.950 469.050 109.050 ;
        RECT 458.400 103.350 459.600 105.600 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 433.950 97.800 436.050 99.900 ;
        RECT 448.950 97.950 451.050 100.050 ;
        RECT 455.400 98.400 456.600 100.650 ;
        RECT 461.400 99.900 462.600 100.650 ;
        RECT 467.400 99.900 468.450 106.950 ;
        RECT 479.400 105.600 480.450 115.950 ;
        RECT 485.400 105.600 486.450 179.400 ;
        RECT 488.400 177.900 489.300 188.400 ;
        RECT 491.100 182.400 493.200 184.500 ;
        RECT 488.400 175.800 490.500 177.900 ;
        RECT 494.100 177.000 495.300 189.300 ;
        RECT 488.400 169.200 489.300 175.800 ;
        RECT 493.800 174.900 495.900 177.000 ;
        RECT 488.400 167.100 490.500 169.200 ;
        RECT 494.100 167.700 495.300 174.900 ;
        RECT 496.800 171.600 498.300 189.300 ;
        RECT 496.800 169.500 498.900 171.600 ;
        RECT 493.800 165.600 495.900 167.700 ;
        RECT 496.800 164.700 498.300 169.500 ;
        RECT 500.100 167.700 501.300 189.300 ;
        RECT 496.200 162.600 498.300 164.700 ;
        RECT 499.200 162.600 501.300 167.700 ;
        RECT 502.200 189.300 504.300 191.400 ;
        RECT 502.200 171.600 503.700 189.300 ;
        RECT 506.400 184.050 507.450 220.950 ;
        RECT 509.400 208.050 510.450 271.950 ;
        RECT 515.400 258.600 516.450 274.950 ;
        RECT 547.950 268.950 550.050 271.050 ;
        RECT 548.400 261.600 549.450 268.950 ;
        RECT 569.400 265.050 570.450 283.950 ;
        RECT 572.400 277.050 573.450 290.400 ;
        RECT 571.950 274.950 574.050 277.050 ;
        RECT 575.400 268.050 576.450 361.950 ;
        RECT 578.400 349.050 579.450 365.400 ;
        RECT 577.950 346.950 580.050 349.050 ;
        RECT 583.950 346.950 586.050 349.050 ;
        RECT 578.400 331.050 579.450 346.950 ;
        RECT 584.400 343.050 585.450 346.950 ;
        RECT 583.950 340.950 586.050 343.050 ;
        RECT 587.400 342.450 588.450 376.950 ;
        RECT 590.400 346.050 591.450 427.950 ;
        RECT 598.950 417.000 601.050 421.050 ;
        RECT 605.400 417.600 606.450 469.950 ;
        RECT 608.400 466.050 609.450 494.400 ;
        RECT 607.950 463.950 610.050 466.050 ;
        RECT 611.400 463.050 612.450 511.950 ;
        RECT 635.400 511.050 636.450 536.400 ;
        RECT 638.400 513.450 639.450 544.950 ;
        RECT 640.950 526.950 643.050 529.050 ;
        RECT 650.400 528.600 651.450 547.950 ;
        RECT 656.400 540.450 657.450 562.800 ;
        RECT 665.400 556.050 666.450 566.400 ;
        RECT 670.950 565.800 673.050 567.900 ;
        RECT 676.950 565.800 679.050 567.900 ;
        RECT 682.950 565.800 685.050 567.900 ;
        RECT 667.950 562.950 670.050 565.050 ;
        RECT 664.950 553.950 667.050 556.050 ;
        RECT 665.400 547.050 666.450 553.950 ;
        RECT 668.400 553.050 669.450 562.950 ;
        RECT 676.950 559.950 679.050 562.050 ;
        RECT 667.950 550.950 670.050 553.050 ;
        RECT 667.950 547.800 670.050 549.900 ;
        RECT 664.950 544.950 667.050 547.050 ;
        RECT 661.950 543.450 664.050 544.050 ;
        RECT 668.400 543.450 669.450 547.800 ;
        RECT 677.400 544.050 678.450 559.950 ;
        RECT 679.950 550.950 682.050 553.050 ;
        RECT 661.950 542.400 669.450 543.450 ;
        RECT 661.950 541.950 664.050 542.400 ;
        RECT 676.950 541.950 679.050 544.050 ;
        RECT 656.400 539.400 660.450 540.450 ;
        RECT 655.950 532.950 658.050 535.050 ;
        RECT 656.400 528.600 657.450 532.950 ;
        RECT 659.400 532.050 660.450 539.400 ;
        RECT 661.950 538.800 664.050 540.900 ;
        RECT 658.950 529.950 661.050 532.050 ;
        RECT 662.400 529.050 663.450 538.800 ;
        RECT 670.950 535.950 673.050 538.050 ;
        RECT 680.400 537.450 681.450 550.950 ;
        RECT 677.400 536.400 681.450 537.450 ;
        RECT 667.950 529.950 670.050 532.050 ;
        RECT 641.400 517.050 642.450 526.950 ;
        RECT 650.400 526.350 651.600 528.600 ;
        RECT 656.400 526.350 657.600 528.600 ;
        RECT 662.400 526.950 667.050 529.050 ;
        RECT 662.400 526.350 663.600 526.950 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 653.400 521.400 654.600 523.650 ;
        RECT 659.400 522.000 660.600 523.650 ;
        RECT 653.400 517.050 654.450 521.400 ;
        RECT 658.950 517.950 661.050 522.000 ;
        RECT 668.400 517.050 669.450 529.950 ;
        RECT 671.400 520.050 672.450 535.950 ;
        RECT 677.400 532.050 678.450 536.400 ;
        RECT 679.950 532.950 682.050 535.050 ;
        RECT 673.950 529.950 676.050 532.050 ;
        RECT 676.950 529.950 679.050 532.050 ;
        RECT 670.950 517.950 673.050 520.050 ;
        RECT 640.950 514.950 643.050 517.050 ;
        RECT 652.950 514.950 655.050 517.050 ;
        RECT 667.950 514.950 670.050 517.050 ;
        RECT 638.400 512.400 642.450 513.450 ;
        RECT 635.400 509.400 640.050 511.050 ;
        RECT 636.000 508.950 640.050 509.400 ;
        RECT 631.950 499.950 634.050 502.050 ;
        RECT 632.400 499.200 633.600 499.950 ;
        RECT 613.950 496.950 616.050 499.050 ;
        RECT 616.950 496.950 619.050 499.050 ;
        RECT 610.950 460.950 613.050 463.050 ;
        RECT 610.950 454.950 613.050 457.050 ;
        RECT 611.400 450.600 612.450 454.950 ;
        RECT 614.400 454.050 615.450 496.950 ;
        RECT 613.950 451.950 616.050 454.050 ;
        RECT 617.400 450.600 618.450 496.950 ;
        RECT 627.900 495.900 630.000 497.700 ;
        RECT 631.800 496.800 633.900 498.900 ;
        RECT 635.100 498.300 637.200 500.400 ;
        RECT 626.400 494.700 635.100 495.900 ;
        RECT 623.100 490.950 625.200 493.050 ;
        RECT 623.400 489.450 624.600 490.650 ;
        RECT 620.400 488.400 624.600 489.450 ;
        RECT 620.400 481.050 621.450 488.400 ;
        RECT 626.400 485.700 627.300 494.700 ;
        RECT 633.000 493.800 635.100 494.700 ;
        RECT 636.000 492.900 636.900 498.300 ;
        RECT 638.400 495.450 639.600 495.600 ;
        RECT 641.400 495.450 642.450 512.400 ;
        RECT 643.950 511.950 646.050 514.050 ;
        RECT 644.400 496.050 645.450 511.950 ;
        RECT 674.400 508.050 675.450 529.950 ;
        RECT 680.400 528.600 681.450 532.950 ;
        RECT 683.400 532.050 684.450 565.800 ;
        RECT 686.400 556.050 687.450 607.950 ;
        RECT 689.400 600.900 690.450 614.400 ;
        RECT 703.950 613.950 706.050 616.050 ;
        RECT 697.950 610.950 700.050 613.050 ;
        RECT 698.400 606.600 699.450 610.950 ;
        RECT 704.400 606.600 705.450 613.950 ;
        RECT 707.400 610.050 708.450 634.950 ;
        RECT 710.400 625.050 711.450 637.950 ;
        RECT 712.950 634.800 715.050 636.900 ;
        RECT 709.950 622.950 712.050 625.050 ;
        RECT 713.400 619.050 714.450 634.800 ;
        RECT 716.400 634.050 717.450 691.950 ;
        RECT 719.400 685.050 720.450 691.950 ;
        RECT 725.400 691.050 726.450 721.950 ;
        RECT 727.950 718.800 730.050 720.900 ;
        RECT 728.400 712.050 729.450 718.800 ;
        RECT 727.950 709.950 730.050 712.050 ;
        RECT 731.400 694.050 732.450 781.950 ;
        RECT 733.950 763.950 736.050 766.050 ;
        RECT 730.950 691.950 733.050 694.050 ;
        RECT 721.950 689.550 726.450 691.050 ;
        RECT 721.950 688.950 726.000 689.550 ;
        RECT 718.950 682.950 721.050 685.050 ;
        RECT 721.950 684.000 724.050 687.900 ;
        RECT 727.950 684.000 730.050 688.050 ;
        RECT 734.400 684.450 735.450 763.950 ;
        RECT 737.400 763.050 738.450 790.950 ;
        RECT 740.400 766.050 741.450 814.950 ;
        RECT 743.400 793.050 744.450 823.950 ;
        RECT 745.950 806.100 748.050 808.200 ;
        RECT 746.400 802.050 747.450 806.100 ;
        RECT 745.950 799.950 748.050 802.050 ;
        RECT 742.950 790.950 745.050 793.050 ;
        RECT 749.400 790.050 750.450 827.400 ;
        RECT 755.400 811.050 756.450 859.950 ;
        RECT 757.950 847.950 760.050 850.050 ;
        RECT 758.400 817.050 759.450 847.950 ;
        RECT 761.400 847.050 762.450 868.950 ;
        RECT 767.400 862.050 768.450 884.100 ;
        RECT 770.400 868.050 771.450 889.950 ;
        RECT 773.400 874.050 774.450 907.950 ;
        RECT 776.400 892.050 777.450 922.950 ;
        RECT 779.400 892.050 780.450 931.950 ;
        RECT 785.400 918.600 786.450 931.950 ;
        RECT 785.400 916.350 786.600 918.600 ;
        RECT 790.950 917.100 793.050 919.200 ;
        RECT 791.400 916.350 792.600 917.100 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 788.400 912.900 789.600 913.650 ;
        RECT 797.400 913.050 798.450 940.950 ;
        RECT 817.950 931.950 820.050 934.050 ;
        RECT 799.950 925.950 802.050 928.050 ;
        RECT 808.950 925.950 811.050 928.050 ;
        RECT 787.950 910.800 790.050 912.900 ;
        RECT 796.950 910.950 799.050 913.050 ;
        RECT 800.400 910.050 801.450 925.950 ;
        RECT 802.950 917.100 805.050 919.200 ;
        RECT 809.400 918.600 810.450 925.950 ;
        RECT 818.400 918.600 819.450 931.950 ;
        RECT 824.400 925.050 825.450 940.950 ;
        RECT 827.400 937.050 828.450 961.950 ;
        RECT 826.950 934.950 829.050 937.050 ;
        RECT 823.950 922.950 826.050 925.050 ;
        RECT 836.400 919.200 837.450 964.950 ;
        RECT 844.950 962.100 847.050 964.200 ;
        RECT 845.400 961.350 846.600 962.100 ;
        RECT 859.950 961.950 862.050 964.050 ;
        RECT 868.950 962.100 871.050 964.200 ;
        RECT 841.950 958.950 844.050 961.050 ;
        RECT 844.950 958.950 847.050 961.050 ;
        RECT 847.950 958.950 850.050 961.050 ;
        RECT 842.400 957.900 843.600 958.650 ;
        RECT 848.400 957.900 849.600 958.650 ;
        RECT 841.950 955.800 844.050 957.900 ;
        RECT 847.950 955.800 850.050 957.900 ;
        RECT 848.400 930.450 849.450 955.800 ;
        RECT 853.950 940.950 856.050 943.050 ;
        RECT 854.400 934.050 855.450 940.950 ;
        RECT 860.400 937.050 861.450 961.950 ;
        RECT 869.400 961.350 870.600 962.100 ;
        RECT 883.950 961.950 886.050 964.050 ;
        RECT 892.950 962.100 895.050 964.200 ;
        RECT 898.950 963.000 901.050 967.050 ;
        RECT 865.950 958.950 868.050 961.050 ;
        RECT 868.950 958.950 871.050 961.050 ;
        RECT 871.950 958.950 874.050 961.050 ;
        RECT 866.400 956.400 867.600 958.650 ;
        RECT 872.400 956.400 873.600 958.650 ;
        RECT 884.400 957.900 885.450 961.950 ;
        RECT 893.400 961.350 894.600 962.100 ;
        RECT 899.400 961.350 900.600 963.000 ;
        RECT 907.950 961.950 910.050 964.050 ;
        RECT 919.950 962.100 922.050 964.200 ;
        RECT 889.950 958.950 892.050 961.050 ;
        RECT 892.950 958.950 895.050 961.050 ;
        RECT 895.950 958.950 898.050 961.050 ;
        RECT 898.950 958.950 901.050 961.050 ;
        RECT 890.400 957.900 891.600 958.650 ;
        RECT 859.950 934.950 862.050 937.050 ;
        RECT 853.950 931.950 856.050 934.050 ;
        RECT 866.400 931.050 867.450 956.400 ;
        RECT 872.400 954.450 873.450 956.400 ;
        RECT 883.950 955.800 886.050 957.900 ;
        RECT 889.950 955.800 892.050 957.900 ;
        RECT 896.400 956.400 897.600 958.650 ;
        RECT 869.400 953.400 873.450 954.450 ;
        RECT 869.400 946.050 870.450 953.400 ;
        RECT 896.400 952.050 897.450 956.400 ;
        RECT 904.950 952.950 907.050 955.050 ;
        RECT 895.950 949.950 898.050 952.050 ;
        RECT 880.950 946.950 883.050 949.050 ;
        RECT 868.950 943.950 871.050 946.050 ;
        RECT 848.400 929.400 852.450 930.450 ;
        RECT 841.950 922.950 844.050 925.050 ;
        RECT 809.400 918.450 810.600 918.600 ;
        RECT 806.400 917.400 810.600 918.450 ;
        RECT 799.950 907.950 802.050 910.050 ;
        RECT 793.950 892.950 796.050 895.050 ;
        RECT 775.950 889.950 778.050 892.050 ;
        RECT 778.950 889.950 781.050 892.050 ;
        RECT 787.950 889.950 790.050 892.050 ;
        RECT 781.950 884.100 784.050 886.200 ;
        RECT 788.400 885.600 789.450 889.950 ;
        RECT 782.400 883.350 783.600 884.100 ;
        RECT 788.400 883.350 789.600 885.600 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 779.400 878.400 780.600 880.650 ;
        RECT 785.400 879.900 786.600 880.650 ;
        RECT 772.950 871.950 775.050 874.050 ;
        RECT 779.400 868.050 780.450 878.400 ;
        RECT 784.950 874.950 787.050 879.900 ;
        RECT 794.400 877.050 795.450 892.950 ;
        RECT 796.950 886.950 799.050 889.050 ;
        RECT 790.800 874.950 792.900 877.050 ;
        RECT 793.950 874.950 796.050 877.050 ;
        RECT 787.950 871.950 790.050 874.050 ;
        RECT 769.950 865.950 772.050 868.050 ;
        RECT 778.950 865.950 781.050 868.050 ;
        RECT 766.950 859.950 769.050 862.050 ;
        RECT 760.950 844.950 763.050 847.050 ;
        RECT 772.950 844.950 775.050 847.050 ;
        RECT 766.950 839.100 769.050 841.200 ;
        RECT 773.400 840.600 774.450 844.950 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 757.950 814.950 760.050 817.050 ;
        RECT 761.400 814.050 762.450 835.950 ;
        RECT 767.400 826.050 768.450 839.100 ;
        RECT 773.400 838.350 774.600 840.600 ;
        RECT 778.950 839.100 781.050 841.200 ;
        RECT 779.400 838.350 780.600 839.100 ;
        RECT 772.950 835.950 775.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 776.400 834.900 777.600 835.650 ;
        RECT 769.950 831.450 772.050 834.900 ;
        RECT 775.950 832.800 778.050 834.900 ;
        RECT 782.400 834.000 783.600 835.650 ;
        RECT 769.950 831.000 774.450 831.450 ;
        RECT 770.400 830.400 774.450 831.000 ;
        RECT 769.950 826.950 772.050 829.050 ;
        RECT 766.950 823.950 769.050 826.050 ;
        RECT 760.950 811.950 763.050 814.050 ;
        RECT 754.950 808.950 757.050 811.050 ;
        RECT 755.400 807.600 756.450 808.950 ;
        RECT 755.400 805.350 756.600 807.600 ;
        RECT 760.950 806.100 763.050 808.200 ;
        RECT 761.400 805.350 762.600 806.100 ;
        RECT 770.400 805.050 771.450 826.950 ;
        RECT 773.400 817.050 774.450 830.400 ;
        RECT 776.400 829.050 777.450 832.800 ;
        RECT 781.950 829.950 784.050 834.000 ;
        RECT 788.400 832.050 789.450 871.950 ;
        RECT 791.400 838.050 792.450 874.950 ;
        RECT 797.400 868.050 798.450 886.950 ;
        RECT 803.400 886.050 804.450 917.100 ;
        RECT 806.400 907.050 807.450 917.400 ;
        RECT 809.400 916.350 810.600 917.400 ;
        RECT 818.400 916.350 819.600 918.600 ;
        RECT 826.950 916.950 829.050 919.050 ;
        RECT 835.950 917.100 838.050 919.200 ;
        RECT 842.400 918.600 843.450 922.950 ;
        RECT 809.100 913.950 811.200 916.050 ;
        RECT 814.500 913.950 816.600 916.050 ;
        RECT 817.800 913.950 819.900 916.050 ;
        RECT 815.400 911.400 816.600 913.650 ;
        RECT 815.400 907.050 816.450 911.400 ;
        RECT 823.950 907.950 826.050 910.050 ;
        RECT 805.950 904.950 808.050 907.050 ;
        RECT 814.950 904.950 817.050 907.050 ;
        RECT 802.950 883.950 805.050 886.050 ;
        RECT 808.950 884.100 811.050 886.200 ;
        RECT 815.400 885.600 816.450 904.950 ;
        RECT 809.400 883.350 810.600 884.100 ;
        RECT 815.400 883.350 816.600 885.600 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 799.950 877.950 802.050 880.050 ;
        RECT 806.400 878.400 807.600 880.650 ;
        RECT 812.400 878.400 813.600 880.650 ;
        RECT 800.400 871.050 801.450 877.950 ;
        RECT 806.400 877.050 807.450 878.400 ;
        RECT 805.950 871.950 808.050 877.050 ;
        RECT 812.400 871.050 813.450 878.400 ;
        RECT 799.950 868.950 802.050 871.050 ;
        RECT 811.950 868.950 814.050 871.050 ;
        RECT 793.800 865.950 796.050 868.050 ;
        RECT 796.950 865.950 799.050 868.050 ;
        RECT 799.950 862.950 802.050 867.900 ;
        RECT 793.950 853.950 796.050 856.050 ;
        RECT 790.950 835.950 793.050 838.050 ;
        RECT 794.400 834.450 795.450 853.950 ;
        RECT 824.400 853.050 825.450 907.950 ;
        RECT 827.400 877.050 828.450 916.950 ;
        RECT 836.400 916.350 837.600 917.100 ;
        RECT 842.400 916.350 843.600 918.600 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 838.950 913.950 841.050 916.050 ;
        RECT 841.950 913.950 844.050 916.050 ;
        RECT 844.950 913.950 847.050 916.050 ;
        RECT 839.400 911.400 840.600 913.650 ;
        RECT 845.400 912.900 846.600 913.650 ;
        RECT 835.950 898.950 838.050 901.050 ;
        RECT 836.400 889.200 837.450 898.950 ;
        RECT 839.400 895.050 840.450 911.400 ;
        RECT 844.950 910.800 847.050 912.900 ;
        RECT 841.950 901.950 844.050 904.050 ;
        RECT 838.950 892.950 841.050 895.050 ;
        RECT 835.950 887.100 838.050 889.200 ;
        RECT 835.950 883.950 838.050 886.050 ;
        RECT 842.400 885.600 843.450 901.950 ;
        RECT 847.950 894.450 850.050 895.050 ;
        RECT 851.400 894.450 852.450 929.400 ;
        RECT 865.950 928.950 868.050 931.050 ;
        RECT 856.950 925.950 859.050 928.050 ;
        RECT 853.950 916.950 856.050 919.050 ;
        RECT 854.400 907.050 855.450 916.950 ;
        RECT 857.400 912.900 858.450 925.950 ;
        RECT 869.400 919.200 870.450 943.950 ;
        RECT 877.950 928.950 880.050 931.050 ;
        RECT 859.950 918.600 864.000 919.050 ;
        RECT 859.950 916.950 864.600 918.600 ;
        RECT 868.950 917.100 871.050 919.200 ;
        RECT 863.400 916.350 864.600 916.950 ;
        RECT 869.400 916.350 870.600 917.100 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 865.950 913.950 868.050 916.050 ;
        RECT 868.950 913.950 871.050 916.050 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 866.400 912.900 867.600 913.650 ;
        RECT 856.950 910.800 859.050 912.900 ;
        RECT 865.950 910.800 868.050 912.900 ;
        RECT 872.400 911.400 873.600 913.650 ;
        RECT 872.400 907.050 873.450 911.400 ;
        RECT 853.950 904.950 856.050 907.050 ;
        RECT 871.950 904.950 874.050 907.050 ;
        RECT 878.400 904.050 879.450 928.950 ;
        RECT 877.950 901.950 880.050 904.050 ;
        RECT 881.400 898.050 882.450 946.950 ;
        RECT 883.950 934.950 886.050 937.050 ;
        RECT 884.400 912.900 885.450 934.950 ;
        RECT 905.400 925.050 906.450 952.950 ;
        RECT 889.950 922.950 892.050 925.050 ;
        RECT 904.950 922.950 907.050 925.050 ;
        RECT 890.400 918.600 891.450 922.950 ;
        RECT 908.400 922.050 909.450 961.950 ;
        RECT 920.400 961.350 921.600 962.100 ;
        RECT 931.800 961.950 933.900 964.050 ;
        RECT 934.950 962.100 937.050 964.200 ;
        RECT 943.950 962.100 946.050 964.200 ;
        RECT 950.400 963.600 951.450 967.950 ;
        RECT 916.950 958.950 919.050 961.050 ;
        RECT 919.950 958.950 922.050 961.050 ;
        RECT 922.950 958.950 925.050 961.050 ;
        RECT 917.400 956.400 918.600 958.650 ;
        RECT 923.400 957.000 924.600 958.650 ;
        RECT 932.400 957.900 933.450 961.950 ;
        RECT 917.400 937.050 918.450 956.400 ;
        RECT 922.950 952.950 925.050 957.000 ;
        RECT 931.950 955.800 934.050 957.900 ;
        RECT 935.400 946.050 936.450 962.100 ;
        RECT 944.400 961.350 945.600 962.100 ;
        RECT 950.400 961.350 951.600 963.600 ;
        RECT 970.950 963.000 973.050 967.050 ;
        RECT 974.400 964.050 975.450 968.400 ;
        RECT 979.950 964.950 982.050 967.050 ;
        RECT 971.400 961.350 972.600 963.000 ;
        RECT 973.950 961.950 976.050 964.050 ;
        RECT 940.950 958.950 943.050 961.050 ;
        RECT 943.950 958.950 946.050 961.050 ;
        RECT 946.950 958.950 949.050 961.050 ;
        RECT 949.950 958.950 952.050 961.050 ;
        RECT 967.950 958.950 970.050 961.050 ;
        RECT 970.950 958.950 973.050 961.050 ;
        RECT 941.400 957.900 942.600 958.650 ;
        RECT 940.950 955.800 943.050 957.900 ;
        RECT 947.400 956.400 948.600 958.650 ;
        RECT 968.400 957.000 969.600 958.650 ;
        RECT 934.950 943.950 937.050 946.050 ;
        RECT 947.400 940.050 948.450 956.400 ;
        RECT 955.950 952.950 958.050 955.050 ;
        RECT 967.950 952.950 970.050 957.000 ;
        RECT 946.950 937.950 949.050 940.050 ;
        RECT 916.950 934.950 919.050 937.050 ;
        RECT 907.950 919.950 910.050 922.050 ;
        RECT 890.400 916.350 891.600 918.600 ;
        RECT 895.950 917.100 898.050 919.200 ;
        RECT 904.950 917.100 907.050 919.200 ;
        RECT 910.950 917.100 913.050 919.200 ;
        RECT 916.950 918.000 919.050 922.050 ;
        RECT 952.950 919.950 955.050 922.050 ;
        RECT 896.400 916.350 897.600 917.100 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 892.950 913.950 895.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 893.400 912.900 894.600 913.650 ;
        RECT 883.950 910.800 886.050 912.900 ;
        RECT 892.950 910.800 895.050 912.900 ;
        RECT 899.400 911.400 900.600 913.650 ;
        RECT 892.950 898.950 895.050 901.050 ;
        RECT 859.950 895.950 862.050 898.050 ;
        RECT 880.950 895.950 883.050 898.050 ;
        RECT 847.950 893.400 852.450 894.450 ;
        RECT 847.950 892.950 850.050 893.400 ;
        RECT 836.400 883.350 837.600 883.950 ;
        RECT 842.400 883.350 843.600 885.600 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 838.950 880.950 841.050 883.050 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 833.400 878.400 834.600 880.650 ;
        RECT 839.400 878.400 840.600 880.650 ;
        RECT 826.950 874.950 829.050 877.050 ;
        RECT 823.950 850.950 826.050 853.050 ;
        RECT 827.400 850.050 828.450 874.950 ;
        RECT 833.400 871.050 834.450 878.400 ;
        RECT 839.400 874.050 840.450 878.400 ;
        RECT 838.950 871.950 841.050 874.050 ;
        RECT 832.950 868.950 835.050 871.050 ;
        RECT 833.400 850.050 834.450 868.950 ;
        RECT 839.400 856.050 840.450 871.950 ;
        RECT 844.950 862.950 847.050 865.050 ;
        RECT 838.950 853.950 841.050 856.050 ;
        RECT 826.950 847.950 829.050 850.050 ;
        RECT 832.950 847.950 835.050 850.050 ;
        RECT 841.950 847.950 844.050 850.050 ;
        RECT 805.950 844.950 808.050 847.050 ;
        RECT 806.400 841.200 807.450 844.950 ;
        RECT 820.950 841.950 823.050 844.050 ;
        RECT 799.950 839.100 802.050 841.200 ;
        RECT 805.950 839.100 808.050 841.200 ;
        RECT 814.950 839.100 817.050 841.200 ;
        RECT 800.400 838.350 801.600 839.100 ;
        RECT 806.400 838.350 807.600 839.100 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 805.950 835.950 808.050 838.050 ;
        RECT 808.950 835.950 811.050 838.050 ;
        RECT 794.400 833.400 798.450 834.450 ;
        RECT 787.800 829.950 789.900 832.050 ;
        RECT 790.950 829.950 793.050 832.050 ;
        RECT 775.950 826.950 778.050 829.050 ;
        RECT 781.950 820.950 784.050 823.050 ;
        RECT 772.950 814.950 775.050 817.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 763.950 802.950 766.050 805.050 ;
        RECT 769.950 802.950 772.050 805.050 ;
        RECT 758.400 801.900 759.600 802.650 ;
        RECT 757.950 799.800 760.050 801.900 ;
        RECT 764.400 800.400 765.600 802.650 ;
        RECT 748.950 787.950 751.050 790.050 ;
        RECT 757.950 787.950 760.050 790.050 ;
        RECT 748.950 772.950 751.050 775.050 ;
        RECT 739.950 763.950 742.050 766.050 ;
        RECT 736.950 760.950 739.050 763.050 ;
        RECT 742.950 761.100 745.050 763.200 ;
        RECT 749.400 763.050 750.450 772.950 ;
        RECT 758.400 769.050 759.450 787.950 ;
        RECT 764.400 772.050 765.450 800.400 ;
        RECT 766.950 790.950 769.050 793.050 ;
        RECT 763.950 769.950 766.050 772.050 ;
        RECT 757.950 766.950 760.050 769.050 ;
        RECT 743.400 760.350 744.600 761.100 ;
        RECT 748.950 760.950 751.050 763.050 ;
        RECT 751.950 760.950 754.050 763.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 740.400 756.900 741.600 757.650 ;
        RECT 739.950 754.800 742.050 756.900 ;
        RECT 746.400 755.400 747.600 757.650 ;
        RECT 736.950 742.950 739.050 745.050 ;
        RECT 737.400 727.050 738.450 742.950 ;
        RECT 739.950 739.950 742.050 742.050 ;
        RECT 740.400 730.050 741.450 739.950 ;
        RECT 746.400 739.050 747.450 755.400 ;
        RECT 745.950 736.950 748.050 739.050 ;
        RECT 739.950 727.950 742.050 730.050 ;
        RECT 742.950 729.000 745.050 733.050 ;
        RECT 752.400 732.450 753.450 760.950 ;
        RECT 754.950 757.950 757.050 760.050 ;
        RECT 755.400 751.050 756.450 757.950 ;
        RECT 754.950 748.950 757.050 751.050 ;
        RECT 758.400 741.450 759.450 766.950 ;
        RECT 767.400 762.600 768.450 790.950 ;
        RECT 769.950 784.950 772.050 787.050 ;
        RECT 770.400 766.050 771.450 784.950 ;
        RECT 773.400 784.050 774.450 814.950 ;
        RECT 775.950 806.100 778.050 808.200 ;
        RECT 782.400 807.600 783.450 820.950 ;
        RECT 791.400 814.050 792.450 829.950 ;
        RECT 793.950 826.950 796.050 829.050 ;
        RECT 790.950 811.950 793.050 814.050 ;
        RECT 776.400 796.050 777.450 806.100 ;
        RECT 782.400 805.350 783.600 807.600 ;
        RECT 787.950 806.100 790.050 808.200 ;
        RECT 794.400 808.050 795.450 826.950 ;
        RECT 788.400 805.350 789.600 806.100 ;
        RECT 793.950 805.950 796.050 808.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 785.400 801.900 786.600 802.650 ;
        RECT 784.950 799.800 787.050 801.900 ;
        RECT 791.400 801.000 792.600 802.650 ;
        RECT 797.400 801.450 798.450 833.400 ;
        RECT 803.400 833.400 804.600 835.650 ;
        RECT 809.400 834.900 810.600 835.650 ;
        RECT 803.400 829.050 804.450 833.400 ;
        RECT 808.950 832.800 811.050 834.900 ;
        RECT 802.950 826.950 805.050 829.050 ;
        RECT 799.950 823.950 802.050 826.050 ;
        RECT 800.400 817.050 801.450 823.950 ;
        RECT 815.400 820.050 816.450 839.100 ;
        RECT 821.400 826.050 822.450 841.950 ;
        RECT 826.950 840.000 829.050 844.050 ;
        RECT 827.400 838.350 828.600 840.000 ;
        RECT 832.950 839.100 835.050 841.200 ;
        RECT 833.400 838.350 834.600 839.100 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 829.950 835.950 832.050 838.050 ;
        RECT 832.950 835.950 835.050 838.050 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 830.400 834.900 831.600 835.650 ;
        RECT 829.950 832.800 832.050 834.900 ;
        RECT 836.400 833.400 837.600 835.650 ;
        RECT 842.400 835.050 843.450 847.950 ;
        RECT 845.400 835.050 846.450 862.950 ;
        RECT 826.950 829.950 829.050 832.050 ;
        RECT 820.950 823.950 823.050 826.050 ;
        RECT 817.950 820.950 820.050 823.050 ;
        RECT 802.950 817.950 805.050 820.050 ;
        RECT 814.950 817.950 817.050 820.050 ;
        RECT 799.950 814.950 802.050 817.050 ;
        RECT 803.400 813.450 804.450 817.950 ;
        RECT 818.400 817.050 819.450 820.950 ;
        RECT 820.950 817.950 823.050 820.050 ;
        RECT 817.950 814.950 820.050 817.050 ;
        RECT 821.400 813.450 822.450 817.950 ;
        RECT 827.400 814.050 828.450 829.950 ;
        RECT 829.950 817.950 832.050 820.050 ;
        RECT 775.950 793.950 778.050 796.050 ;
        RECT 785.400 790.050 786.450 799.800 ;
        RECT 790.950 796.950 793.050 801.000 ;
        RECT 794.400 800.400 798.450 801.450 ;
        RECT 800.400 812.400 804.450 813.450 ;
        RECT 818.400 812.400 822.450 813.450 ;
        RECT 787.950 793.950 790.050 796.050 ;
        RECT 784.950 787.950 787.050 790.050 ;
        RECT 772.950 781.950 775.050 784.050 ;
        RECT 778.950 781.950 781.050 784.050 ;
        RECT 769.950 763.950 772.050 766.050 ;
        RECT 767.400 760.350 768.600 762.600 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 760.950 754.950 763.050 757.050 ;
        RECT 764.400 756.900 765.600 757.650 ;
        RECT 773.400 757.050 774.450 781.950 ;
        RECT 749.400 731.400 753.450 732.450 ;
        RECT 755.400 740.400 759.450 741.450 ;
        RECT 749.400 729.600 750.450 731.400 ;
        RECT 755.400 730.050 756.450 740.400 ;
        RECT 757.950 733.950 760.050 739.050 ;
        RECT 743.400 727.350 744.600 729.000 ;
        RECT 749.400 727.350 750.600 729.600 ;
        RECT 754.950 727.950 757.050 730.050 ;
        RECT 757.950 727.950 760.050 730.050 ;
        RECT 736.950 724.950 739.050 727.050 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 746.400 723.900 747.600 724.650 ;
        RECT 752.400 724.050 753.600 724.650 ;
        RECT 736.800 721.800 738.900 723.900 ;
        RECT 737.400 712.050 738.450 721.800 ;
        RECT 739.950 718.950 742.050 723.900 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 752.400 722.400 757.050 724.050 ;
        RECT 753.000 721.950 757.050 722.400 ;
        RECT 758.400 718.050 759.450 727.950 ;
        RECT 761.400 724.050 762.450 754.950 ;
        RECT 763.950 754.800 766.050 756.900 ;
        RECT 772.950 754.950 775.050 757.050 ;
        RECT 766.950 736.950 769.050 739.050 ;
        RECT 763.950 730.950 766.050 733.050 ;
        RECT 760.950 721.950 763.050 724.050 ;
        RECT 757.950 715.950 760.050 718.050 ;
        RECT 739.950 712.950 742.050 715.050 ;
        RECT 745.950 712.950 748.050 715.050 ;
        RECT 736.950 709.950 739.050 712.050 ;
        RECT 740.400 709.050 741.450 712.950 ;
        RECT 739.950 706.950 742.050 709.050 ;
        RECT 736.950 697.950 739.050 703.050 ;
        RECT 742.950 700.950 745.050 703.050 ;
        RECT 739.950 685.950 742.050 688.050 ;
        RECT 722.400 682.350 723.600 684.000 ;
        RECT 728.400 682.350 729.600 684.000 ;
        RECT 734.400 683.400 738.450 684.450 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 718.950 676.950 721.050 679.050 ;
        RECT 725.400 677.400 726.600 679.650 ;
        RECT 731.400 678.900 732.600 679.650 ;
        RECT 715.950 631.950 718.050 634.050 ;
        RECT 712.950 616.950 715.050 619.050 ;
        RECT 706.950 607.950 709.050 610.050 ;
        RECT 712.950 607.950 715.050 610.050 ;
        RECT 698.400 604.350 699.600 606.600 ;
        RECT 704.400 604.350 705.600 606.600 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 697.950 601.950 700.050 604.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 695.400 600.900 696.600 601.650 ;
        RECT 688.950 595.950 691.050 600.900 ;
        RECT 694.950 598.800 697.050 600.900 ;
        RECT 701.400 599.400 702.600 601.650 ;
        RECT 707.400 600.000 708.600 601.650 ;
        RECT 713.400 601.050 714.450 607.950 ;
        RECT 691.950 592.950 694.050 595.050 ;
        RECT 688.950 580.950 691.050 583.050 ;
        RECT 689.400 562.050 690.450 580.950 ;
        RECT 692.400 574.050 693.450 592.950 ;
        RECT 695.400 577.050 696.450 598.800 ;
        RECT 694.950 574.950 697.050 577.050 ;
        RECT 701.400 576.450 702.450 599.400 ;
        RECT 706.950 595.950 709.050 600.000 ;
        RECT 712.950 598.950 715.050 601.050 ;
        RECT 712.950 595.800 715.050 597.900 ;
        RECT 713.400 589.050 714.450 595.800 ;
        RECT 712.950 586.950 715.050 589.050 ;
        RECT 701.400 575.400 705.450 576.450 ;
        RECT 691.950 571.950 694.050 574.050 ;
        RECT 697.950 572.100 700.050 574.200 ;
        RECT 704.400 573.600 705.450 575.400 ;
        RECT 712.950 574.950 715.050 577.050 ;
        RECT 698.400 571.350 699.600 572.100 ;
        RECT 704.400 571.350 705.600 573.600 ;
        RECT 709.950 571.950 712.050 574.050 ;
        RECT 694.950 568.950 697.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 695.400 567.900 696.600 568.650 ;
        RECT 701.400 567.900 702.600 568.650 ;
        RECT 694.950 565.800 697.050 567.900 ;
        RECT 700.950 565.800 703.050 567.900 ;
        RECT 688.950 559.950 691.050 562.050 ;
        RECT 694.950 559.950 697.050 562.050 ;
        RECT 685.950 553.950 688.050 556.050 ;
        RECT 691.950 550.950 694.050 553.050 ;
        RECT 692.400 541.050 693.450 550.950 ;
        RECT 691.950 538.950 694.050 541.050 ;
        RECT 695.400 532.050 696.450 559.950 ;
        RECT 710.400 559.050 711.450 571.950 ;
        RECT 713.400 565.050 714.450 574.950 ;
        RECT 712.950 562.950 715.050 565.050 ;
        RECT 709.950 556.950 712.050 559.050 ;
        RECT 700.950 553.950 703.050 556.050 ;
        RECT 697.950 541.950 700.050 544.050 ;
        RECT 682.950 529.950 685.050 532.050 ;
        RECT 680.400 526.350 681.600 528.600 ;
        RECT 685.950 528.000 688.050 532.050 ;
        RECT 694.950 529.950 697.050 532.050 ;
        RECT 686.400 526.350 687.600 528.000 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 694.950 523.950 697.050 526.050 ;
        RECT 676.950 520.950 679.050 523.050 ;
        RECT 683.400 521.400 684.600 523.650 ;
        RECT 689.400 521.400 690.600 523.650 ;
        RECT 677.400 508.050 678.450 520.950 ;
        RECT 683.400 514.050 684.450 521.400 ;
        RECT 689.400 517.050 690.450 521.400 ;
        RECT 688.950 514.950 691.050 517.050 ;
        RECT 682.950 511.950 685.050 514.050 ;
        RECT 695.400 508.050 696.450 523.950 ;
        RECT 698.400 523.050 699.450 541.950 ;
        RECT 697.950 520.950 700.050 523.050 ;
        RECT 701.400 522.450 702.450 553.950 ;
        RECT 706.950 550.950 709.050 553.050 ;
        RECT 703.950 547.950 706.050 550.050 ;
        RECT 704.400 544.050 705.450 547.950 ;
        RECT 703.950 541.950 706.050 544.050 ;
        RECT 707.400 541.050 708.450 550.950 ;
        RECT 709.950 547.950 712.050 550.050 ;
        RECT 710.400 544.050 711.450 547.950 ;
        RECT 709.950 541.950 712.050 544.050 ;
        RECT 703.950 538.800 706.050 540.900 ;
        RECT 706.950 538.950 709.050 541.050 ;
        RECT 716.400 540.450 717.450 631.950 ;
        RECT 719.400 628.050 720.450 676.950 ;
        RECT 725.400 667.050 726.450 677.400 ;
        RECT 730.950 676.800 733.050 678.900 ;
        RECT 733.950 673.950 736.050 676.050 ;
        RECT 733.950 670.800 736.050 672.900 ;
        RECT 734.400 667.050 735.450 670.800 ;
        RECT 721.800 664.950 723.900 667.050 ;
        RECT 724.950 664.950 727.050 667.050 ;
        RECT 733.950 664.950 736.050 667.050 ;
        RECT 722.400 661.050 723.450 664.950 ;
        RECT 722.400 659.400 727.050 661.050 ;
        RECT 723.000 658.950 727.050 659.400 ;
        RECT 733.950 658.950 736.050 661.050 ;
        RECT 721.950 655.950 724.050 658.050 ;
        RECT 722.400 652.050 723.450 655.950 ;
        RECT 721.950 649.950 724.050 652.050 ;
        RECT 727.950 651.000 730.050 655.050 ;
        RECT 734.400 651.600 735.450 658.950 ;
        RECT 737.400 658.050 738.450 683.400 ;
        RECT 740.400 673.050 741.450 685.950 ;
        RECT 743.400 682.050 744.450 700.950 ;
        RECT 746.400 700.050 747.450 712.950 ;
        RECT 745.950 697.950 748.050 700.050 ;
        RECT 760.950 697.950 763.050 700.050 ;
        RECT 757.950 694.950 760.050 697.050 ;
        RECT 745.950 685.950 748.050 691.050 ;
        RECT 751.950 683.100 754.050 685.200 ;
        RECT 758.400 684.600 759.450 694.950 ;
        RECT 761.400 685.050 762.450 697.950 ;
        RECT 752.400 682.350 753.600 683.100 ;
        RECT 758.400 682.350 759.600 684.600 ;
        RECT 760.950 682.950 763.050 685.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 751.950 679.950 754.050 682.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 749.400 678.450 750.600 679.650 ;
        RECT 746.400 677.400 750.600 678.450 ;
        RECT 755.400 677.400 756.600 679.650 ;
        RECT 742.950 673.950 745.050 676.050 ;
        RECT 739.950 670.950 742.050 673.050 ;
        RECT 743.400 670.050 744.450 673.950 ;
        RECT 746.400 673.050 747.450 677.400 ;
        RECT 745.950 670.950 748.050 673.050 ;
        RECT 755.400 670.050 756.450 677.400 ;
        RECT 739.800 669.000 741.900 669.900 ;
        RECT 739.800 667.800 742.050 669.000 ;
        RECT 742.950 667.950 745.050 670.050 ;
        RECT 754.950 667.950 757.050 670.050 ;
        RECT 739.950 666.450 742.050 667.800 ;
        RECT 739.950 666.000 747.450 666.450 ;
        RECT 740.400 665.400 747.450 666.000 ;
        RECT 742.950 661.950 745.050 664.050 ;
        RECT 739.950 658.950 742.050 661.050 ;
        RECT 736.950 655.950 739.050 658.050 ;
        RECT 740.400 655.050 741.450 658.950 ;
        RECT 738.000 654.900 741.450 655.050 ;
        RECT 736.950 653.400 741.450 654.900 ;
        RECT 736.950 652.950 741.000 653.400 ;
        RECT 736.950 652.800 739.050 652.950 ;
        RECT 743.400 652.050 744.450 661.950 ;
        RECT 746.400 655.050 747.450 665.400 ;
        RECT 748.950 661.950 751.050 664.050 ;
        RECT 760.950 661.950 763.050 664.050 ;
        RECT 745.950 652.950 748.050 655.050 ;
        RECT 728.400 649.350 729.600 651.000 ;
        RECT 734.400 649.350 735.600 651.600 ;
        RECT 742.950 649.950 745.050 652.050 ;
        RECT 745.950 649.800 748.050 651.900 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 725.400 645.900 726.600 646.650 ;
        RECT 724.950 643.800 727.050 645.900 ;
        RECT 731.400 644.400 732.600 646.650 ;
        RECT 737.400 645.000 738.600 646.650 ;
        RECT 724.950 642.300 727.050 642.750 ;
        RECT 731.400 642.300 732.450 644.400 ;
        RECT 724.950 641.250 732.450 642.300 ;
        RECT 724.950 640.650 727.050 641.250 ;
        RECT 736.950 640.950 739.050 645.000 ;
        RECT 721.950 637.950 724.050 640.050 ;
        RECT 718.950 625.950 721.050 628.050 ;
        RECT 722.400 622.050 723.450 637.950 ;
        RECT 727.950 625.950 730.050 628.050 ;
        RECT 721.950 619.950 724.050 622.050 ;
        RECT 722.400 606.450 723.450 619.950 ;
        RECT 728.400 610.050 729.450 625.950 ;
        RECT 736.950 613.950 739.050 616.050 ;
        RECT 719.400 605.400 723.450 606.450 ;
        RECT 724.950 606.000 727.050 610.050 ;
        RECT 727.950 607.950 730.050 610.050 ;
        RECT 719.400 598.050 720.450 605.400 ;
        RECT 725.400 604.350 726.600 606.000 ;
        RECT 730.950 605.100 733.050 607.200 ;
        RECT 737.400 606.600 738.450 613.950 ;
        RECT 731.400 604.350 732.600 605.100 ;
        RECT 737.400 604.350 738.600 606.600 ;
        RECT 742.950 604.950 745.050 607.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 721.950 598.800 724.050 601.050 ;
        RECT 728.400 600.900 729.600 601.650 ;
        RECT 727.950 598.800 730.050 600.900 ;
        RECT 734.400 600.000 735.600 601.650 ;
        RECT 718.950 595.950 721.050 598.050 ;
        RECT 727.950 595.650 730.050 597.750 ;
        RECT 733.950 595.950 736.050 600.000 ;
        RECT 718.800 589.950 720.900 592.050 ;
        RECT 721.950 589.950 724.050 595.050 ;
        RECT 719.400 577.050 720.450 589.950 ;
        RECT 728.400 583.050 729.450 595.650 ;
        RECT 733.950 592.800 736.050 594.900 ;
        RECT 727.950 580.950 730.050 583.050 ;
        RECT 718.950 574.950 721.050 577.050 ;
        RECT 724.950 572.100 727.050 574.200 ;
        RECT 725.400 571.350 726.600 572.100 ;
        RECT 722.100 568.950 724.200 571.050 ;
        RECT 725.400 568.950 727.500 571.050 ;
        RECT 730.800 568.950 732.900 571.050 ;
        RECT 722.400 567.900 723.600 568.650 ;
        RECT 731.400 567.900 732.600 568.650 ;
        RECT 721.950 565.800 724.050 567.900 ;
        RECT 730.950 565.800 733.050 567.900 ;
        RECT 724.950 562.950 727.050 565.050 ;
        RECT 716.400 539.400 720.450 540.450 ;
        RECT 704.400 529.050 705.450 538.800 ;
        RECT 715.950 535.950 718.050 538.050 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 709.950 527.100 712.050 529.200 ;
        RECT 716.400 528.600 717.450 535.950 ;
        RECT 719.400 535.050 720.450 539.400 ;
        RECT 718.950 532.950 721.050 535.050 ;
        RECT 718.950 529.800 721.050 531.900 ;
        RECT 710.400 526.350 711.600 527.100 ;
        RECT 716.400 526.350 717.600 528.600 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 707.400 522.900 708.600 523.650 ;
        RECT 701.400 521.400 705.450 522.450 ;
        RECT 697.950 517.800 700.050 519.900 ;
        RECT 652.950 505.950 655.050 508.050 ;
        RECT 670.950 506.400 675.450 508.050 ;
        RECT 670.950 505.950 675.000 506.400 ;
        RECT 676.950 505.950 679.050 508.050 ;
        RECT 694.950 505.950 697.050 508.050 ;
        RECT 638.400 494.400 642.450 495.450 ;
        RECT 638.400 493.350 639.600 494.400 ;
        RECT 643.950 493.950 646.050 496.050 ;
        RECT 630.000 491.700 636.900 492.900 ;
        RECT 630.000 489.300 630.900 491.700 ;
        RECT 628.800 487.200 630.900 489.300 ;
        RECT 631.800 487.950 633.900 490.050 ;
        RECT 625.500 483.600 627.600 485.700 ;
        RECT 632.400 485.400 633.600 487.650 ;
        RECT 635.700 484.500 636.900 491.700 ;
        RECT 637.800 490.950 639.900 493.050 ;
        RECT 643.800 487.950 645.900 490.050 ;
        RECT 649.800 487.950 651.900 490.050 ;
        RECT 644.400 485.400 645.600 487.650 ;
        RECT 635.100 482.400 637.200 484.500 ;
        RECT 619.950 478.950 622.050 481.050 ;
        RECT 625.950 472.950 628.050 475.050 ;
        RECT 611.400 448.350 612.600 450.600 ;
        RECT 617.400 448.350 618.600 450.600 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 614.400 443.400 615.600 445.650 ;
        RECT 620.400 444.900 621.600 445.650 ;
        RECT 610.950 433.950 613.050 436.050 ;
        RECT 599.400 415.350 600.600 417.000 ;
        RECT 605.400 415.350 606.600 417.600 ;
        RECT 607.950 415.950 610.050 421.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 596.400 410.400 597.600 412.650 ;
        RECT 602.400 410.400 603.600 412.650 ;
        RECT 596.400 403.050 597.450 410.400 ;
        RECT 595.950 400.950 598.050 403.050 ;
        RECT 602.400 391.050 603.450 410.400 ;
        RECT 601.950 388.950 604.050 391.050 ;
        RECT 592.950 385.950 595.050 388.050 ;
        RECT 593.400 364.050 594.450 385.950 ;
        RECT 601.950 372.000 604.050 376.050 ;
        RECT 602.400 370.350 603.600 372.000 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 599.400 366.900 600.600 367.650 ;
        RECT 605.400 366.900 606.600 367.650 ;
        RECT 611.400 366.900 612.450 433.950 ;
        RECT 614.400 433.050 615.450 443.400 ;
        RECT 619.950 442.800 622.050 444.900 ;
        RECT 613.950 430.950 616.050 433.050 ;
        RECT 626.400 424.050 627.450 472.950 ;
        RECT 644.400 466.050 645.450 485.400 ;
        RECT 646.950 484.950 649.050 487.050 ;
        RECT 643.950 463.950 646.050 466.050 ;
        RECT 631.950 454.950 634.050 457.050 ;
        RECT 632.400 433.050 633.450 454.950 ;
        RECT 647.400 454.050 648.450 484.950 ;
        RECT 649.950 481.950 652.050 484.050 ;
        RECT 646.950 451.950 649.050 454.050 ;
        RECT 640.950 449.100 643.050 451.200 ;
        RECT 641.400 448.350 642.600 449.100 ;
        RECT 646.950 448.800 649.050 450.900 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 638.400 444.900 639.600 445.650 ;
        RECT 647.400 444.900 648.450 448.800 ;
        RECT 637.950 442.800 640.050 444.900 ;
        RECT 646.950 442.800 649.050 444.900 ;
        RECT 650.400 436.050 651.450 481.950 ;
        RECT 653.400 475.050 654.450 505.950 ;
        RECT 656.700 501.300 658.800 503.400 ;
        RECT 659.700 501.300 661.800 503.400 ;
        RECT 662.700 501.300 664.800 503.400 ;
        RECT 657.300 497.700 658.500 501.300 ;
        RECT 656.400 495.600 658.500 497.700 ;
        RECT 656.400 476.700 657.900 495.600 ;
        RECT 660.300 484.800 661.500 501.300 ;
        RECT 659.400 482.700 661.500 484.800 ;
        RECT 660.300 476.700 661.500 482.700 ;
        RECT 662.700 479.700 663.900 501.300 ;
        RECT 670.800 500.400 672.900 502.500 ;
        RECT 676.200 501.300 678.300 503.400 ;
        RECT 679.200 501.300 681.300 503.400 ;
        RECT 682.200 501.300 684.300 503.400 ;
        RECT 667.800 493.950 669.900 496.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 668.400 491.400 669.600 493.650 ;
        RECT 665.400 484.050 666.450 490.950 ;
        RECT 664.950 481.950 667.050 484.050 ;
        RECT 662.700 477.600 664.800 479.700 ;
        RECT 652.950 472.950 655.050 475.050 ;
        RECT 656.400 474.600 659.400 476.700 ;
        RECT 660.300 474.600 662.400 476.700 ;
        RECT 668.400 472.050 669.450 491.400 ;
        RECT 671.400 489.900 672.300 500.400 ;
        RECT 674.100 494.400 676.200 496.500 ;
        RECT 671.400 487.800 673.500 489.900 ;
        RECT 677.100 489.000 678.300 501.300 ;
        RECT 671.400 481.200 672.300 487.800 ;
        RECT 676.800 486.900 678.900 489.000 ;
        RECT 671.400 479.100 673.500 481.200 ;
        RECT 677.100 479.700 678.300 486.900 ;
        RECT 679.800 483.600 681.300 501.300 ;
        RECT 679.800 481.500 681.900 483.600 ;
        RECT 670.950 475.950 673.050 478.050 ;
        RECT 676.800 477.600 678.900 479.700 ;
        RECT 679.800 476.700 681.300 481.500 ;
        RECT 683.100 479.700 684.300 501.300 ;
        RECT 667.950 469.950 670.050 472.050 ;
        RECT 671.400 463.050 672.450 475.950 ;
        RECT 679.200 474.600 681.300 476.700 ;
        RECT 682.200 474.600 684.300 479.700 ;
        RECT 685.200 501.300 687.300 503.400 ;
        RECT 685.200 483.600 686.700 501.300 ;
        RECT 695.400 492.450 696.600 492.600 ;
        RECT 689.400 491.400 696.600 492.450 ;
        RECT 689.400 487.050 690.450 491.400 ;
        RECT 695.400 490.350 696.600 491.400 ;
        RECT 694.800 487.950 696.900 490.050 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 685.200 481.500 687.300 483.600 ;
        RECT 685.200 476.700 686.700 481.500 ;
        RECT 685.200 474.600 687.300 476.700 ;
        RECT 685.950 469.950 688.050 472.050 ;
        RECT 682.950 466.950 685.050 469.050 ;
        RECT 670.950 460.950 673.050 463.050 ;
        RECT 652.950 449.100 655.050 451.200 ;
        RECT 658.950 450.000 661.050 454.050 ;
        RECT 653.400 439.050 654.450 449.100 ;
        RECT 659.400 448.350 660.600 450.000 ;
        RECT 664.950 449.100 667.050 451.200 ;
        RECT 683.400 451.050 684.450 466.950 ;
        RECT 665.400 448.350 666.600 449.100 ;
        RECT 682.950 448.950 685.050 451.050 ;
        RECT 686.400 450.600 687.450 469.950 ;
        RECT 698.400 456.450 699.450 517.800 ;
        RECT 704.400 492.600 705.450 521.400 ;
        RECT 706.950 520.800 709.050 522.900 ;
        RECT 713.400 521.400 714.600 523.650 ;
        RECT 719.400 521.400 720.600 523.650 ;
        RECT 713.400 517.050 714.450 521.400 ;
        RECT 712.950 514.950 715.050 517.050 ;
        RECT 709.950 511.950 712.050 514.050 ;
        RECT 704.400 492.450 705.600 492.600 ;
        RECT 704.400 491.400 708.450 492.450 ;
        RECT 704.400 490.350 705.600 491.400 ;
        RECT 703.800 487.950 705.900 490.050 ;
        RECT 707.400 483.450 708.450 491.400 ;
        RECT 704.400 482.400 708.450 483.450 ;
        RECT 698.400 455.400 702.450 456.450 ;
        RECT 686.400 448.350 687.600 450.600 ;
        RECT 691.950 450.000 694.050 454.050 ;
        RECT 697.950 451.950 700.050 454.050 ;
        RECT 692.400 448.350 693.600 450.000 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 662.400 444.900 663.600 445.650 ;
        RECT 661.950 442.800 664.050 444.900 ;
        RECT 668.400 443.400 669.600 445.650 ;
        RECT 652.950 436.950 655.050 439.050 ;
        RECT 664.950 436.950 667.050 439.050 ;
        RECT 649.950 433.950 652.050 436.050 ;
        RECT 631.950 430.950 634.050 433.050 ;
        RECT 640.950 427.950 643.050 430.050 ;
        RECT 625.950 421.950 628.050 424.050 ;
        RECT 628.950 420.450 633.000 421.050 ;
        RECT 628.950 418.950 633.450 420.450 ;
        RECT 625.950 416.100 628.050 418.200 ;
        RECT 632.400 417.600 633.450 418.950 ;
        RECT 626.400 415.350 627.600 416.100 ;
        RECT 632.400 415.350 633.600 417.600 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 623.400 410.400 624.600 412.650 ;
        RECT 629.400 411.900 630.600 412.650 ;
        RECT 623.400 385.050 624.450 410.400 ;
        RECT 628.950 409.800 631.050 411.900 ;
        RECT 638.400 400.050 639.450 412.950 ;
        RECT 637.950 397.950 640.050 400.050 ;
        RECT 622.950 382.950 625.050 385.050 ;
        RECT 616.950 373.950 619.050 376.050 ;
        RECT 617.400 366.900 618.450 373.950 ;
        RECT 625.950 371.100 628.050 373.200 ;
        RECT 626.400 370.350 627.600 371.100 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 623.400 366.900 624.600 367.650 ;
        RECT 629.400 366.900 630.600 367.650 ;
        RECT 598.950 364.800 601.050 366.900 ;
        RECT 604.950 364.800 607.050 366.900 ;
        RECT 610.950 364.800 613.050 366.900 ;
        RECT 616.950 364.800 619.050 366.900 ;
        RECT 622.950 364.800 625.050 366.900 ;
        RECT 628.950 364.800 631.050 366.900 ;
        RECT 592.950 361.950 595.050 364.050 ;
        RECT 599.400 361.050 600.450 364.800 ;
        RECT 598.950 358.950 601.050 361.050 ;
        RECT 589.950 343.950 592.050 346.050 ;
        RECT 601.950 343.950 604.050 346.050 ;
        RECT 587.400 341.400 591.450 342.450 ;
        RECT 580.950 337.950 583.050 340.050 ;
        RECT 590.400 339.600 591.450 341.400 ;
        RECT 581.400 333.900 582.450 337.950 ;
        RECT 590.400 337.350 591.600 339.600 ;
        RECT 595.950 338.100 598.050 340.200 ;
        RECT 596.400 337.350 597.600 338.100 ;
        RECT 602.400 337.050 603.450 343.950 ;
        RECT 605.400 340.200 606.450 364.800 ;
        RECT 641.400 364.050 642.450 427.950 ;
        RECT 665.400 427.050 666.450 436.950 ;
        RECT 668.400 433.050 669.450 443.400 ;
        RECT 667.950 430.950 670.050 433.050 ;
        RECT 664.950 424.950 667.050 427.050 ;
        RECT 643.950 415.950 646.050 418.050 ;
        RECT 652.950 417.000 655.050 421.050 ;
        RECT 644.400 403.050 645.450 415.950 ;
        RECT 653.400 415.350 654.600 417.000 ;
        RECT 649.950 412.950 652.050 415.050 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 650.400 411.900 651.600 412.650 ;
        RECT 649.950 409.800 652.050 411.900 ;
        RECT 665.400 411.450 666.450 424.950 ;
        RECT 680.400 421.050 681.450 445.950 ;
        RECT 689.400 443.400 690.600 445.650 ;
        RECT 698.400 444.900 699.450 451.950 ;
        RECT 673.950 417.000 676.050 421.050 ;
        RECT 679.950 418.950 682.050 421.050 ;
        RECT 685.950 418.950 688.050 421.050 ;
        RECT 680.400 417.600 681.450 418.950 ;
        RECT 674.400 415.350 675.600 417.000 ;
        RECT 680.400 415.350 681.600 417.600 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 671.400 411.450 672.600 412.650 ;
        RECT 677.400 411.900 678.600 412.650 ;
        RECT 665.400 410.400 672.600 411.450 ;
        RECT 643.950 400.950 646.050 403.050 ;
        RECT 655.950 397.950 658.050 400.050 ;
        RECT 643.950 388.950 646.050 391.050 ;
        RECT 644.400 364.050 645.450 388.950 ;
        RECT 646.950 371.100 649.050 373.200 ;
        RECT 656.400 372.600 657.450 397.950 ;
        RECT 661.950 385.950 664.050 388.050 ;
        RECT 662.400 379.050 663.450 385.950 ;
        RECT 661.950 376.950 664.050 379.050 ;
        RECT 658.950 373.950 661.050 376.050 ;
        RECT 664.950 373.950 667.050 376.050 ;
        RECT 647.400 370.350 648.600 371.100 ;
        RECT 656.400 370.350 657.600 372.600 ;
        RECT 647.100 367.950 649.200 370.050 ;
        RECT 652.500 367.950 654.600 370.050 ;
        RECT 655.800 367.950 657.900 370.050 ;
        RECT 653.400 365.400 654.600 367.650 ;
        RECT 659.400 366.900 660.450 373.950 ;
        RECT 628.950 361.650 631.050 363.750 ;
        RECT 640.950 361.950 643.050 364.050 ;
        RECT 643.950 361.950 646.050 364.050 ;
        RECT 607.950 358.950 610.050 361.050 ;
        RECT 604.950 338.100 607.050 340.200 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 587.400 333.900 588.600 334.650 ;
        RECT 580.950 331.800 583.050 333.900 ;
        RECT 586.950 331.800 589.050 333.900 ;
        RECT 593.400 332.400 594.600 334.650 ;
        RECT 577.950 328.950 580.050 331.050 ;
        RECT 593.400 319.050 594.450 332.400 ;
        RECT 595.950 319.950 598.050 322.050 ;
        RECT 592.950 316.950 595.050 319.050 ;
        RECT 583.950 304.950 586.050 307.050 ;
        RECT 580.800 292.950 582.900 295.050 ;
        RECT 581.400 291.900 582.600 292.650 ;
        RECT 580.950 289.800 583.050 291.900 ;
        RECT 577.950 274.950 580.050 277.050 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 556.950 262.950 559.050 265.050 ;
        RECT 568.950 262.950 571.050 265.050 ;
        RECT 548.400 259.350 549.600 261.600 ;
        RECT 515.400 256.350 516.600 258.600 ;
        RECT 517.950 256.800 520.050 258.900 ;
        RECT 524.400 258.450 525.600 258.600 ;
        RECT 524.400 258.000 528.450 258.450 ;
        RECT 524.400 257.400 529.050 258.000 ;
        RECT 514.800 253.950 516.900 256.050 ;
        RECT 511.950 244.950 514.050 247.050 ;
        RECT 512.400 220.050 513.450 244.950 ;
        RECT 518.400 244.050 519.450 256.800 ;
        RECT 524.400 256.350 525.600 257.400 ;
        RECT 523.800 253.950 525.900 256.050 ;
        RECT 526.950 253.950 529.050 257.400 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 545.400 255.900 546.600 256.650 ;
        RECT 551.400 255.900 552.600 256.650 ;
        RECT 557.400 255.900 558.450 262.950 ;
        RECT 569.400 261.600 570.450 262.950 ;
        RECT 569.400 259.350 570.600 261.600 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 544.950 253.800 547.050 255.900 ;
        RECT 550.950 253.800 553.050 255.900 ;
        RECT 556.950 253.800 559.050 255.900 ;
        RECT 572.400 254.400 573.600 256.650 ;
        RECT 551.400 247.050 552.450 253.800 ;
        RECT 550.950 244.950 553.050 247.050 ;
        RECT 517.950 241.950 520.050 244.050 ;
        RECT 572.400 235.050 573.450 254.400 ;
        RECT 571.950 232.950 574.050 235.050 ;
        RECT 514.950 231.450 517.050 232.050 ;
        RECT 520.950 231.450 523.050 232.050 ;
        RECT 514.950 230.400 523.050 231.450 ;
        RECT 514.950 229.950 517.050 230.400 ;
        RECT 520.950 229.950 523.050 230.400 ;
        RECT 517.950 226.950 520.050 229.050 ;
        RECT 536.400 228.300 539.400 230.400 ;
        RECT 540.300 228.300 542.400 230.400 ;
        RECT 559.200 228.300 561.300 230.400 ;
        RECT 518.400 220.200 519.450 226.950 ;
        RECT 511.950 217.950 514.050 220.050 ;
        RECT 517.950 216.000 520.050 220.200 ;
        RECT 523.950 218.100 526.050 220.200 ;
        RECT 524.400 217.350 525.600 218.100 ;
        RECT 518.400 214.350 519.600 216.000 ;
        RECT 523.800 214.950 525.900 217.050 ;
        RECT 529.800 214.950 531.900 217.050 ;
        RECT 512.400 211.950 514.500 214.050 ;
        RECT 517.800 211.950 519.900 214.050 ;
        RECT 512.400 209.400 513.600 211.650 ;
        RECT 536.400 209.400 537.900 228.300 ;
        RECT 540.300 222.300 541.500 228.300 ;
        RECT 539.400 220.200 541.500 222.300 ;
        RECT 508.950 205.950 511.050 208.050 ;
        RECT 512.400 184.050 513.450 209.400 ;
        RECT 536.400 207.300 538.500 209.400 ;
        RECT 537.300 203.700 538.500 207.300 ;
        RECT 540.300 203.700 541.500 220.200 ;
        RECT 542.700 225.300 544.800 227.400 ;
        RECT 542.700 203.700 543.900 225.300 ;
        RECT 551.400 223.800 553.500 225.900 ;
        RECT 556.800 225.300 558.900 227.400 ;
        RECT 551.400 217.200 552.300 223.800 ;
        RECT 557.100 218.100 558.300 225.300 ;
        RECT 559.800 223.500 561.300 228.300 ;
        RECT 562.200 225.300 564.300 230.400 ;
        RECT 559.800 221.400 561.900 223.500 ;
        RECT 551.400 215.100 553.500 217.200 ;
        RECT 556.800 216.000 558.900 218.100 ;
        RECT 547.950 212.100 550.050 214.200 ;
        RECT 548.400 211.350 549.600 212.100 ;
        RECT 547.800 208.950 549.900 211.050 ;
        RECT 551.400 204.600 552.300 215.100 ;
        RECT 554.100 208.500 556.200 210.600 ;
        RECT 536.700 201.600 538.800 203.700 ;
        RECT 539.700 201.600 541.800 203.700 ;
        RECT 542.700 201.600 544.800 203.700 ;
        RECT 550.800 202.500 552.900 204.600 ;
        RECT 557.100 203.700 558.300 216.000 ;
        RECT 559.800 203.700 561.300 221.400 ;
        RECT 563.100 203.700 564.300 225.300 ;
        RECT 556.200 201.600 558.300 203.700 ;
        RECT 559.200 201.600 561.300 203.700 ;
        RECT 562.200 201.600 564.300 203.700 ;
        RECT 565.200 228.300 567.300 230.400 ;
        RECT 565.200 223.500 566.700 228.300 ;
        RECT 568.950 226.950 571.050 229.050 ;
        RECT 565.200 221.400 567.300 223.500 ;
        RECT 565.200 203.700 566.700 221.400 ;
        RECT 565.200 201.600 567.300 203.700 ;
        RECT 526.950 196.950 529.050 199.050 ;
        RECT 527.400 193.050 528.450 196.950 ;
        RECT 526.950 190.950 529.050 193.050 ;
        RECT 569.400 184.050 570.450 226.950 ;
        RECT 574.800 214.950 576.900 217.050 ;
        RECT 575.400 213.450 576.600 214.650 ;
        RECT 578.400 213.450 579.450 274.950 ;
        RECT 580.950 265.950 583.050 268.050 ;
        RECT 581.400 235.050 582.450 265.950 ;
        RECT 580.950 232.950 583.050 235.050 ;
        RECT 584.400 229.050 585.450 304.950 ;
        RECT 586.950 298.950 589.050 301.050 ;
        RECT 587.400 283.050 588.450 298.950 ;
        RECT 586.950 280.950 589.050 283.050 ;
        RECT 593.400 274.050 594.450 316.950 ;
        RECT 596.400 288.900 597.450 319.950 ;
        RECT 602.400 310.050 603.450 334.950 ;
        RECT 608.400 333.900 609.450 358.950 ;
        RECT 616.950 346.950 619.050 349.050 ;
        RECT 617.400 339.600 618.450 346.950 ;
        RECT 617.400 337.350 618.600 339.600 ;
        RECT 622.950 338.100 625.050 340.200 ;
        RECT 623.400 337.350 624.600 338.100 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 607.950 331.800 610.050 333.900 ;
        RECT 614.400 333.000 615.600 334.650 ;
        RECT 620.400 333.900 621.600 334.650 ;
        RECT 613.950 328.950 616.050 333.000 ;
        RECT 619.950 331.800 622.050 333.900 ;
        RECT 629.400 325.050 630.450 361.650 ;
        RECT 653.400 361.050 654.450 365.400 ;
        RECT 658.950 364.800 661.050 366.900 ;
        RECT 661.950 361.950 664.050 364.050 ;
        RECT 652.950 358.950 655.050 361.050 ;
        RECT 658.950 358.950 661.050 361.050 ;
        RECT 631.950 352.950 634.050 355.050 ;
        RECT 649.950 352.950 652.050 355.050 ;
        RECT 632.400 328.050 633.450 352.950 ;
        RECT 634.950 346.950 637.050 349.050 ;
        RECT 635.400 333.900 636.450 346.950 ;
        RECT 637.950 343.950 640.050 346.050 ;
        RECT 650.400 345.450 651.450 352.950 ;
        RECT 634.950 331.800 637.050 333.900 ;
        RECT 631.950 325.950 634.050 328.050 ;
        RECT 619.950 322.950 622.050 325.050 ;
        RECT 628.950 322.950 631.050 325.050 ;
        RECT 613.950 316.950 616.050 319.050 ;
        RECT 601.950 307.950 604.050 310.050 ;
        RECT 607.950 307.950 610.050 310.050 ;
        RECT 602.400 297.450 603.450 307.950 ;
        RECT 608.400 298.050 609.450 307.950 ;
        RECT 602.400 296.400 606.450 297.450 ;
        RECT 605.400 294.600 606.450 296.400 ;
        RECT 607.950 295.950 610.050 298.050 ;
        RECT 605.400 292.350 606.600 294.600 ;
        RECT 610.950 294.450 613.050 295.200 ;
        RECT 614.400 294.450 615.450 316.950 ;
        RECT 610.950 293.400 615.450 294.450 ;
        RECT 610.950 293.100 613.050 293.400 ;
        RECT 611.400 292.350 612.600 293.100 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 610.950 289.950 613.050 292.050 ;
        RECT 602.400 288.900 603.600 289.650 ;
        RECT 608.400 288.900 609.600 289.650 ;
        RECT 595.950 286.800 598.050 288.900 ;
        RECT 601.950 286.800 604.050 288.900 ;
        RECT 607.950 286.800 610.050 288.900 ;
        RECT 592.950 271.950 595.050 274.050 ;
        RECT 604.950 271.950 607.050 274.050 ;
        RECT 589.950 260.100 592.050 262.200 ;
        RECT 590.400 259.350 591.600 260.100 ;
        RECT 598.950 259.950 601.050 262.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 593.400 254.400 594.600 256.650 ;
        RECT 593.400 250.050 594.450 254.400 ;
        RECT 592.950 247.950 595.050 250.050 ;
        RECT 599.400 244.050 600.450 259.950 ;
        RECT 598.950 241.950 601.050 244.050 ;
        RECT 598.950 232.950 601.050 235.050 ;
        RECT 583.950 226.950 586.050 229.050 ;
        RECT 586.950 223.950 589.050 226.050 ;
        RECT 583.800 214.950 585.900 217.050 ;
        RECT 575.400 212.400 579.450 213.450 ;
        RECT 584.400 213.450 585.600 214.650 ;
        RECT 587.400 213.450 588.450 223.950 ;
        RECT 589.950 214.950 592.050 217.050 ;
        RECT 584.400 212.400 588.450 213.450 ;
        RECT 574.950 205.950 577.050 208.050 ;
        RECT 505.950 181.950 508.050 184.050 ;
        RECT 511.950 181.950 514.050 184.050 ;
        RECT 568.950 181.950 571.050 184.050 ;
        RECT 502.200 169.500 504.300 171.600 ;
        RECT 502.200 164.700 503.700 169.500 ;
        RECT 502.200 162.600 504.300 164.700 ;
        RECT 493.950 145.950 496.050 148.050 ;
        RECT 494.400 132.450 495.450 145.950 ;
        RECT 506.400 145.050 507.450 181.950 ;
        RECT 512.400 180.450 513.600 180.600 ;
        RECT 521.400 180.450 522.600 180.600 ;
        RECT 512.400 180.000 516.450 180.450 ;
        RECT 512.400 179.400 517.050 180.000 ;
        RECT 512.400 178.350 513.600 179.400 ;
        RECT 511.800 175.950 513.900 178.050 ;
        RECT 514.950 175.950 517.050 179.400 ;
        RECT 521.400 179.400 525.450 180.450 ;
        RECT 521.400 178.350 522.600 179.400 ;
        RECT 520.800 175.950 522.900 178.050 ;
        RECT 515.400 166.050 516.450 175.950 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 517.950 154.950 520.050 157.050 ;
        RECT 514.950 148.950 517.050 151.050 ;
        RECT 500.100 142.500 502.200 144.600 ;
        RECT 505.950 142.950 508.050 145.050 ;
        RECT 497.100 133.950 499.200 136.050 ;
        RECT 500.100 135.900 501.000 142.500 ;
        RECT 509.100 142.200 511.200 144.300 ;
        RECT 503.400 139.350 504.600 141.600 ;
        RECT 502.800 136.950 504.900 139.050 ;
        RECT 507.000 135.900 509.100 136.200 ;
        RECT 500.100 135.000 509.100 135.900 ;
        RECT 497.400 132.450 498.600 133.650 ;
        RECT 494.400 131.400 498.600 132.450 ;
        RECT 500.100 129.900 501.000 135.000 ;
        RECT 507.000 134.100 509.100 135.000 ;
        RECT 501.900 133.200 504.000 134.100 ;
        RECT 501.900 132.000 509.100 133.200 ;
        RECT 507.000 131.100 509.100 132.000 ;
        RECT 499.500 127.800 501.600 129.900 ;
        RECT 502.800 128.100 504.900 130.200 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 503.400 126.450 504.600 127.800 ;
        RECT 505.950 126.450 508.050 130.050 ;
        RECT 510.000 129.600 510.900 142.200 ;
        RECT 515.400 142.050 516.450 148.950 ;
        RECT 514.950 139.950 517.050 142.050 ;
        RECT 511.950 138.450 514.050 139.200 ;
        RECT 511.950 137.400 516.450 138.450 ;
        RECT 511.950 137.100 514.050 137.400 ;
        RECT 512.400 136.350 513.600 137.100 ;
        RECT 511.800 133.950 513.900 136.050 ;
        RECT 509.400 127.500 511.500 129.600 ;
        RECT 503.400 126.000 508.050 126.450 ;
        RECT 503.400 125.400 507.450 126.000 ;
        RECT 491.400 105.600 492.450 124.950 ;
        RECT 515.400 124.050 516.450 137.400 ;
        RECT 518.400 130.050 519.450 154.950 ;
        RECT 520.950 139.950 523.050 142.050 ;
        RECT 521.400 132.900 522.450 139.950 ;
        RECT 520.950 130.800 523.050 132.900 ;
        RECT 517.950 127.950 520.050 130.050 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 508.950 118.950 511.050 121.050 ;
        RECT 509.400 105.600 510.450 118.950 ;
        RECT 514.950 109.950 517.050 112.050 ;
        RECT 515.400 105.600 516.450 109.950 ;
        RECT 479.400 103.350 480.600 105.600 ;
        RECT 485.400 103.350 486.600 105.600 ;
        RECT 491.400 103.350 492.600 105.600 ;
        RECT 509.400 103.350 510.600 105.600 ;
        RECT 515.400 103.350 516.600 105.600 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 517.950 100.950 520.050 103.050 ;
        RECT 424.950 94.950 427.050 97.050 ;
        RECT 425.400 88.050 426.450 94.950 ;
        RECT 424.950 85.950 427.050 88.050 ;
        RECT 439.950 73.950 442.050 76.050 ;
        RECT 424.950 64.950 427.050 67.050 ;
        RECT 403.950 61.950 406.050 64.050 ;
        RECT 380.400 52.050 381.450 59.100 ;
        RECT 386.400 58.350 387.600 60.600 ;
        RECT 391.950 59.100 394.050 61.200 ;
        RECT 400.950 59.100 403.050 61.200 ;
        RECT 392.400 58.350 393.600 59.100 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 389.400 54.900 390.600 55.650 ;
        RECT 388.950 52.800 391.050 54.900 ;
        RECT 379.950 49.950 382.050 52.050 ;
        RECT 397.950 46.950 400.050 49.050 ;
        RECT 391.950 34.950 394.050 37.050 ;
        RECT 367.950 28.950 370.050 31.050 ;
        RECT 376.950 28.950 379.050 31.050 ;
        RECT 368.400 24.600 369.450 28.950 ;
        RECT 368.400 22.350 369.600 24.600 ;
        RECT 370.950 23.100 373.050 25.200 ;
        RECT 376.950 23.100 379.050 25.200 ;
        RECT 367.800 19.950 369.900 22.050 ;
        RECT 361.950 16.800 364.050 18.900 ;
        RECT 358.200 13.500 360.300 15.600 ;
        RECT 358.200 8.700 359.700 13.500 ;
        RECT 371.400 13.050 372.450 23.100 ;
        RECT 377.400 22.350 378.600 23.100 ;
        RECT 376.800 19.950 378.900 22.050 ;
        RECT 392.400 21.900 393.450 34.950 ;
        RECT 398.400 27.600 399.450 46.950 ;
        RECT 401.400 40.050 402.450 59.100 ;
        RECT 404.400 55.050 405.450 61.950 ;
        RECT 409.950 60.000 412.050 64.050 ;
        RECT 418.950 61.950 421.050 64.050 ;
        RECT 410.400 58.350 411.600 60.000 ;
        RECT 415.950 59.100 418.050 61.200 ;
        RECT 416.400 58.350 417.600 59.100 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 413.400 54.900 414.600 55.650 ;
        RECT 412.950 52.800 415.050 54.900 ;
        RECT 421.950 46.950 424.050 49.050 ;
        RECT 403.950 40.950 406.050 43.050 ;
        RECT 400.950 37.950 403.050 40.050 ;
        RECT 404.400 37.050 405.450 40.950 ;
        RECT 403.950 34.950 406.050 37.050 ;
        RECT 398.400 25.350 399.600 27.600 ;
        RECT 403.950 26.100 406.050 28.200 ;
        RECT 404.400 25.350 405.600 26.100 ;
        RECT 418.950 25.950 421.050 28.050 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 401.400 21.900 402.600 22.650 ;
        RECT 407.400 21.900 408.600 22.650 ;
        RECT 391.950 19.800 394.050 21.900 ;
        RECT 400.950 19.800 403.050 21.900 ;
        RECT 406.950 19.800 409.050 21.900 ;
        RECT 419.400 13.050 420.450 25.950 ;
        RECT 422.400 21.450 423.450 46.950 ;
        RECT 425.400 46.050 426.450 64.950 ;
        RECT 427.950 61.950 430.050 64.050 ;
        RECT 424.950 43.950 427.050 46.050 ;
        RECT 428.400 34.050 429.450 61.950 ;
        RECT 433.950 59.100 436.050 61.200 ;
        RECT 440.400 60.600 441.450 73.950 ;
        RECT 434.400 58.350 435.600 59.100 ;
        RECT 440.400 58.350 441.600 60.600 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 437.400 53.400 438.600 55.650 ;
        RECT 443.400 54.900 444.600 55.650 ;
        RECT 455.400 55.050 456.450 98.400 ;
        RECT 460.950 97.800 463.050 99.900 ;
        RECT 466.950 97.800 469.050 99.900 ;
        RECT 482.400 98.400 483.600 100.650 ;
        RECT 488.400 98.400 489.600 100.650 ;
        RECT 512.400 98.400 513.600 100.650 ;
        RECT 518.400 98.400 519.600 100.650 ;
        RECT 461.400 76.050 462.450 97.800 ;
        RECT 460.950 73.950 463.050 76.050 ;
        RECT 482.400 73.050 483.450 98.400 ;
        RECT 488.400 94.050 489.450 98.400 ;
        RECT 512.400 97.050 513.450 98.400 ;
        RECT 511.950 94.950 514.050 97.050 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 488.400 85.050 489.450 91.950 ;
        RECT 487.950 82.950 490.050 85.050 ;
        RECT 490.950 73.950 493.050 76.050 ;
        RECT 481.950 70.950 484.050 73.050 ;
        RECT 463.800 64.200 465.900 66.300 ;
        RECT 472.800 64.500 474.900 66.600 ;
        RECT 461.400 60.450 462.600 60.600 ;
        RECT 458.400 59.400 462.600 60.450 ;
        RECT 437.400 49.050 438.450 53.400 ;
        RECT 442.950 52.800 445.050 54.900 ;
        RECT 454.950 52.950 457.050 55.050 ;
        RECT 436.950 46.950 439.050 49.050 ;
        RECT 433.950 37.950 436.050 40.050 ;
        RECT 427.950 31.950 430.050 34.050 ;
        RECT 434.400 33.450 435.450 37.950 ;
        RECT 434.400 31.200 435.600 33.450 ;
        RECT 429.900 27.900 432.000 29.700 ;
        RECT 433.800 28.800 435.900 30.900 ;
        RECT 437.100 30.300 439.200 32.400 ;
        RECT 442.950 31.950 445.050 34.050 ;
        RECT 428.400 26.700 437.100 27.900 ;
        RECT 425.100 22.950 427.200 25.050 ;
        RECT 425.400 21.450 426.600 22.650 ;
        RECT 422.400 20.400 426.600 21.450 ;
        RECT 428.400 17.700 429.300 26.700 ;
        RECT 435.000 25.800 437.100 26.700 ;
        RECT 438.000 24.900 438.900 30.300 ;
        RECT 440.400 27.450 441.600 27.600 ;
        RECT 443.400 27.450 444.450 31.950 ;
        RECT 455.400 30.450 456.450 52.950 ;
        RECT 458.400 49.050 459.450 59.400 ;
        RECT 461.400 58.350 462.600 59.400 ;
        RECT 461.100 55.950 463.200 58.050 ;
        RECT 464.100 51.600 465.000 64.200 ;
        RECT 470.400 61.350 471.600 63.600 ;
        RECT 470.100 58.950 472.200 61.050 ;
        RECT 465.900 57.900 468.000 58.200 ;
        RECT 474.000 57.900 474.900 64.500 ;
        RECT 465.900 57.000 474.900 57.900 ;
        RECT 465.900 56.100 468.000 57.000 ;
        RECT 471.000 55.200 473.100 56.100 ;
        RECT 465.900 54.000 473.100 55.200 ;
        RECT 465.900 53.100 468.000 54.000 ;
        RECT 463.500 49.500 465.600 51.600 ;
        RECT 470.100 50.100 472.200 52.200 ;
        RECT 474.000 51.900 474.900 57.000 ;
        RECT 475.800 55.950 477.900 58.050 ;
        RECT 476.400 54.450 477.600 55.650 ;
        RECT 476.400 53.400 480.450 54.450 ;
        RECT 473.400 49.800 475.500 51.900 ;
        RECT 470.400 49.050 471.600 49.800 ;
        RECT 457.950 46.950 460.050 49.050 ;
        RECT 469.950 46.950 472.050 49.050 ;
        RECT 479.400 40.050 480.450 53.400 ;
        RECT 472.950 37.950 475.050 40.050 ;
        RECT 478.950 37.950 481.050 40.050 ;
        RECT 455.400 29.400 459.450 30.450 ;
        RECT 440.400 26.400 444.450 27.450 ;
        RECT 440.400 25.350 441.600 26.400 ;
        RECT 432.000 23.700 438.900 24.900 ;
        RECT 432.000 21.300 432.900 23.700 ;
        RECT 430.800 19.200 432.900 21.300 ;
        RECT 433.800 19.950 435.900 22.050 ;
        RECT 427.500 15.600 429.600 17.700 ;
        RECT 434.400 17.400 435.600 19.650 ;
        RECT 437.700 16.500 438.900 23.700 ;
        RECT 439.800 22.950 441.900 25.050 ;
        RECT 443.400 21.900 444.450 26.400 ;
        RECT 458.400 27.600 459.450 29.400 ;
        RECT 458.400 25.350 459.600 27.600 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 442.950 19.800 445.050 21.900 ;
        RECT 461.400 20.400 462.600 22.650 ;
        RECT 473.400 21.900 474.450 37.950 ;
        RECT 491.400 31.050 492.450 73.950 ;
        RECT 505.950 70.950 508.050 73.050 ;
        RECT 493.950 64.950 496.050 67.050 ;
        RECT 494.400 60.600 495.450 64.950 ;
        RECT 494.400 58.350 495.600 60.600 ;
        RECT 503.400 60.450 504.600 60.600 ;
        RECT 506.400 60.450 507.450 70.950 ;
        RECT 503.400 59.400 507.450 60.450 ;
        RECT 503.400 58.350 504.600 59.400 ;
        RECT 494.100 55.950 496.200 58.050 ;
        RECT 499.500 55.950 501.600 58.050 ;
        RECT 502.800 55.950 504.900 58.050 ;
        RECT 500.400 54.900 501.600 55.650 ;
        RECT 499.950 52.800 502.050 54.900 ;
        RECT 506.400 49.050 507.450 59.400 ;
        RECT 505.950 46.950 508.050 49.050 ;
        RECT 512.400 46.050 513.450 94.950 ;
        RECT 518.400 91.050 519.450 98.400 ;
        RECT 517.950 88.950 520.050 91.050 ;
        RECT 524.400 79.050 525.450 179.400 ;
        RECT 545.100 178.950 547.200 181.050 ;
        RECT 563.100 178.950 565.200 181.050 ;
        RECT 545.400 177.900 546.600 178.650 ;
        RECT 544.950 175.800 547.050 177.900 ;
        RECT 569.400 166.050 570.450 181.950 ;
        RECT 568.950 163.950 571.050 166.050 ;
        RECT 538.950 160.950 541.050 163.050 ;
        RECT 532.950 137.100 535.050 139.200 ;
        RECT 539.400 138.600 540.450 160.950 ;
        RECT 553.950 148.950 556.050 151.050 ;
        RECT 533.400 136.350 534.600 137.100 ;
        RECT 539.400 136.350 540.600 138.600 ;
        RECT 550.950 137.100 553.050 139.200 ;
        RECT 554.400 138.450 555.450 148.950 ;
        RECT 559.500 141.300 561.600 143.400 ;
        RECT 569.100 142.500 571.200 144.600 ;
        RECT 557.400 138.450 558.600 138.600 ;
        RECT 554.400 137.400 558.600 138.450 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 530.400 132.900 531.600 133.650 ;
        RECT 529.950 130.800 532.050 132.900 ;
        RECT 536.400 131.400 537.600 133.650 ;
        RECT 536.400 124.050 537.450 131.400 ;
        RECT 535.950 121.950 538.050 124.050 ;
        RECT 538.950 109.950 541.050 112.050 ;
        RECT 539.400 105.600 540.450 109.950 ;
        RECT 539.400 103.350 540.600 105.600 ;
        RECT 544.950 105.000 547.050 109.050 ;
        RECT 545.400 103.350 546.600 105.000 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 541.950 100.950 544.050 103.050 ;
        RECT 544.950 100.950 547.050 103.050 ;
        RECT 536.400 99.000 537.600 100.650 ;
        RECT 542.400 99.900 543.600 100.650 ;
        RECT 535.950 94.950 538.050 99.000 ;
        RECT 541.950 97.800 544.050 99.900 ;
        RECT 551.400 99.450 552.450 137.100 ;
        RECT 557.400 136.350 558.600 137.400 ;
        RECT 557.100 133.950 559.200 136.050 ;
        RECT 560.400 132.300 561.300 141.300 ;
        RECT 562.800 137.700 564.900 139.800 ;
        RECT 566.400 139.350 567.600 141.600 ;
        RECT 564.000 135.300 564.900 137.700 ;
        RECT 565.800 136.950 567.900 139.050 ;
        RECT 569.700 135.300 570.900 142.500 ;
        RECT 564.000 134.100 570.900 135.300 ;
        RECT 567.000 132.300 569.100 133.200 ;
        RECT 560.400 131.100 569.100 132.300 ;
        RECT 561.900 129.300 564.000 131.100 ;
        RECT 565.800 128.100 567.900 130.200 ;
        RECT 570.000 128.700 570.900 134.100 ;
        RECT 571.800 133.950 573.900 136.050 ;
        RECT 572.400 132.900 573.600 133.650 ;
        RECT 571.950 130.800 574.050 132.900 ;
        RECT 575.400 130.050 576.450 205.950 ;
        RECT 583.950 199.950 586.050 202.050 ;
        RECT 577.950 187.950 580.050 190.050 ;
        RECT 578.400 157.050 579.450 187.950 ;
        RECT 584.400 183.600 585.450 199.950 ;
        RECT 590.400 183.600 591.450 214.950 ;
        RECT 599.400 210.900 600.450 232.950 ;
        RECT 605.400 229.050 606.450 271.950 ;
        RECT 620.400 271.050 621.450 322.950 ;
        RECT 628.950 313.950 631.050 316.050 ;
        RECT 629.400 307.050 630.450 313.950 ;
        RECT 628.950 304.950 631.050 307.050 ;
        RECT 638.400 298.050 639.450 343.950 ;
        RECT 643.500 341.400 645.600 343.500 ;
        RECT 650.400 343.200 651.600 345.450 ;
        RECT 641.100 334.950 643.200 337.050 ;
        RECT 641.400 333.900 642.600 334.650 ;
        RECT 640.950 331.800 643.050 333.900 ;
        RECT 644.100 328.800 645.000 341.400 ;
        RECT 650.100 340.800 652.200 342.900 ;
        RECT 653.400 341.100 655.500 343.200 ;
        RECT 645.900 339.000 648.000 339.900 ;
        RECT 645.900 337.800 653.100 339.000 ;
        RECT 651.000 336.900 653.100 337.800 ;
        RECT 645.900 336.000 648.000 336.900 ;
        RECT 654.000 336.000 654.900 341.100 ;
        RECT 656.400 339.450 657.600 339.600 ;
        RECT 659.400 339.450 660.450 358.950 ;
        RECT 656.400 338.400 660.450 339.450 ;
        RECT 656.400 337.350 657.600 338.400 ;
        RECT 645.900 335.100 654.900 336.000 ;
        RECT 645.900 334.800 648.000 335.100 ;
        RECT 650.100 331.950 652.200 334.050 ;
        RECT 646.950 328.950 649.050 331.050 ;
        RECT 650.400 329.400 651.600 331.650 ;
        RECT 643.800 326.700 645.900 328.800 ;
        RECT 643.950 319.950 646.050 322.050 ;
        RECT 637.950 295.950 640.050 298.050 ;
        RECT 622.950 293.100 625.050 295.200 ;
        RECT 628.950 293.100 631.050 295.200 ;
        RECT 634.950 293.100 637.050 295.200 ;
        RECT 623.400 289.050 624.450 293.100 ;
        RECT 629.400 292.350 630.600 293.100 ;
        RECT 635.400 292.350 636.600 293.100 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 622.950 286.950 625.050 289.050 ;
        RECT 632.400 287.400 633.600 289.650 ;
        RECT 638.400 288.900 639.600 289.650 ;
        RECT 632.400 283.050 633.450 287.400 ;
        RECT 637.950 286.800 640.050 288.900 ;
        RECT 631.950 280.950 634.050 283.050 ;
        RECT 644.400 274.050 645.450 319.950 ;
        RECT 647.400 310.050 648.450 328.950 ;
        RECT 654.000 328.500 654.900 335.100 ;
        RECT 655.800 334.950 657.900 337.050 ;
        RECT 658.950 334.950 661.050 337.050 ;
        RECT 652.800 326.400 654.900 328.500 ;
        RECT 646.950 307.950 649.050 310.050 ;
        RECT 646.950 295.950 649.050 298.050 ;
        RECT 647.400 288.900 648.450 295.950 ;
        RECT 649.950 293.100 652.050 295.200 ;
        RECT 659.400 294.600 660.450 334.950 ;
        RECT 662.400 304.050 663.450 361.950 ;
        RECT 661.950 301.950 664.050 304.050 ;
        RECT 665.400 295.200 666.450 373.950 ;
        RECT 668.400 367.050 669.450 410.400 ;
        RECT 676.950 409.800 679.050 411.900 ;
        RECT 677.400 379.050 678.450 409.800 ;
        RECT 682.950 397.950 685.050 400.050 ;
        RECT 683.400 391.050 684.450 397.950 ;
        RECT 682.950 388.950 685.050 391.050 ;
        RECT 676.950 376.950 679.050 379.050 ;
        RECT 682.950 376.950 685.050 379.050 ;
        RECT 673.950 375.450 678.000 376.050 ;
        RECT 673.950 373.950 678.450 375.450 ;
        RECT 677.400 372.600 678.450 373.950 ;
        RECT 683.400 373.050 684.450 376.950 ;
        RECT 686.400 373.050 687.450 418.950 ;
        RECT 689.400 393.450 690.450 443.400 ;
        RECT 697.950 442.800 700.050 444.900 ;
        RECT 701.400 427.050 702.450 455.400 ;
        RECT 704.400 444.450 705.450 482.400 ;
        RECT 710.400 453.450 711.450 511.950 ;
        RECT 719.400 508.050 720.450 521.400 ;
        RECT 721.950 508.950 724.050 511.050 ;
        RECT 718.950 505.950 721.050 508.050 ;
        RECT 715.950 502.950 718.050 505.050 ;
        RECT 712.950 457.950 715.050 460.050 ;
        RECT 707.400 453.000 711.450 453.450 ;
        RECT 706.950 452.400 711.450 453.000 ;
        RECT 706.950 448.950 709.050 452.400 ;
        RECT 713.400 450.600 714.450 457.950 ;
        RECT 716.400 454.050 717.450 502.950 ;
        RECT 718.950 469.950 721.050 472.050 ;
        RECT 719.400 457.050 720.450 469.950 ;
        RECT 722.400 460.050 723.450 508.950 ;
        RECT 725.400 469.050 726.450 562.950 ;
        RECT 727.950 547.950 730.050 550.050 ;
        RECT 728.400 529.200 729.450 547.950 ;
        RECT 734.400 538.050 735.450 592.800 ;
        RECT 743.400 576.450 744.450 604.950 ;
        RECT 740.400 575.400 744.450 576.450 ;
        RECT 736.950 572.100 739.050 574.200 ;
        RECT 737.400 562.050 738.450 572.100 ;
        RECT 740.400 567.900 741.450 575.400 ;
        RECT 746.400 573.450 747.450 649.800 ;
        RECT 749.400 622.050 750.450 661.950 ;
        RECT 751.950 655.950 754.050 658.050 ;
        RECT 752.400 652.050 753.450 655.950 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 754.950 650.100 757.050 655.050 ;
        RECT 761.400 651.600 762.450 661.950 ;
        RECT 764.400 658.050 765.450 730.950 ;
        RECT 772.950 728.100 775.050 730.200 ;
        RECT 779.400 729.600 780.450 781.950 ;
        RECT 788.400 762.600 789.450 793.950 ;
        RECT 794.400 793.050 795.450 800.400 ;
        RECT 796.950 795.450 799.050 796.050 ;
        RECT 800.400 795.450 801.450 812.400 ;
        RECT 802.950 806.100 805.050 808.200 ;
        RECT 811.950 806.100 814.050 808.200 ;
        RECT 818.400 807.600 819.450 812.400 ;
        RECT 826.950 811.950 829.050 814.050 ;
        RECT 803.400 799.050 804.450 806.100 ;
        RECT 812.400 805.350 813.600 806.100 ;
        RECT 818.400 805.350 819.600 807.600 ;
        RECT 823.950 805.950 826.050 811.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 809.400 801.000 810.600 802.650 ;
        RECT 815.400 801.900 816.600 802.650 ;
        RECT 802.950 796.950 805.050 799.050 ;
        RECT 808.950 796.950 811.050 801.000 ;
        RECT 814.950 796.950 817.050 801.900 ;
        RECT 820.950 796.950 823.050 799.050 ;
        RECT 796.950 794.400 801.450 795.450 ;
        RECT 796.950 793.950 799.050 794.400 ;
        RECT 793.950 790.950 796.050 793.050 ;
        RECT 797.400 784.050 798.450 793.950 ;
        RECT 799.950 790.800 802.050 792.900 ;
        RECT 796.950 781.950 799.050 784.050 ;
        RECT 796.950 775.950 799.050 778.050 ;
        RECT 788.400 760.350 789.600 762.600 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 781.950 754.950 784.050 757.050 ;
        RECT 785.400 755.400 786.600 757.650 ;
        RECT 791.400 756.900 792.600 757.650 ;
        RECT 797.400 756.900 798.450 775.950 ;
        RECT 782.400 751.050 783.450 754.950 ;
        RECT 781.950 748.950 784.050 751.050 ;
        RECT 785.400 745.050 786.450 755.400 ;
        RECT 790.950 754.800 793.050 756.900 ;
        RECT 796.950 754.800 799.050 756.900 ;
        RECT 800.400 748.050 801.450 790.800 ;
        RECT 805.950 787.950 808.050 790.050 ;
        RECT 806.400 784.050 807.450 787.950 ;
        RECT 821.400 784.050 822.450 796.950 ;
        RECT 805.950 781.950 808.050 784.050 ;
        RECT 820.950 781.950 823.050 784.050 ;
        RECT 805.950 775.950 808.050 778.050 ;
        RECT 806.400 766.050 807.450 775.950 ;
        RECT 814.950 766.950 817.050 769.050 ;
        RECT 805.950 763.950 808.050 766.050 ;
        RECT 808.950 761.100 811.050 763.200 ;
        RECT 815.400 762.600 816.450 766.950 ;
        RECT 809.400 760.350 810.600 761.100 ;
        RECT 815.400 760.350 816.600 762.600 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 812.400 755.400 813.600 757.650 ;
        RECT 821.400 757.050 822.450 781.950 ;
        RECT 823.950 778.950 826.050 781.050 ;
        RECT 808.950 751.950 811.050 754.050 ;
        RECT 799.950 745.950 802.050 748.050 ;
        RECT 784.950 744.450 787.050 745.050 ;
        RECT 784.950 743.400 789.450 744.450 ;
        RECT 784.950 742.950 787.050 743.400 ;
        RECT 773.400 727.350 774.600 728.100 ;
        RECT 779.400 727.350 780.600 729.600 ;
        RECT 784.950 728.100 787.050 730.200 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 766.950 721.950 769.050 724.050 ;
        RECT 770.400 722.400 771.600 724.650 ;
        RECT 776.400 723.900 777.600 724.650 ;
        RECT 767.400 679.050 768.450 721.950 ;
        RECT 770.400 718.050 771.450 722.400 ;
        RECT 775.950 718.950 778.050 723.900 ;
        RECT 769.950 715.950 772.050 718.050 ;
        RECT 775.950 715.800 778.050 717.900 ;
        RECT 781.950 715.950 784.050 718.050 ;
        RECT 776.400 712.050 777.450 715.800 ;
        RECT 785.400 715.050 786.450 728.100 ;
        RECT 784.950 712.950 787.050 715.050 ;
        RECT 769.950 709.950 772.050 712.050 ;
        RECT 775.950 709.950 778.050 712.050 ;
        RECT 781.950 709.950 784.050 712.050 ;
        RECT 770.400 700.050 771.450 709.950 ;
        RECT 788.400 700.050 789.450 743.400 ;
        RECT 790.950 736.950 793.050 739.050 ;
        RECT 791.400 721.050 792.450 736.950 ;
        RECT 793.950 727.950 796.050 730.050 ;
        RECT 800.400 729.600 801.450 745.950 ;
        RECT 800.400 727.350 801.600 729.600 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 797.400 724.050 798.600 724.650 ;
        RECT 793.950 722.400 798.600 724.050 ;
        RECT 803.400 723.000 804.600 724.650 ;
        RECT 793.950 721.950 798.000 722.400 ;
        RECT 790.950 718.950 793.050 721.050 ;
        RECT 802.950 718.950 805.050 723.000 ;
        RECT 805.950 721.800 808.050 723.900 ;
        RECT 793.950 715.950 796.050 718.050 ;
        RECT 790.950 709.950 793.050 712.050 ;
        RECT 794.400 703.050 795.450 715.950 ;
        RECT 802.950 715.800 805.050 717.900 ;
        RECT 803.400 712.050 804.450 715.800 ;
        RECT 802.950 709.950 805.050 712.050 ;
        RECT 799.950 703.950 802.050 706.050 ;
        RECT 793.950 700.950 796.050 703.050 ;
        RECT 769.950 697.950 772.050 700.050 ;
        RECT 787.950 697.950 790.050 700.050 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 763.950 655.950 766.050 658.050 ;
        RECT 755.400 649.350 756.600 650.100 ;
        RECT 761.400 649.350 762.600 651.600 ;
        RECT 767.400 651.450 768.600 651.600 ;
        RECT 770.400 651.450 771.450 697.950 ;
        RECT 781.950 694.950 784.050 697.050 ;
        RECT 775.950 683.100 778.050 685.200 ;
        RECT 782.400 684.600 783.450 694.950 ;
        RECT 800.400 688.050 801.450 703.950 ;
        RECT 806.400 700.050 807.450 721.800 ;
        RECT 809.400 714.450 810.450 751.950 ;
        RECT 812.400 730.200 813.450 755.400 ;
        RECT 817.950 754.950 820.050 757.050 ;
        RECT 820.950 754.950 823.050 757.050 ;
        RECT 818.400 735.450 819.450 754.950 ;
        RECT 824.400 748.050 825.450 778.950 ;
        RECT 827.400 763.200 828.450 811.950 ;
        RECT 830.400 796.050 831.450 817.950 ;
        RECT 836.400 814.050 837.450 833.400 ;
        RECT 841.950 832.950 844.050 835.050 ;
        RECT 844.950 832.950 847.050 835.050 ;
        RECT 844.950 828.450 847.050 829.050 ;
        RECT 848.400 828.450 849.450 892.950 ;
        RECT 860.400 885.600 861.450 895.950 ;
        RECT 860.400 883.350 861.600 885.600 ;
        RECT 877.950 884.100 880.050 886.200 ;
        RECT 886.950 884.100 889.050 886.200 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 859.950 880.950 862.050 883.050 ;
        RECT 862.950 880.950 865.050 883.050 ;
        RECT 857.400 878.400 858.600 880.650 ;
        RECT 863.400 878.400 864.600 880.650 ;
        RECT 857.400 874.050 858.450 878.400 ;
        RECT 856.950 871.950 859.050 874.050 ;
        RECT 863.400 868.050 864.450 878.400 ;
        RECT 878.400 868.050 879.450 884.100 ;
        RECT 887.400 883.350 888.600 884.100 ;
        RECT 881.100 880.950 883.200 883.050 ;
        RECT 886.500 880.950 888.600 883.050 ;
        RECT 889.800 880.950 891.900 883.050 ;
        RECT 881.400 878.400 882.600 880.650 ;
        RECT 890.400 878.400 891.600 880.650 ;
        RECT 881.400 874.050 882.450 878.400 ;
        RECT 890.400 877.050 891.450 878.400 ;
        RECT 893.400 877.050 894.450 898.950 ;
        RECT 899.400 885.450 900.450 911.400 ;
        RECT 905.400 907.050 906.450 917.100 ;
        RECT 904.950 904.950 907.050 907.050 ;
        RECT 907.950 892.950 910.050 895.050 ;
        RECT 908.400 889.050 909.450 892.950 ;
        RECT 907.950 886.950 910.050 889.050 ;
        RECT 911.400 886.200 912.450 917.100 ;
        RECT 917.400 916.350 918.600 918.000 ;
        RECT 922.950 917.100 925.050 919.200 ;
        RECT 934.950 917.100 937.050 919.200 ;
        RECT 940.950 917.100 943.050 919.200 ;
        RECT 946.950 917.100 949.050 919.200 ;
        RECT 923.400 916.350 924.600 917.100 ;
        RECT 916.950 913.950 919.050 916.050 ;
        RECT 919.950 913.950 922.050 916.050 ;
        RECT 922.950 913.950 925.050 916.050 ;
        RECT 925.950 913.950 928.050 916.050 ;
        RECT 920.400 911.400 921.600 913.650 ;
        RECT 926.400 912.900 927.600 913.650 ;
        RECT 935.400 913.050 936.450 917.100 ;
        RECT 941.400 916.350 942.600 917.100 ;
        RECT 947.400 916.350 948.600 917.100 ;
        RECT 940.950 913.950 943.050 916.050 ;
        RECT 943.950 913.950 946.050 916.050 ;
        RECT 946.950 913.950 949.050 916.050 ;
        RECT 920.400 901.050 921.450 911.400 ;
        RECT 925.950 910.800 928.050 912.900 ;
        RECT 934.950 912.450 937.050 913.050 ;
        RECT 932.400 911.400 937.050 912.450 ;
        RECT 922.950 901.950 925.050 904.050 ;
        RECT 919.950 898.950 922.050 901.050 ;
        RECT 899.400 884.400 903.450 885.450 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 890.400 875.400 895.050 877.050 ;
        RECT 891.000 874.950 895.050 875.400 ;
        RECT 895.950 874.950 898.050 877.050 ;
        RECT 880.950 871.950 883.050 874.050 ;
        RECT 862.950 865.950 865.050 868.050 ;
        RECT 877.950 865.950 880.050 868.050 ;
        RECT 865.950 859.950 868.050 862.050 ;
        RECT 856.950 839.100 859.050 841.200 ;
        RECT 857.400 838.350 858.600 839.100 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 850.950 834.450 853.050 835.050 ;
        RECT 854.400 834.450 855.600 835.650 ;
        RECT 850.950 833.400 855.600 834.450 ;
        RECT 860.400 833.400 861.600 835.650 ;
        RECT 866.400 835.050 867.450 859.950 ;
        RECT 868.950 853.950 871.050 856.050 ;
        RECT 869.400 835.050 870.450 853.950 ;
        RECT 881.400 850.050 882.450 871.950 ;
        RECT 886.950 865.950 889.050 868.050 ;
        RECT 880.950 847.950 883.050 850.050 ;
        RECT 871.950 838.950 874.050 841.050 ;
        RECT 880.950 839.100 883.050 841.200 ;
        RECT 887.400 840.600 888.450 865.950 ;
        RECT 892.950 850.950 895.050 853.050 ;
        RECT 896.400 852.450 897.450 874.950 ;
        RECT 899.400 874.050 900.450 880.950 ;
        RECT 902.400 877.050 903.450 884.400 ;
        RECT 910.950 884.100 913.050 886.200 ;
        RECT 916.950 884.100 919.050 886.200 ;
        RECT 911.400 883.350 912.600 884.100 ;
        RECT 917.400 883.350 918.600 884.100 ;
        RECT 907.950 880.950 910.050 883.050 ;
        RECT 910.950 880.950 913.050 883.050 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 908.400 879.000 909.600 880.650 ;
        RECT 914.400 879.000 915.600 880.650 ;
        RECT 901.950 874.950 904.050 877.050 ;
        RECT 907.950 874.950 910.050 879.000 ;
        RECT 913.950 874.950 916.050 879.000 ;
        RECT 919.950 877.950 922.050 880.050 ;
        RECT 898.950 871.950 901.050 874.050 ;
        RECT 920.400 865.050 921.450 877.950 ;
        RECT 919.950 862.950 922.050 865.050 ;
        RECT 913.950 856.950 916.050 859.050 ;
        RECT 914.400 853.050 915.450 856.950 ;
        RECT 923.400 856.050 924.450 901.950 ;
        RECT 928.950 895.950 931.050 898.050 ;
        RECT 925.950 883.950 928.050 886.050 ;
        RECT 922.950 853.950 925.050 856.050 ;
        RECT 896.400 851.400 900.450 852.450 ;
        RECT 850.950 832.950 853.050 833.400 ;
        RECT 844.950 827.400 849.450 828.450 ;
        RECT 844.950 826.950 847.050 827.400 ;
        RECT 845.400 820.050 846.450 826.950 ;
        RECT 851.400 826.050 852.450 832.950 ;
        RECT 853.950 829.950 856.050 832.050 ;
        RECT 850.950 823.950 853.050 826.050 ;
        RECT 847.950 820.950 850.050 823.050 ;
        RECT 844.950 817.950 847.050 820.050 ;
        RECT 844.950 814.800 847.050 816.900 ;
        RECT 835.950 811.950 838.050 814.050 ;
        RECT 838.950 807.000 841.050 811.050 ;
        RECT 845.400 807.600 846.450 814.800 ;
        RECT 848.400 808.050 849.450 820.950 ;
        RECT 850.950 817.950 853.050 820.050 ;
        RECT 839.400 805.350 840.600 807.000 ;
        RECT 845.400 805.350 846.600 807.600 ;
        RECT 847.950 805.950 850.050 808.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 841.950 802.950 844.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 836.400 801.000 837.600 802.650 ;
        RECT 835.950 796.950 838.050 801.000 ;
        RECT 842.400 800.400 843.600 802.650 ;
        RECT 829.950 793.950 832.050 796.050 ;
        RECT 842.400 784.050 843.450 800.400 ;
        RECT 851.400 799.050 852.450 817.950 ;
        RECT 847.950 793.950 850.050 799.050 ;
        RECT 850.950 796.950 853.050 799.050 ;
        RECT 850.950 787.950 853.050 790.050 ;
        RECT 847.950 784.950 850.050 787.050 ;
        RECT 841.950 781.950 844.050 784.050 ;
        RECT 842.400 772.050 843.450 781.950 ;
        RECT 848.400 778.050 849.450 784.950 ;
        RECT 847.950 775.950 850.050 778.050 ;
        RECT 841.950 769.950 844.050 772.050 ;
        RECT 826.950 761.100 829.050 763.200 ;
        RECT 835.950 761.100 838.050 763.200 ;
        RECT 841.950 761.100 844.050 763.200 ;
        RECT 827.400 757.050 828.450 761.100 ;
        RECT 836.400 760.350 837.600 761.100 ;
        RECT 842.400 760.350 843.600 761.100 ;
        RECT 847.950 760.950 850.050 763.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 826.950 754.950 829.050 757.050 ;
        RECT 833.400 756.900 834.600 757.650 ;
        RECT 839.400 756.900 840.600 757.650 ;
        RECT 832.950 754.800 835.050 756.900 ;
        RECT 838.950 754.800 841.050 756.900 ;
        RECT 844.950 754.950 847.050 757.050 ;
        RECT 823.950 745.950 826.050 748.050 ;
        RECT 829.950 742.950 832.050 745.050 ;
        RECT 841.950 742.950 844.050 745.050 ;
        RECT 830.400 739.050 831.450 742.950 ;
        RECT 829.950 736.950 832.050 739.050 ;
        RECT 815.400 734.400 819.450 735.450 ;
        RECT 811.950 728.100 814.050 730.200 ;
        RECT 815.400 723.450 816.450 734.400 ;
        RECT 823.950 728.100 826.050 730.200 ;
        RECT 829.950 728.100 832.050 730.200 ;
        RECT 824.400 727.350 825.600 728.100 ;
        RECT 830.400 727.350 831.600 728.100 ;
        RECT 838.950 727.950 841.050 730.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 815.400 722.400 819.450 723.450 ;
        RECT 814.950 718.950 817.050 721.050 ;
        RECT 811.950 714.450 814.050 715.050 ;
        RECT 809.400 713.400 814.050 714.450 ;
        RECT 811.950 712.950 814.050 713.400 ;
        RECT 805.950 697.950 808.050 700.050 ;
        RECT 805.950 694.800 808.050 696.900 ;
        RECT 802.950 688.950 805.050 691.050 ;
        RECT 784.950 685.950 787.050 688.050 ;
        RECT 799.950 685.950 802.050 688.050 ;
        RECT 776.400 682.350 777.600 683.100 ;
        RECT 782.400 682.350 783.600 684.600 ;
        RECT 787.950 683.100 790.050 685.200 ;
        RECT 788.400 682.350 789.600 683.100 ;
        RECT 796.950 682.950 799.050 685.050 ;
        RECT 803.400 684.450 804.450 688.950 ;
        RECT 800.400 683.400 804.450 684.450 ;
        RECT 806.400 684.600 807.450 694.800 ;
        RECT 812.400 685.050 813.450 712.950 ;
        RECT 815.400 703.050 816.450 718.950 ;
        RECT 814.950 700.950 817.050 703.050 ;
        RECT 814.950 694.950 817.050 697.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 787.950 679.950 790.050 682.050 ;
        RECT 779.400 678.900 780.600 679.650 ;
        RECT 778.950 676.800 781.050 678.900 ;
        RECT 785.400 678.000 786.600 679.650 ;
        RECT 784.950 673.950 787.050 678.000 ;
        RECT 793.950 676.950 796.050 679.050 ;
        RECT 790.950 673.950 793.050 676.050 ;
        RECT 791.400 661.050 792.450 673.950 ;
        RECT 794.400 673.050 795.450 676.950 ;
        RECT 793.950 670.950 796.050 673.050 ;
        RECT 797.400 664.050 798.450 682.950 ;
        RECT 800.400 675.450 801.450 683.400 ;
        RECT 806.400 682.350 807.600 684.600 ;
        RECT 811.950 682.950 814.050 685.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 809.400 678.000 810.600 679.650 ;
        RECT 802.950 675.450 805.050 676.050 ;
        RECT 808.950 675.450 811.050 678.000 ;
        RECT 811.950 676.950 814.050 679.050 ;
        RECT 800.400 674.400 805.050 675.450 ;
        RECT 806.400 675.000 811.050 675.450 ;
        RECT 802.950 673.950 805.050 674.400 ;
        RECT 805.950 674.400 811.050 675.000 ;
        RECT 796.950 661.950 799.050 664.050 ;
        RECT 775.950 658.950 778.050 661.050 ;
        RECT 790.950 658.950 793.050 661.050 ;
        RECT 767.400 650.400 774.450 651.450 ;
        RECT 767.400 649.350 768.600 650.400 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 751.950 643.950 754.050 646.050 ;
        RECT 758.400 644.400 759.600 646.650 ;
        RECT 764.400 644.400 765.600 646.650 ;
        RECT 748.950 619.950 751.050 622.050 ;
        RECT 752.400 613.050 753.450 643.950 ;
        RECT 758.400 643.050 759.450 644.400 ;
        RECT 757.950 642.450 760.050 643.050 ;
        RECT 757.950 642.000 762.450 642.450 ;
        RECT 757.950 641.400 763.050 642.000 ;
        RECT 757.950 640.950 760.050 641.400 ;
        RECT 760.950 637.950 763.050 641.400 ;
        RECT 764.400 633.450 765.450 644.400 ;
        RECT 769.950 643.800 772.050 645.900 ;
        RECT 766.950 640.950 769.050 643.050 ;
        RECT 767.400 637.050 768.450 640.950 ;
        RECT 766.950 634.950 769.050 637.050 ;
        RECT 770.400 634.050 771.450 643.800 ;
        RECT 764.400 632.400 768.450 633.450 ;
        RECT 757.950 619.950 760.050 622.050 ;
        RECT 763.950 619.950 766.050 622.050 ;
        RECT 751.950 610.950 754.050 613.050 ;
        RECT 748.950 604.950 751.050 607.050 ;
        RECT 758.400 606.600 759.450 619.950 ;
        RECT 764.400 606.600 765.450 619.950 ;
        RECT 767.400 619.050 768.450 632.400 ;
        RECT 769.950 631.950 772.050 634.050 ;
        RECT 773.400 631.050 774.450 650.400 ;
        RECT 769.950 628.800 772.050 630.900 ;
        RECT 772.950 628.950 775.050 631.050 ;
        RECT 766.950 616.950 769.050 619.050 ;
        RECT 770.400 615.450 771.450 628.800 ;
        RECT 776.400 621.450 777.450 658.950 ;
        RECT 778.950 652.950 781.050 655.050 ;
        RECT 791.400 654.450 792.450 658.950 ;
        RECT 788.400 653.400 792.450 654.450 ;
        RECT 779.400 640.050 780.450 652.950 ;
        RECT 788.400 651.600 789.450 653.400 ;
        RECT 788.400 649.350 789.600 651.600 ;
        RECT 793.950 650.100 796.050 652.200 ;
        RECT 794.400 649.350 795.600 650.100 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 785.400 645.900 786.600 646.650 ;
        RECT 784.950 643.800 787.050 645.900 ;
        RECT 791.400 644.400 792.600 646.650 ;
        RECT 797.400 645.900 798.600 646.650 ;
        RECT 786.000 642.750 789.000 643.050 ;
        RECT 784.950 642.300 789.000 642.750 ;
        RECT 784.950 640.950 789.450 642.300 ;
        RECT 784.950 640.650 787.050 640.950 ;
        RECT 778.950 637.950 781.050 640.050 ;
        RECT 784.950 633.450 787.050 637.050 ;
        RECT 782.400 633.000 787.050 633.450 ;
        RECT 781.950 632.400 786.450 633.000 ;
        RECT 778.950 628.950 781.050 631.050 ;
        RECT 781.950 628.950 784.050 632.400 ;
        RECT 767.400 614.400 771.450 615.450 ;
        RECT 773.400 620.400 777.450 621.450 ;
        RECT 767.400 607.050 768.450 614.400 ;
        RECT 769.950 610.950 772.050 613.050 ;
        RECT 749.400 589.050 750.450 604.950 ;
        RECT 758.400 604.350 759.600 606.600 ;
        RECT 764.400 604.350 765.600 606.600 ;
        RECT 766.950 604.950 769.050 607.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 763.950 601.950 766.050 604.050 ;
        RECT 751.950 598.800 754.050 600.900 ;
        RECT 755.400 599.400 756.600 601.650 ;
        RECT 761.400 600.900 762.600 601.650 ;
        RECT 748.950 586.950 751.050 589.050 ;
        RECT 743.400 572.400 747.450 573.450 ;
        RECT 752.400 573.600 753.450 598.800 ;
        RECT 755.400 580.050 756.450 599.400 ;
        RECT 760.950 598.800 763.050 600.900 ;
        RECT 763.950 595.950 766.050 598.050 ;
        RECT 760.950 580.950 763.050 583.050 ;
        RECT 754.950 577.950 757.050 580.050 ;
        RECT 739.950 565.800 742.050 567.900 ;
        RECT 736.950 559.950 739.050 562.050 ;
        RECT 743.400 559.050 744.450 572.400 ;
        RECT 752.400 571.350 753.600 573.600 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 749.400 567.900 750.600 568.650 ;
        RECT 748.950 565.800 751.050 567.900 ;
        RECT 755.400 566.400 756.600 568.650 ;
        RECT 755.400 562.050 756.450 566.400 ;
        RECT 754.950 559.950 757.050 562.050 ;
        RECT 742.950 556.950 745.050 559.050 ;
        RECT 761.400 556.050 762.450 580.950 ;
        RECT 764.400 567.900 765.450 595.950 ;
        RECT 766.950 592.950 769.050 595.050 ;
        RECT 763.950 565.800 766.050 567.900 ;
        RECT 760.950 553.950 763.050 556.050 ;
        RECT 767.400 546.450 768.450 592.950 ;
        RECT 770.400 589.050 771.450 610.950 ;
        RECT 773.400 595.050 774.450 620.400 ;
        RECT 775.950 616.950 778.050 619.050 ;
        RECT 772.950 592.950 775.050 595.050 ;
        RECT 772.950 589.800 775.050 591.900 ;
        RECT 769.950 586.950 772.050 589.050 ;
        RECT 773.400 577.050 774.450 589.800 ;
        RECT 776.400 586.050 777.450 616.950 ;
        RECT 779.400 598.050 780.450 628.950 ;
        RECT 788.400 613.050 789.450 640.950 ;
        RECT 791.400 622.050 792.450 644.400 ;
        RECT 796.950 643.800 799.050 645.900 ;
        RECT 799.950 643.950 802.050 646.050 ;
        RECT 793.950 640.950 796.050 643.050 ;
        RECT 790.950 619.950 793.050 622.050 ;
        RECT 787.950 610.950 790.050 613.050 ;
        RECT 781.950 606.000 784.050 610.050 ;
        RECT 790.950 606.000 793.050 610.050 ;
        RECT 782.400 604.350 783.600 606.000 ;
        RECT 791.400 604.350 792.600 606.000 ;
        RECT 782.100 601.950 784.200 604.050 ;
        RECT 787.500 601.950 789.600 604.050 ;
        RECT 790.800 601.950 792.900 604.050 ;
        RECT 788.400 600.900 789.600 601.650 ;
        RECT 787.950 598.800 790.050 600.900 ;
        RECT 778.950 595.950 781.050 598.050 ;
        RECT 794.400 597.450 795.450 640.950 ;
        RECT 797.400 640.050 798.450 643.800 ;
        RECT 796.950 637.950 799.050 640.050 ;
        RECT 796.950 631.950 799.050 634.050 ;
        RECT 791.400 596.400 795.450 597.450 ;
        RECT 787.950 586.950 790.050 589.050 ;
        RECT 775.950 583.950 778.050 586.050 ;
        RECT 772.950 574.950 775.050 577.050 ;
        RECT 775.950 572.100 778.050 574.200 ;
        RECT 776.400 571.350 777.600 572.100 ;
        RECT 784.950 571.950 787.050 574.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 773.400 567.900 774.600 568.650 ;
        RECT 772.950 565.800 775.050 567.900 ;
        RECT 779.400 566.400 780.600 568.650 ;
        RECT 775.950 562.950 778.050 565.050 ;
        RECT 772.950 550.950 775.050 553.050 ;
        RECT 767.400 545.400 771.450 546.450 ;
        RECT 770.400 541.050 771.450 545.400 ;
        RECT 769.950 538.950 772.050 541.050 ;
        RECT 733.950 535.950 736.050 538.050 ;
        RECT 754.950 535.950 757.050 538.050 ;
        RECT 730.800 532.950 732.900 535.050 ;
        RECT 727.950 527.100 730.050 529.200 ;
        RECT 731.400 496.050 732.450 532.950 ;
        RECT 733.950 529.950 736.050 534.900 ;
        RECT 739.500 531.300 741.600 533.400 ;
        RECT 749.100 532.500 751.200 534.600 ;
        RECT 736.950 527.100 739.050 529.200 ;
        RECT 737.400 526.350 738.600 527.100 ;
        RECT 737.100 523.950 739.200 526.050 ;
        RECT 733.950 520.800 736.050 522.900 ;
        RECT 740.400 522.300 741.300 531.300 ;
        RECT 742.800 527.700 744.900 529.800 ;
        RECT 746.400 529.350 747.600 531.600 ;
        RECT 744.000 525.300 744.900 527.700 ;
        RECT 745.800 526.950 747.900 529.050 ;
        RECT 749.700 525.300 750.900 532.500 ;
        RECT 744.000 524.100 750.900 525.300 ;
        RECT 747.000 522.300 749.100 523.200 ;
        RECT 740.400 521.100 749.100 522.300 ;
        RECT 730.950 493.950 733.050 496.050 ;
        RECT 728.100 490.950 730.200 493.050 ;
        RECT 728.400 488.400 729.600 490.650 ;
        RECT 728.400 487.050 729.450 488.400 ;
        RECT 727.950 484.950 730.050 487.050 ;
        RECT 724.950 466.950 727.050 469.050 ;
        RECT 721.950 457.950 724.050 460.050 ;
        RECT 718.950 454.950 721.050 457.050 ;
        RECT 715.950 451.950 718.050 454.050 ;
        RECT 719.400 450.600 720.450 454.950 ;
        RECT 722.400 451.050 723.450 457.950 ;
        RECT 728.400 454.050 729.450 484.950 ;
        RECT 734.400 480.450 735.450 520.800 ;
        RECT 741.900 519.300 744.000 521.100 ;
        RECT 745.800 518.100 747.900 520.200 ;
        RECT 750.000 518.700 750.900 524.100 ;
        RECT 751.800 523.950 753.900 526.050 ;
        RECT 752.400 522.900 753.600 523.650 ;
        RECT 751.950 520.800 754.050 522.900 ;
        RECT 755.400 520.050 756.450 535.950 ;
        RECT 769.950 532.950 772.050 535.050 ;
        RECT 757.950 529.950 760.050 532.050 ;
        RECT 746.400 515.550 747.600 517.800 ;
        RECT 749.100 516.600 751.200 518.700 ;
        RECT 754.950 517.950 757.050 520.050 ;
        RECT 746.400 511.050 747.450 515.550 ;
        RECT 745.950 508.950 748.050 511.050 ;
        RECT 739.950 493.950 742.050 496.050 ;
        RECT 734.400 479.400 738.450 480.450 ;
        RECT 737.400 454.050 738.450 479.400 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 736.950 451.950 739.050 454.050 ;
        RECT 713.400 448.350 714.600 450.600 ;
        RECT 719.400 448.350 720.600 450.600 ;
        RECT 721.950 448.950 724.050 451.050 ;
        RECT 725.100 448.950 727.200 451.050 ;
        RECT 734.100 448.950 736.200 451.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 712.950 445.950 715.050 448.050 ;
        RECT 715.950 445.950 718.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 725.400 446.400 726.600 448.650 ;
        RECT 734.400 447.900 735.600 448.650 ;
        RECT 704.400 443.400 708.450 444.450 ;
        RECT 703.950 439.950 706.050 442.050 ;
        RECT 691.950 424.950 694.050 427.050 ;
        RECT 700.950 424.950 703.050 427.050 ;
        RECT 692.400 411.900 693.450 424.950 ;
        RECT 704.400 418.200 705.450 439.950 ;
        RECT 694.950 417.600 699.000 418.050 ;
        RECT 694.950 415.950 699.600 417.600 ;
        RECT 703.950 416.100 706.050 418.200 ;
        RECT 698.400 415.350 699.600 415.950 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 701.400 411.900 702.600 412.650 ;
        RECT 707.400 412.050 708.450 443.400 ;
        RECT 710.400 443.400 711.600 445.650 ;
        RECT 716.400 444.900 717.600 445.650 ;
        RECT 691.950 409.800 694.050 411.900 ;
        RECT 700.950 409.800 703.050 411.900 ;
        RECT 703.950 409.950 706.050 412.050 ;
        RECT 706.950 409.950 709.050 412.050 ;
        RECT 701.400 406.050 702.450 409.800 ;
        RECT 700.950 403.950 703.050 406.050 ;
        RECT 689.400 392.400 693.450 393.450 ;
        RECT 688.950 388.950 691.050 391.050 ;
        RECT 677.400 370.350 678.600 372.600 ;
        RECT 682.800 370.950 684.900 373.050 ;
        RECT 685.950 370.950 688.050 373.050 ;
        RECT 673.950 367.950 676.050 370.050 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 685.950 367.800 688.050 369.900 ;
        RECT 667.950 364.950 670.050 367.050 ;
        RECT 674.400 366.900 675.600 367.650 ;
        RECT 673.950 364.800 676.050 366.900 ;
        RECT 680.400 366.000 681.600 367.650 ;
        RECT 679.950 361.950 682.050 366.000 ;
        RECT 686.400 364.050 687.450 367.800 ;
        RECT 689.400 367.050 690.450 388.950 ;
        RECT 688.950 364.950 691.050 367.050 ;
        RECT 685.950 361.950 688.050 364.050 ;
        RECT 688.950 358.950 691.050 361.050 ;
        RECT 674.400 353.400 681.450 354.450 ;
        RECT 674.400 346.050 675.450 353.400 ;
        RECT 676.950 349.950 679.050 352.050 ;
        RECT 673.950 343.950 676.050 346.050 ;
        RECT 677.400 343.050 678.450 349.950 ;
        RECT 680.400 349.050 681.450 353.400 ;
        RECT 679.950 346.950 682.050 349.050 ;
        RECT 676.950 340.950 679.050 343.050 ;
        RECT 667.950 338.100 670.050 340.200 ;
        RECT 673.950 338.100 676.050 340.200 ;
        RECT 679.950 338.100 682.050 340.200 ;
        RECT 668.400 322.050 669.450 338.100 ;
        RECT 674.400 337.350 675.600 338.100 ;
        RECT 680.400 337.350 681.600 338.100 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 676.950 334.950 679.050 337.050 ;
        RECT 679.950 334.950 682.050 337.050 ;
        RECT 682.950 334.950 685.050 337.050 ;
        RECT 670.950 331.950 673.050 334.050 ;
        RECT 677.400 333.900 678.600 334.650 ;
        RECT 667.950 319.950 670.050 322.050 ;
        RECT 646.950 286.800 649.050 288.900 ;
        RECT 643.950 271.950 646.050 274.050 ;
        RECT 619.950 268.950 622.050 271.050 ;
        RECT 622.950 265.950 625.050 268.050 ;
        RECT 613.950 260.100 616.050 262.200 ;
        RECT 614.400 259.350 615.600 260.100 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 611.400 254.400 612.600 256.650 ;
        RECT 617.400 254.400 618.600 256.650 ;
        RECT 611.400 250.050 612.450 254.400 ;
        RECT 610.950 247.950 613.050 250.050 ;
        RECT 617.400 238.050 618.450 254.400 ;
        RECT 616.950 235.950 619.050 238.050 ;
        RECT 604.950 226.950 607.050 229.050 ;
        RECT 619.950 220.950 622.050 223.050 ;
        RECT 607.950 215.100 610.050 217.200 ;
        RECT 608.400 214.350 609.600 215.100 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 605.400 210.900 606.600 211.650 ;
        RECT 598.950 208.800 601.050 210.900 ;
        RECT 604.950 208.800 607.050 210.900 ;
        RECT 611.400 209.400 612.600 211.650 ;
        RECT 599.400 184.200 600.450 208.800 ;
        RECT 611.400 190.050 612.450 209.400 ;
        RECT 620.400 199.050 621.450 220.950 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 610.950 187.950 613.050 190.050 ;
        RECT 584.400 181.350 585.600 183.600 ;
        RECT 590.400 181.350 591.600 183.600 ;
        RECT 598.950 182.100 601.050 184.200 ;
        RECT 611.400 183.450 612.600 183.600 ;
        RECT 605.400 182.400 612.600 183.450 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 587.400 176.400 588.600 178.650 ;
        RECT 593.400 176.400 594.600 178.650 ;
        RECT 587.400 172.050 588.450 176.400 ;
        RECT 586.950 169.950 589.050 172.050 ;
        RECT 577.950 154.950 580.050 157.050 ;
        RECT 593.400 151.050 594.450 176.400 ;
        RECT 601.950 169.950 604.050 172.050 ;
        RECT 592.950 148.950 595.050 151.050 ;
        RECT 598.950 145.950 601.050 148.050 ;
        RECT 592.950 137.100 595.050 139.200 ;
        RECT 599.400 139.050 600.450 145.950 ;
        RECT 593.400 136.350 594.600 137.100 ;
        RECT 598.950 136.950 601.050 139.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 590.400 132.000 591.600 133.650 ;
        RECT 566.400 126.000 567.600 127.800 ;
        RECT 569.100 126.600 571.200 128.700 ;
        RECT 574.950 127.950 577.050 130.050 ;
        RECT 565.950 121.950 568.050 126.000 ;
        RECT 578.400 118.050 579.450 130.800 ;
        RECT 583.950 127.950 586.050 130.050 ;
        RECT 589.950 127.950 592.050 132.000 ;
        RECT 577.950 115.950 580.050 118.050 ;
        RECT 571.950 112.950 574.050 115.050 ;
        RECT 553.950 106.950 556.050 109.050 ;
        RECT 554.400 99.900 555.450 106.950 ;
        RECT 556.950 104.100 559.050 106.200 ;
        RECT 565.950 104.100 568.050 106.200 ;
        RECT 572.400 105.600 573.450 112.950 ;
        RECT 574.950 109.950 577.050 112.050 ;
        RECT 575.400 106.050 576.450 109.950 ;
        RECT 548.400 98.400 552.450 99.450 ;
        RECT 548.400 88.050 549.450 98.400 ;
        RECT 553.950 97.800 556.050 99.900 ;
        RECT 547.950 85.950 550.050 88.050 ;
        RECT 557.400 85.050 558.450 104.100 ;
        RECT 566.400 103.350 567.600 104.100 ;
        RECT 572.400 103.350 573.600 105.600 ;
        RECT 574.950 103.950 577.050 106.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 565.950 100.950 568.050 103.050 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 563.400 99.900 564.600 100.650 ;
        RECT 562.950 97.800 565.050 99.900 ;
        RECT 569.400 98.400 570.600 100.650 ;
        RECT 532.950 82.950 535.050 85.050 ;
        RECT 556.950 82.950 559.050 85.050 ;
        RECT 523.950 76.950 526.050 79.050 ;
        RECT 514.950 64.950 517.050 67.050 ;
        RECT 505.950 43.800 508.050 45.900 ;
        RECT 511.950 43.950 514.050 46.050 ;
        RECT 490.950 28.950 493.050 31.050 ;
        RECT 481.950 26.100 484.050 28.200 ;
        RECT 506.400 27.600 507.450 43.800 ;
        RECT 515.400 34.050 516.450 64.950 ;
        RECT 521.400 60.450 522.600 60.600 ;
        RECT 518.400 59.400 522.600 60.450 ;
        RECT 518.400 37.050 519.450 59.400 ;
        RECT 521.400 58.350 522.600 59.400 ;
        RECT 530.400 60.450 531.600 60.600 ;
        RECT 533.400 60.450 534.450 82.950 ;
        RECT 544.950 79.950 547.050 82.050 ;
        RECT 541.950 61.950 544.050 64.050 ;
        RECT 530.400 59.400 534.450 60.450 ;
        RECT 530.400 58.350 531.600 59.400 ;
        RECT 521.100 55.950 523.200 58.050 ;
        RECT 526.500 55.950 528.600 58.050 ;
        RECT 529.800 55.950 531.900 58.050 ;
        RECT 527.400 54.900 528.600 55.650 ;
        RECT 526.950 52.800 529.050 54.900 ;
        RECT 533.400 46.050 534.450 59.400 ;
        RECT 532.950 43.950 535.050 46.050 ;
        RECT 517.950 34.950 520.050 37.050 ;
        RECT 514.950 31.950 517.050 34.050 ;
        RECT 482.400 25.350 483.600 26.100 ;
        RECT 506.400 25.350 507.600 27.600 ;
        RECT 526.950 27.000 529.050 31.050 ;
        RECT 538.950 28.950 541.050 31.050 ;
        RECT 527.400 25.350 528.600 27.000 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 479.400 21.900 480.600 22.650 ;
        RECT 437.100 14.400 439.200 16.500 ;
        RECT 461.400 16.050 462.450 20.400 ;
        RECT 472.950 19.800 475.050 21.900 ;
        RECT 478.950 19.800 481.050 21.900 ;
        RECT 485.400 20.400 486.600 22.650 ;
        RECT 503.400 20.400 504.600 22.650 ;
        RECT 509.400 21.900 510.600 22.650 ;
        RECT 530.400 21.900 531.600 22.650 ;
        RECT 485.400 16.050 486.450 20.400 ;
        RECT 503.400 16.050 504.450 20.400 ;
        RECT 508.950 19.800 511.050 21.900 ;
        RECT 529.950 19.800 532.050 21.900 ;
        RECT 530.400 16.050 531.450 19.800 ;
        RECT 539.400 19.050 540.450 28.950 ;
        RECT 538.950 16.950 541.050 19.050 ;
        RECT 460.950 13.950 463.050 16.050 ;
        RECT 484.950 13.950 487.050 16.050 ;
        RECT 502.950 13.950 505.050 16.050 ;
        RECT 529.950 13.950 532.050 16.050 ;
        RECT 370.950 10.950 373.050 13.050 ;
        RECT 418.950 10.950 421.050 13.050 ;
        RECT 358.200 6.600 360.300 8.700 ;
        RECT 371.400 7.050 372.450 10.950 ;
        RECT 542.400 7.050 543.450 61.950 ;
        RECT 545.400 54.900 546.450 79.950 ;
        RECT 569.400 73.050 570.450 98.400 ;
        RECT 568.950 70.950 571.050 73.050 ;
        RECT 578.400 67.050 579.450 115.950 ;
        RECT 580.950 103.950 583.050 106.050 ;
        RECT 581.400 82.050 582.450 103.950 ;
        RECT 584.400 99.900 585.450 127.950 ;
        RECT 592.950 124.950 595.050 127.050 ;
        RECT 593.400 105.600 594.450 124.950 ;
        RECT 599.400 106.050 600.450 136.950 ;
        RECT 593.400 103.350 594.600 105.600 ;
        RECT 598.950 103.950 601.050 106.050 ;
        RECT 589.950 100.950 592.050 103.050 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 590.400 99.900 591.600 100.650 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 589.950 97.800 592.050 99.900 ;
        RECT 596.400 98.400 597.600 100.650 ;
        RECT 584.400 91.050 585.450 97.800 ;
        RECT 583.950 88.950 586.050 91.050 ;
        RECT 596.400 85.050 597.450 98.400 ;
        RECT 602.400 97.050 603.450 169.950 ;
        RECT 605.400 145.050 606.450 182.400 ;
        RECT 611.400 181.350 612.600 182.400 ;
        RECT 616.950 182.100 619.050 184.200 ;
        RECT 617.400 181.350 618.600 182.100 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 614.400 177.900 615.600 178.650 ;
        RECT 613.950 175.800 616.050 177.900 ;
        RECT 619.950 157.950 622.050 160.050 ;
        RECT 613.950 154.950 616.050 157.050 ;
        RECT 604.950 142.950 607.050 145.050 ;
        RECT 614.400 138.600 615.450 154.950 ;
        RECT 620.400 138.600 621.450 157.950 ;
        RECT 623.400 139.200 624.450 265.950 ;
        RECT 644.400 262.200 645.450 271.950 ;
        RECT 628.950 259.950 631.050 262.050 ;
        RECT 637.950 260.100 640.050 262.200 ;
        RECT 643.950 260.100 646.050 262.200 ;
        RECT 629.400 216.600 630.450 259.950 ;
        RECT 638.400 259.350 639.600 260.100 ;
        RECT 644.400 259.350 645.600 260.100 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 640.950 256.950 643.050 259.050 ;
        RECT 643.950 256.950 646.050 259.050 ;
        RECT 635.400 254.400 636.600 256.650 ;
        RECT 641.400 255.900 642.600 256.650 ;
        RECT 635.400 226.050 636.450 254.400 ;
        RECT 640.950 253.800 643.050 255.900 ;
        RECT 650.400 244.050 651.450 293.100 ;
        RECT 659.400 292.350 660.600 294.600 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 665.400 292.350 666.600 293.100 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 656.400 287.400 657.600 289.650 ;
        RECT 662.400 288.900 663.600 289.650 ;
        RECT 656.400 274.050 657.450 287.400 ;
        RECT 661.950 286.800 664.050 288.900 ;
        RECT 655.950 271.950 658.050 274.050 ;
        RECT 671.400 268.050 672.450 331.950 ;
        RECT 676.950 331.800 679.050 333.900 ;
        RECT 683.400 332.400 684.600 334.650 ;
        RECT 683.400 331.050 684.450 332.400 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 679.950 328.950 684.450 331.050 ;
        RECT 679.950 322.950 682.050 325.050 ;
        RECT 680.400 316.050 681.450 322.950 ;
        RECT 679.950 313.950 682.050 316.050 ;
        RECT 683.400 307.050 684.450 328.950 ;
        RECT 682.950 304.950 685.050 307.050 ;
        RECT 676.950 298.950 679.050 301.050 ;
        RECT 673.950 292.950 676.050 295.050 ;
        RECT 655.950 265.950 658.050 268.050 ;
        RECT 670.950 265.950 673.050 268.050 ;
        RECT 656.400 255.900 657.450 265.950 ;
        RECT 661.950 260.100 664.050 262.200 ;
        RECT 667.950 260.100 670.050 262.200 ;
        RECT 674.400 261.450 675.450 292.950 ;
        RECT 677.400 268.050 678.450 298.950 ;
        RECT 686.400 297.450 687.450 331.950 ;
        RECT 689.400 298.200 690.450 358.950 ;
        RECT 692.400 301.050 693.450 392.400 ;
        RECT 704.400 385.050 705.450 409.950 ;
        RECT 710.400 391.050 711.450 443.400 ;
        RECT 715.950 442.800 718.050 444.900 ;
        RECT 725.400 439.050 726.450 446.400 ;
        RECT 733.800 445.800 735.900 447.900 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 727.950 439.950 730.050 442.050 ;
        RECT 724.950 436.950 727.050 439.050 ;
        RECT 724.950 430.950 727.050 433.050 ;
        RECT 725.400 424.050 726.450 430.950 ;
        RECT 715.950 421.950 718.050 424.050 ;
        RECT 724.950 421.950 727.050 424.050 ;
        RECT 728.400 423.450 729.450 439.950 ;
        RECT 712.950 412.950 715.050 418.050 ;
        RECT 712.950 409.800 715.050 411.900 ;
        RECT 713.400 400.050 714.450 409.800 ;
        RECT 712.950 397.950 715.050 400.050 ;
        RECT 709.950 388.950 712.050 391.050 ;
        RECT 694.950 382.950 697.050 385.050 ;
        RECT 703.950 382.950 706.050 385.050 ;
        RECT 695.400 313.050 696.450 382.950 ;
        RECT 700.800 376.500 702.900 378.600 ;
        RECT 698.100 367.950 700.200 370.050 ;
        RECT 701.100 369.300 702.300 376.500 ;
        RECT 704.400 373.350 705.600 375.600 ;
        RECT 710.400 375.300 712.500 377.400 ;
        RECT 704.100 370.950 706.200 373.050 ;
        RECT 707.100 371.700 709.200 373.800 ;
        RECT 707.100 369.300 708.000 371.700 ;
        RECT 701.100 368.100 708.000 369.300 ;
        RECT 698.400 366.900 699.600 367.650 ;
        RECT 697.950 364.800 700.050 366.900 ;
        RECT 701.100 362.700 702.000 368.100 ;
        RECT 702.900 366.300 705.000 367.200 ;
        RECT 710.700 366.300 711.600 375.300 ;
        RECT 712.950 371.100 715.050 373.200 ;
        RECT 713.400 370.350 714.600 371.100 ;
        RECT 712.800 367.950 714.900 370.050 ;
        RECT 702.900 365.100 711.600 366.300 ;
        RECT 700.800 360.600 702.900 362.700 ;
        RECT 704.100 362.100 706.200 364.200 ;
        RECT 708.000 363.300 710.100 365.100 ;
        RECT 704.400 361.050 705.600 361.800 ;
        RECT 703.950 358.950 706.050 361.050 ;
        RECT 697.950 352.950 700.050 355.050 ;
        RECT 698.400 339.450 699.450 352.950 ;
        RECT 716.400 349.050 717.450 421.950 ;
        RECT 728.400 421.200 729.600 423.450 ;
        RECT 723.900 417.900 726.000 419.700 ;
        RECT 727.800 418.800 729.900 420.900 ;
        RECT 731.100 420.300 733.200 422.400 ;
        RECT 722.400 416.700 731.100 417.900 ;
        RECT 719.100 412.950 721.200 415.050 ;
        RECT 719.400 411.900 720.600 412.650 ;
        RECT 718.950 409.800 721.050 411.900 ;
        RECT 722.400 407.700 723.300 416.700 ;
        RECT 729.000 415.800 731.100 416.700 ;
        RECT 732.000 414.900 732.900 420.300 ;
        RECT 733.950 416.100 736.050 418.200 ;
        RECT 734.400 415.350 735.600 416.100 ;
        RECT 726.000 413.700 732.900 414.900 ;
        RECT 726.000 411.300 726.900 413.700 ;
        RECT 724.800 409.200 726.900 411.300 ;
        RECT 727.800 409.950 729.900 412.050 ;
        RECT 721.500 405.600 723.600 407.700 ;
        RECT 728.400 407.400 729.600 409.650 ;
        RECT 731.700 406.500 732.900 413.700 ;
        RECT 733.800 412.950 735.900 415.050 ;
        RECT 731.100 404.400 733.200 406.500 ;
        RECT 737.400 400.050 738.450 445.950 ;
        RECT 740.400 442.050 741.450 493.950 ;
        RECT 758.400 493.050 759.450 529.950 ;
        RECT 770.400 528.600 771.450 532.950 ;
        RECT 773.400 532.050 774.450 550.950 ;
        RECT 776.400 544.050 777.450 562.950 ;
        RECT 779.400 559.050 780.450 566.400 ;
        RECT 781.950 565.950 784.050 568.050 ;
        RECT 782.400 562.050 783.450 565.950 ;
        RECT 781.950 559.950 784.050 562.050 ;
        RECT 778.800 556.950 780.900 559.050 ;
        RECT 781.950 556.800 784.050 558.900 ;
        RECT 775.950 541.950 778.050 544.050 ;
        RECT 772.950 529.950 775.050 532.050 ;
        RECT 770.400 526.350 771.600 528.600 ;
        RECT 778.950 528.450 781.050 529.200 ;
        RECT 782.400 528.450 783.450 556.800 ;
        RECT 785.400 553.050 786.450 571.950 ;
        RECT 784.950 550.950 787.050 553.050 ;
        RECT 778.950 527.400 783.450 528.450 ;
        RECT 778.950 527.100 781.050 527.400 ;
        RECT 779.400 526.350 780.600 527.100 ;
        RECT 770.100 523.950 772.200 526.050 ;
        RECT 775.500 523.950 777.600 526.050 ;
        RECT 778.800 523.950 780.900 526.050 ;
        RECT 776.400 521.400 777.600 523.650 ;
        RECT 782.400 523.050 783.450 527.400 ;
        RECT 784.950 526.950 787.050 529.050 ;
        RECT 776.400 520.050 777.450 521.400 ;
        RECT 781.950 520.950 784.050 523.050 ;
        RECT 785.400 520.050 786.450 526.950 ;
        RECT 788.400 526.050 789.450 586.950 ;
        RECT 787.950 523.950 790.050 526.050 ;
        RECT 776.400 518.400 781.050 520.050 ;
        RECT 777.000 517.950 781.050 518.400 ;
        RECT 784.950 517.950 787.050 520.050 ;
        RECT 785.400 514.050 786.450 517.950 ;
        RECT 784.950 511.950 787.050 514.050 ;
        RECT 791.400 511.050 792.450 596.400 ;
        RECT 797.400 592.050 798.450 631.950 ;
        RECT 800.400 607.200 801.450 643.950 ;
        RECT 803.400 628.050 804.450 673.950 ;
        RECT 805.950 670.950 808.050 674.400 ;
        RECT 808.950 673.950 811.050 674.400 ;
        RECT 802.950 625.950 805.050 628.050 ;
        RECT 803.400 622.050 804.450 625.950 ;
        RECT 802.950 619.950 805.050 622.050 ;
        RECT 802.950 616.800 805.050 618.900 ;
        RECT 799.950 605.100 802.050 607.200 ;
        RECT 800.400 601.050 801.450 605.100 ;
        RECT 799.950 598.950 802.050 601.050 ;
        RECT 796.950 589.950 799.050 592.050 ;
        RECT 799.950 583.950 802.050 586.050 ;
        RECT 800.400 573.600 801.450 583.950 ;
        RECT 800.400 571.350 801.600 573.600 ;
        RECT 803.400 573.450 804.450 616.800 ;
        RECT 806.400 616.050 807.450 670.950 ;
        RECT 808.950 670.800 811.050 672.900 ;
        RECT 809.400 643.050 810.450 670.800 ;
        RECT 812.400 652.050 813.450 676.950 ;
        RECT 815.400 676.050 816.450 694.950 ;
        RECT 814.950 673.950 817.050 676.050 ;
        RECT 818.400 673.050 819.450 722.400 ;
        RECT 821.400 722.400 822.600 724.650 ;
        RECT 827.400 723.000 828.600 724.650 ;
        RECT 821.400 694.050 822.450 722.400 ;
        RECT 826.950 718.950 829.050 723.000 ;
        RECT 826.950 706.950 829.050 709.050 ;
        RECT 823.950 694.950 826.050 697.050 ;
        RECT 820.950 691.950 823.050 694.050 ;
        RECT 817.950 670.950 820.050 673.050 ;
        RECT 821.400 670.050 822.450 691.950 ;
        RECT 824.400 685.050 825.450 694.950 ;
        RECT 827.400 691.050 828.450 706.950 ;
        RECT 839.400 694.050 840.450 727.950 ;
        RECT 838.950 691.950 841.050 694.050 ;
        RECT 826.950 688.950 829.050 691.050 ;
        RECT 823.800 682.950 825.900 685.050 ;
        RECT 826.950 683.100 829.050 685.200 ;
        RECT 827.400 682.350 828.600 683.100 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 830.400 678.900 831.600 679.650 ;
        RECT 829.950 676.800 832.050 678.900 ;
        RECT 823.950 673.950 829.050 676.050 ;
        RECT 823.950 670.800 826.050 672.900 ;
        RECT 820.950 667.950 823.050 670.050 ;
        RECT 814.950 664.950 817.050 667.050 ;
        RECT 815.400 652.200 816.450 664.950 ;
        RECT 811.950 649.950 814.050 652.050 ;
        RECT 814.950 650.100 817.050 652.200 ;
        RECT 820.950 651.000 823.050 655.050 ;
        RECT 824.400 652.050 825.450 670.800 ;
        RECT 836.400 661.050 837.450 679.950 ;
        RECT 838.950 676.800 841.050 678.900 ;
        RECT 826.950 658.950 829.050 661.050 ;
        RECT 835.950 658.950 838.050 661.050 ;
        RECT 815.400 649.350 816.600 650.100 ;
        RECT 821.400 649.350 822.600 651.000 ;
        RECT 823.950 649.950 826.050 652.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 818.400 644.400 819.600 646.650 ;
        RECT 808.950 640.950 811.050 643.050 ;
        RECT 818.400 640.050 819.450 644.400 ;
        RECT 820.950 640.950 823.050 643.050 ;
        RECT 817.950 637.950 820.050 640.050 ;
        RECT 805.950 613.950 808.050 616.050 ;
        RECT 805.950 606.600 810.000 607.050 ;
        RECT 805.950 604.950 810.600 606.600 ;
        RECT 814.950 605.100 817.050 607.200 ;
        RECT 809.400 604.350 810.600 604.950 ;
        RECT 815.400 604.350 816.600 605.100 ;
        RECT 821.400 604.050 822.450 640.950 ;
        RECT 827.400 613.050 828.450 658.950 ;
        RECT 832.950 652.950 835.050 655.050 ;
        RECT 829.950 649.950 832.050 652.050 ;
        RECT 826.950 610.950 829.050 613.050 ;
        RECT 823.950 604.950 826.050 607.050 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 805.950 598.950 808.050 601.050 ;
        RECT 812.400 599.400 813.600 601.650 ;
        RECT 806.400 576.450 807.450 598.950 ;
        RECT 812.400 598.050 813.450 599.400 ;
        RECT 817.950 598.950 820.050 601.050 ;
        RECT 812.400 596.400 817.050 598.050 ;
        RECT 813.000 595.950 817.050 596.400 ;
        RECT 818.400 594.450 819.450 598.950 ;
        RECT 815.400 593.400 819.450 594.450 ;
        RECT 811.950 577.950 814.050 580.050 ;
        RECT 806.400 575.400 810.450 576.450 ;
        RECT 803.400 572.400 807.450 573.450 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 797.400 566.400 798.600 568.650 ;
        RECT 797.400 546.450 798.450 566.400 ;
        RECT 794.400 545.400 798.450 546.450 ;
        RECT 794.400 529.050 795.450 545.400 ;
        RECT 799.950 544.950 802.050 547.050 ;
        RECT 793.950 526.950 796.050 529.050 ;
        RECT 800.400 528.600 801.450 544.950 ;
        RECT 806.400 529.050 807.450 572.400 ;
        RECT 809.400 565.050 810.450 575.400 ;
        RECT 812.400 567.900 813.450 577.950 ;
        RECT 811.950 565.800 814.050 567.900 ;
        RECT 808.950 562.950 811.050 565.050 ;
        RECT 808.950 559.800 811.050 561.900 ;
        RECT 800.400 526.350 801.600 528.600 ;
        RECT 805.950 526.950 808.050 529.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 793.950 520.800 796.050 523.050 ;
        RECT 797.400 522.000 798.600 523.650 ;
        RECT 803.400 522.900 804.600 523.650 ;
        RECT 809.400 523.050 810.450 559.800 ;
        RECT 812.400 538.050 813.450 565.800 ;
        RECT 815.400 562.050 816.450 593.400 ;
        RECT 817.950 589.950 820.050 592.050 ;
        RECT 818.400 577.050 819.450 589.950 ;
        RECT 821.400 580.050 822.450 601.950 ;
        RECT 824.400 601.050 825.450 604.950 ;
        RECT 827.400 604.050 828.450 610.950 ;
        RECT 830.400 607.050 831.450 649.950 ;
        RECT 833.400 610.050 834.450 652.950 ;
        RECT 839.400 652.050 840.450 676.800 ;
        RECT 842.400 655.050 843.450 742.950 ;
        RECT 845.400 739.050 846.450 754.950 ;
        RECT 844.950 736.950 847.050 739.050 ;
        RECT 848.400 736.050 849.450 760.950 ;
        RECT 851.400 745.050 852.450 787.950 ;
        RECT 854.400 769.050 855.450 829.950 ;
        RECT 860.400 829.050 861.450 833.400 ;
        RECT 862.950 832.950 865.050 835.050 ;
        RECT 865.950 832.950 868.050 835.050 ;
        RECT 868.950 832.950 871.050 835.050 ;
        RECT 859.950 826.950 862.050 829.050 ;
        RECT 856.950 823.950 859.050 826.050 ;
        RECT 857.400 808.200 858.450 823.950 ;
        RECT 863.400 820.050 864.450 832.950 ;
        RECT 868.950 823.950 871.050 826.050 ;
        RECT 865.950 820.950 868.050 823.050 ;
        RECT 862.950 817.950 865.050 820.050 ;
        RECT 866.400 811.050 867.450 820.950 ;
        RECT 865.950 808.950 868.050 811.050 ;
        RECT 856.950 806.100 859.050 808.200 ;
        RECT 862.950 806.100 865.050 808.200 ;
        RECT 869.400 807.600 870.450 823.950 ;
        RECT 872.400 823.050 873.450 838.950 ;
        RECT 881.400 838.350 882.600 839.100 ;
        RECT 887.400 838.350 888.600 840.600 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 878.400 833.400 879.600 835.650 ;
        RECT 884.400 834.900 885.600 835.650 ;
        RECT 871.950 820.950 874.050 823.050 ;
        RECT 878.400 817.050 879.450 833.400 ;
        RECT 883.950 832.800 886.050 834.900 ;
        RECT 880.950 829.950 883.050 832.050 ;
        RECT 889.950 829.950 892.050 832.050 ;
        RECT 877.950 814.950 880.050 817.050 ;
        RECT 877.950 808.950 880.050 811.050 ;
        RECT 857.400 796.050 858.450 806.100 ;
        RECT 863.400 805.350 864.600 806.100 ;
        RECT 869.400 805.350 870.600 807.600 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 865.950 802.950 868.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 859.950 799.950 862.050 802.050 ;
        RECT 866.400 801.000 867.600 802.650 ;
        RECT 856.950 793.950 859.050 796.050 ;
        RECT 856.950 790.800 859.050 792.900 ;
        RECT 857.400 781.050 858.450 790.800 ;
        RECT 860.400 786.450 861.450 799.950 ;
        RECT 865.950 796.950 868.050 801.000 ;
        RECT 872.400 800.400 873.600 802.650 ;
        RECT 868.950 796.950 871.050 799.050 ;
        RECT 860.400 785.400 864.450 786.450 ;
        RECT 859.950 781.950 862.050 784.050 ;
        RECT 856.950 778.950 859.050 781.050 ;
        RECT 853.950 766.950 856.050 769.050 ;
        RECT 853.800 761.100 855.900 763.200 ;
        RECT 850.950 742.950 853.050 745.050 ;
        RECT 854.400 742.050 855.450 761.100 ;
        RECT 856.950 760.950 859.050 763.050 ;
        RECT 860.400 762.600 861.450 781.950 ;
        RECT 863.400 781.050 864.450 785.400 ;
        RECT 862.950 778.950 865.050 781.050 ;
        RECT 865.950 766.950 868.050 769.050 ;
        RECT 860.400 760.350 861.600 762.600 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 863.400 756.900 864.600 757.650 ;
        RECT 862.950 754.800 865.050 756.900 ;
        RECT 869.400 754.050 870.450 796.950 ;
        RECT 872.400 775.050 873.450 800.400 ;
        RECT 881.400 799.050 882.450 829.950 ;
        RECT 886.950 826.950 889.050 829.050 ;
        RECT 887.400 814.050 888.450 826.950 ;
        RECT 890.400 820.050 891.450 829.950 ;
        RECT 889.950 817.950 892.050 820.050 ;
        RECT 893.400 817.050 894.450 850.950 ;
        RECT 895.950 847.950 898.050 850.050 ;
        RECT 896.400 835.050 897.450 847.950 ;
        RECT 895.950 832.950 898.050 835.050 ;
        RECT 892.950 814.950 895.050 817.050 ;
        RECT 886.950 811.950 889.050 814.050 ;
        RECT 889.950 806.100 892.050 811.050 ;
        RECT 895.950 807.000 898.050 811.050 ;
        RECT 899.400 807.450 900.450 851.400 ;
        RECT 913.950 850.950 916.050 853.050 ;
        RECT 914.400 841.200 915.450 850.950 ;
        RECT 926.400 847.050 927.450 883.950 ;
        RECT 929.400 879.900 930.450 895.950 ;
        RECT 932.400 886.050 933.450 911.400 ;
        RECT 934.950 910.950 937.050 911.400 ;
        RECT 944.400 911.400 945.600 913.650 ;
        RECT 944.400 910.050 945.450 911.400 ;
        RECT 949.950 910.950 952.050 913.050 ;
        RECT 944.400 908.400 949.050 910.050 ;
        RECT 945.000 907.950 949.050 908.400 ;
        RECT 950.400 892.050 951.450 910.950 ;
        RECT 940.950 889.950 943.050 892.050 ;
        RECT 949.950 889.950 952.050 892.050 ;
        RECT 931.800 883.950 933.900 886.050 ;
        RECT 934.950 884.100 937.050 886.200 ;
        RECT 941.400 885.600 942.450 889.950 ;
        RECT 935.400 883.350 936.600 884.100 ;
        RECT 941.400 883.350 942.600 885.600 ;
        RECT 949.950 883.950 952.050 886.050 ;
        RECT 934.950 880.950 937.050 883.050 ;
        RECT 937.950 880.950 940.050 883.050 ;
        RECT 940.950 880.950 943.050 883.050 ;
        RECT 943.950 880.950 946.050 883.050 ;
        RECT 938.400 879.900 939.600 880.650 ;
        RECT 944.400 879.900 945.600 880.650 ;
        RECT 928.950 877.800 931.050 879.900 ;
        RECT 937.950 877.800 940.050 879.900 ;
        RECT 943.950 877.800 946.050 879.900 ;
        RECT 950.400 874.050 951.450 883.950 ;
        RECT 953.400 877.050 954.450 919.950 ;
        RECT 952.950 874.950 955.050 877.050 ;
        RECT 928.950 871.950 931.050 874.050 ;
        RECT 949.950 871.950 952.050 874.050 ;
        RECT 929.400 862.050 930.450 871.950 ;
        RECT 956.400 871.050 957.450 952.950 ;
        RECT 973.950 925.950 976.050 928.050 ;
        RECT 958.950 917.100 961.050 919.200 ;
        RECT 967.950 917.100 970.050 919.200 ;
        RECT 974.400 918.600 975.450 925.950 ;
        RECT 959.400 910.050 960.450 917.100 ;
        RECT 968.400 916.350 969.600 917.100 ;
        RECT 974.400 916.350 975.600 918.600 ;
        RECT 964.950 913.950 967.050 916.050 ;
        RECT 967.950 913.950 970.050 916.050 ;
        RECT 970.950 913.950 973.050 916.050 ;
        RECT 973.950 913.950 976.050 916.050 ;
        RECT 965.400 911.400 966.600 913.650 ;
        RECT 971.400 911.400 972.600 913.650 ;
        RECT 958.950 907.950 961.050 910.050 ;
        RECT 965.400 904.050 966.450 911.400 ;
        RECT 971.400 907.050 972.450 911.400 ;
        RECT 970.950 904.950 973.050 907.050 ;
        RECT 964.950 901.950 967.050 904.050 ;
        RECT 964.950 892.950 967.050 895.050 ;
        RECT 965.400 885.600 966.450 892.950 ;
        RECT 965.400 883.350 966.600 885.600 ;
        RECT 970.950 884.100 973.050 886.200 ;
        RECT 971.400 883.350 972.600 884.100 ;
        RECT 976.950 883.950 979.050 886.050 ;
        RECT 961.950 880.950 964.050 883.050 ;
        RECT 964.950 880.950 967.050 883.050 ;
        RECT 967.950 880.950 970.050 883.050 ;
        RECT 970.950 880.950 973.050 883.050 ;
        RECT 962.400 878.400 963.600 880.650 ;
        RECT 968.400 879.900 969.600 880.650 ;
        RECT 962.400 871.050 963.450 878.400 ;
        RECT 967.950 877.800 970.050 879.900 ;
        RECT 977.400 877.050 978.450 883.950 ;
        RECT 976.950 874.950 979.050 877.050 ;
        RECT 967.950 871.950 970.050 874.050 ;
        RECT 943.950 865.950 946.050 871.050 ;
        RECT 949.950 868.800 952.050 870.900 ;
        RECT 955.950 868.950 958.050 871.050 ;
        RECT 961.950 868.950 964.050 871.050 ;
        RECT 928.950 859.950 931.050 862.050 ;
        RECT 946.950 853.950 949.050 856.050 ;
        RECT 919.950 844.950 922.050 847.050 ;
        RECT 925.950 844.950 928.050 847.050 ;
        RECT 907.950 839.100 910.050 841.200 ;
        RECT 913.950 839.100 916.050 841.200 ;
        RECT 908.400 838.350 909.600 839.100 ;
        RECT 914.400 838.350 915.600 839.100 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 907.950 835.950 910.050 838.050 ;
        RECT 910.950 835.950 913.050 838.050 ;
        RECT 913.950 835.950 916.050 838.050 ;
        RECT 905.400 833.400 906.600 835.650 ;
        RECT 911.400 833.400 912.600 835.650 ;
        RECT 905.400 823.050 906.450 833.400 ;
        RECT 904.950 820.950 907.050 823.050 ;
        RECT 904.950 814.950 907.050 817.050 ;
        RECT 890.400 805.350 891.600 806.100 ;
        RECT 896.400 805.350 897.600 807.000 ;
        RECT 899.400 806.400 903.450 807.450 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 895.950 802.950 898.050 805.050 ;
        RECT 886.950 799.950 889.050 802.050 ;
        RECT 893.400 801.900 894.600 802.650 ;
        RECT 880.950 796.950 883.050 799.050 ;
        RECT 877.950 793.950 880.050 796.050 ;
        RECT 871.950 772.950 874.050 775.050 ;
        RECT 874.950 766.950 877.050 772.050 ;
        RECT 871.950 763.950 874.050 766.050 ;
        RECT 868.950 751.950 871.050 754.050 ;
        RECT 872.400 751.050 873.450 763.950 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 871.950 748.950 874.050 751.050 ;
        RECT 865.950 745.950 868.050 748.050 ;
        RECT 859.950 742.950 862.050 745.050 ;
        RECT 853.950 739.950 856.050 742.050 ;
        RECT 847.950 733.950 850.050 736.050 ;
        RECT 853.950 733.950 856.050 736.050 ;
        RECT 847.950 728.100 850.050 730.200 ;
        RECT 854.400 729.600 855.450 733.950 ;
        RECT 848.400 727.350 849.600 728.100 ;
        RECT 854.400 727.350 855.600 729.600 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 851.400 723.900 852.600 724.650 ;
        RECT 850.950 721.800 853.050 723.900 ;
        RECT 847.950 718.950 850.050 721.050 ;
        RECT 848.400 709.050 849.450 718.950 ;
        RECT 847.950 706.950 850.050 709.050 ;
        RECT 844.950 703.950 847.050 706.050 ;
        RECT 845.400 688.050 846.450 703.950 ;
        RECT 847.950 700.950 850.050 703.050 ;
        RECT 848.400 697.050 849.450 700.950 ;
        RECT 847.950 694.950 850.050 697.050 ;
        RECT 856.950 694.950 859.050 697.050 ;
        RECT 844.950 682.950 847.050 688.050 ;
        RECT 847.950 683.100 850.050 685.200 ;
        RECT 853.950 683.100 856.050 685.200 ;
        RECT 857.400 685.050 858.450 694.950 ;
        RECT 848.400 682.350 849.600 683.100 ;
        RECT 854.400 682.350 855.600 683.100 ;
        RECT 856.950 682.950 859.050 685.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 851.400 678.000 852.600 679.650 ;
        RECT 850.950 673.950 853.050 678.000 ;
        RECT 856.950 676.950 859.050 679.050 ;
        RECT 853.950 673.950 856.050 676.050 ;
        RECT 854.400 663.450 855.450 673.950 ;
        RECT 857.400 673.050 858.450 676.950 ;
        RECT 856.950 670.950 859.050 673.050 ;
        RECT 851.400 662.400 855.450 663.450 ;
        RECT 841.950 652.950 844.050 655.050 ;
        RECT 835.950 651.600 840.450 652.050 ;
        RECT 835.950 649.950 840.600 651.600 ;
        RECT 844.950 651.000 847.050 655.050 ;
        RECT 851.400 652.050 852.450 662.400 ;
        RECT 853.950 658.950 856.050 661.050 ;
        RECT 839.400 649.350 840.600 649.950 ;
        RECT 845.400 649.350 846.600 651.000 ;
        RECT 850.950 649.950 853.050 652.050 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 835.950 643.950 838.050 646.050 ;
        RECT 842.400 645.900 843.600 646.650 ;
        RECT 836.400 613.050 837.450 643.950 ;
        RECT 841.950 643.800 844.050 645.900 ;
        RECT 848.400 644.400 849.600 646.650 ;
        RECT 844.950 637.950 847.050 640.050 ;
        RECT 845.400 628.050 846.450 637.950 ;
        RECT 844.950 625.950 847.050 628.050 ;
        RECT 848.400 625.050 849.450 644.400 ;
        RECT 850.950 643.950 853.050 646.050 ;
        RECT 851.400 631.050 852.450 643.950 ;
        RECT 850.950 628.950 853.050 631.050 ;
        RECT 847.950 622.950 850.050 625.050 ;
        RECT 844.950 619.950 847.050 622.050 ;
        RECT 835.950 610.950 838.050 613.050 ;
        RECT 841.950 610.950 844.050 613.050 ;
        RECT 832.950 607.950 835.050 610.050 ;
        RECT 829.950 604.950 832.050 607.050 ;
        RECT 835.950 605.100 838.050 607.200 ;
        RECT 842.400 607.050 843.450 610.950 ;
        RECT 836.400 604.350 837.600 605.100 ;
        RECT 841.950 604.950 844.050 607.050 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 833.400 601.050 834.600 601.650 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 829.950 599.400 834.600 601.050 ;
        RECT 839.400 600.000 840.600 601.650 ;
        RECT 829.950 598.950 834.000 599.400 ;
        RECT 832.950 595.950 835.050 598.050 ;
        RECT 835.950 595.950 838.050 598.050 ;
        RECT 838.950 595.950 841.050 600.000 ;
        RECT 841.950 595.950 844.050 601.050 ;
        RECT 829.950 586.950 832.050 592.050 ;
        RECT 833.400 586.050 834.450 595.950 ;
        RECT 826.950 583.950 829.050 586.050 ;
        RECT 832.950 583.950 835.050 586.050 ;
        RECT 820.950 577.950 823.050 580.050 ;
        RECT 827.400 579.450 828.450 583.950 ;
        RECT 827.400 577.200 828.600 579.450 ;
        RECT 817.950 574.950 820.050 577.050 ;
        RECT 822.900 573.900 825.000 575.700 ;
        RECT 826.800 574.800 828.900 576.900 ;
        RECT 830.100 576.300 832.200 578.400 ;
        RECT 821.400 572.700 830.100 573.900 ;
        RECT 818.100 568.950 820.200 571.050 ;
        RECT 818.400 567.900 819.600 568.650 ;
        RECT 817.950 565.800 820.050 567.900 ;
        RECT 821.400 563.700 822.300 572.700 ;
        RECT 828.000 571.800 830.100 572.700 ;
        RECT 831.000 570.900 831.900 576.300 ;
        RECT 833.400 573.450 834.600 573.600 ;
        RECT 836.400 573.450 837.450 595.950 ;
        RECT 845.400 595.050 846.450 619.950 ;
        RECT 851.400 612.450 852.450 628.950 ;
        RECT 854.400 625.050 855.450 658.950 ;
        RECT 857.400 658.050 858.450 670.950 ;
        RECT 856.950 655.950 859.050 658.050 ;
        RECT 856.950 652.800 859.050 654.900 ;
        RECT 853.950 622.950 856.050 625.050 ;
        RECT 857.400 619.050 858.450 652.800 ;
        RECT 856.950 616.950 859.050 619.050 ;
        RECT 860.400 613.050 861.450 742.950 ;
        RECT 862.950 736.950 865.050 739.050 ;
        RECT 863.400 727.050 864.450 736.950 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 866.400 721.050 867.450 745.950 ;
        RECT 875.400 745.050 876.450 757.950 ;
        RECT 878.400 757.050 879.450 793.950 ;
        RECT 880.950 778.950 883.050 781.050 ;
        RECT 881.400 762.600 882.450 778.950 ;
        RECT 883.950 772.950 886.050 775.050 ;
        RECT 884.400 766.050 885.450 772.950 ;
        RECT 887.400 769.050 888.450 799.950 ;
        RECT 892.950 799.800 895.050 801.900 ;
        RECT 889.950 796.950 892.050 799.050 ;
        RECT 886.950 766.950 889.050 769.050 ;
        RECT 883.950 763.950 886.050 766.050 ;
        RECT 890.400 763.200 891.450 796.950 ;
        RECT 902.400 796.050 903.450 806.400 ;
        RECT 901.950 793.950 904.050 796.050 ;
        RECT 898.800 790.950 900.900 793.050 ;
        RECT 895.950 778.950 898.050 781.050 ;
        RECT 892.950 763.950 895.050 766.050 ;
        RECT 881.400 760.350 882.600 762.600 ;
        RECT 889.950 761.100 892.050 763.200 ;
        RECT 890.400 760.350 891.600 761.100 ;
        RECT 881.100 757.950 883.200 760.050 ;
        RECT 886.500 757.950 888.600 760.050 ;
        RECT 889.800 757.950 891.900 760.050 ;
        RECT 877.950 754.950 880.050 757.050 ;
        RECT 887.400 755.400 888.600 757.650 ;
        RECT 887.400 753.450 888.450 755.400 ;
        RECT 887.400 752.400 891.450 753.450 ;
        RECT 886.950 748.950 889.050 751.050 ;
        RECT 874.950 742.950 877.050 745.050 ;
        RECT 874.950 733.950 877.050 736.050 ;
        RECT 883.950 733.950 886.050 736.050 ;
        RECT 875.400 729.600 876.450 733.950 ;
        RECT 883.950 730.800 886.050 732.900 ;
        RECT 875.400 727.350 876.600 729.600 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 877.950 724.950 880.050 727.050 ;
        RECT 872.400 723.000 873.600 724.650 ;
        RECT 878.400 723.000 879.600 724.650 ;
        RECT 865.950 718.950 868.050 721.050 ;
        RECT 871.950 718.950 874.050 723.000 ;
        RECT 877.950 718.950 880.050 723.000 ;
        RECT 877.950 715.800 880.050 717.900 ;
        RECT 874.950 712.950 877.050 715.050 ;
        RECT 865.950 709.950 868.050 712.050 ;
        RECT 862.950 683.100 865.050 685.200 ;
        RECT 863.400 679.050 864.450 683.100 ;
        RECT 862.950 676.950 865.050 679.050 ;
        RECT 862.950 664.950 865.050 667.050 ;
        RECT 863.400 651.450 864.450 664.950 ;
        RECT 866.400 655.050 867.450 709.950 ;
        RECT 871.950 694.950 874.050 697.050 ;
        RECT 868.950 682.950 871.050 688.050 ;
        RECT 872.400 687.450 873.450 694.950 ;
        RECT 875.400 691.050 876.450 712.950 ;
        RECT 878.400 700.050 879.450 715.800 ;
        RECT 880.950 712.950 883.050 715.050 ;
        RECT 877.950 697.950 880.050 700.050 ;
        RECT 874.950 688.950 877.050 691.050 ;
        RECT 881.400 688.050 882.450 712.950 ;
        RECT 884.400 697.050 885.450 730.800 ;
        RECT 883.950 694.950 886.050 697.050 ;
        RECT 872.400 686.400 876.450 687.450 ;
        RECT 875.400 684.600 876.450 686.400 ;
        RECT 880.950 685.950 883.050 688.050 ;
        RECT 875.400 682.350 876.600 684.600 ;
        RECT 881.400 684.450 882.600 684.600 ;
        RECT 887.400 684.450 888.450 748.950 ;
        RECT 890.400 721.050 891.450 752.400 ;
        RECT 893.400 730.050 894.450 763.950 ;
        RECT 896.400 748.050 897.450 778.950 ;
        RECT 899.400 778.050 900.450 790.950 ;
        RECT 901.950 790.800 904.050 792.900 ;
        RECT 898.950 775.950 901.050 778.050 ;
        RECT 898.950 766.950 901.050 769.050 ;
        RECT 895.950 745.950 898.050 748.050 ;
        RECT 899.400 745.050 900.450 766.950 ;
        RECT 898.950 742.950 901.050 745.050 ;
        RECT 902.400 736.050 903.450 790.800 ;
        RECT 905.400 765.450 906.450 814.950 ;
        RECT 911.400 811.050 912.450 833.400 ;
        RECT 920.400 817.050 921.450 844.950 ;
        RECT 922.950 841.950 925.050 844.050 ;
        RECT 923.400 829.050 924.450 841.950 ;
        RECT 925.950 839.100 928.050 841.200 ;
        RECT 931.950 840.000 934.050 844.050 ;
        RECT 943.950 841.950 946.050 844.050 ;
        RECT 926.400 835.050 927.450 839.100 ;
        RECT 932.400 838.350 933.600 840.000 ;
        RECT 937.950 839.100 940.050 841.200 ;
        RECT 938.400 838.350 939.600 839.100 ;
        RECT 931.950 835.950 934.050 838.050 ;
        RECT 934.950 835.950 937.050 838.050 ;
        RECT 937.950 835.950 940.050 838.050 ;
        RECT 925.950 832.950 928.050 835.050 ;
        RECT 935.400 834.900 936.600 835.650 ;
        RECT 934.950 832.800 937.050 834.900 ;
        RECT 940.950 832.950 943.050 835.050 ;
        RECT 922.950 826.950 925.050 829.050 ;
        RECT 941.400 826.050 942.450 832.950 ;
        RECT 944.400 832.050 945.450 841.950 ;
        RECT 943.950 829.950 946.050 832.050 ;
        RECT 940.950 823.950 943.050 826.050 ;
        RECT 928.950 817.950 931.050 820.050 ;
        RECT 920.400 815.400 925.050 817.050 ;
        RECT 921.000 814.950 925.050 815.400 ;
        RECT 910.950 808.950 913.050 811.050 ;
        RECT 925.950 808.950 928.050 811.050 ;
        RECT 907.950 805.950 910.050 808.050 ;
        RECT 916.950 806.100 919.050 808.200 ;
        RECT 908.400 799.050 909.450 805.950 ;
        RECT 917.400 805.350 918.600 806.100 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 919.950 802.950 922.050 805.050 ;
        RECT 914.400 801.000 915.600 802.650 ;
        RECT 907.950 796.950 910.050 799.050 ;
        RECT 913.950 796.950 916.050 801.000 ;
        RECT 920.400 800.400 921.600 802.650 ;
        RECT 920.400 798.450 921.450 800.400 ;
        RECT 917.400 797.400 921.450 798.450 ;
        RECT 913.950 769.950 916.050 772.050 ;
        RECT 914.400 766.050 915.450 769.950 ;
        RECT 907.950 765.450 910.050 766.050 ;
        RECT 905.400 764.400 910.050 765.450 ;
        RECT 907.950 762.000 910.050 764.400 ;
        RECT 913.950 763.950 916.050 766.050 ;
        RECT 908.400 760.350 909.600 762.000 ;
        RECT 907.950 757.950 910.050 760.050 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 911.400 755.400 912.600 757.650 ;
        RECT 917.400 756.450 918.450 797.400 ;
        RECT 922.950 796.950 925.050 799.050 ;
        RECT 919.950 784.950 922.050 787.050 ;
        RECT 920.400 781.050 921.450 784.950 ;
        RECT 919.950 778.950 922.050 781.050 ;
        RECT 919.950 766.950 922.050 772.050 ;
        RECT 919.950 763.800 922.050 765.900 ;
        RECT 914.400 755.400 918.450 756.450 ;
        RECT 911.400 751.050 912.450 755.400 ;
        RECT 910.950 748.950 913.050 751.050 ;
        RECT 910.950 742.950 913.050 745.050 ;
        RECT 895.950 735.450 900.000 736.050 ;
        RECT 895.950 733.950 900.450 735.450 ;
        RECT 901.950 733.950 904.050 736.050 ;
        RECT 907.950 733.950 910.050 736.050 ;
        RECT 892.950 727.950 895.050 730.050 ;
        RECT 895.950 729.000 898.050 732.900 ;
        RECT 899.400 732.450 900.450 733.950 ;
        RECT 899.400 731.400 903.450 732.450 ;
        RECT 902.400 729.600 903.450 731.400 ;
        RECT 896.400 727.350 897.600 729.000 ;
        RECT 902.400 727.350 903.600 729.600 ;
        RECT 904.950 727.950 907.050 733.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 898.950 724.950 901.050 727.050 ;
        RECT 901.950 724.950 904.050 727.050 ;
        RECT 892.950 721.950 895.050 724.050 ;
        RECT 899.400 723.900 900.600 724.650 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 881.400 683.400 888.450 684.450 ;
        RECT 881.400 682.350 882.600 683.400 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 872.400 678.900 873.600 679.650 ;
        RECT 871.950 676.800 874.050 678.900 ;
        RECT 878.400 677.400 879.600 679.650 ;
        RECT 868.950 672.450 873.000 673.050 ;
        RECT 868.950 670.950 873.450 672.450 ;
        RECT 872.400 670.050 873.450 670.950 ;
        RECT 868.800 667.800 870.900 669.900 ;
        RECT 871.950 667.950 874.050 670.050 ;
        RECT 869.400 655.050 870.450 667.800 ;
        RECT 865.950 652.950 868.050 655.050 ;
        RECT 868.950 652.950 871.050 655.050 ;
        RECT 872.400 651.600 873.450 667.950 ;
        RECT 878.400 661.050 879.450 677.400 ;
        RECT 883.950 676.950 886.050 679.050 ;
        RECT 884.400 664.050 885.450 676.950 ;
        RECT 883.950 661.950 886.050 664.050 ;
        RECT 877.950 658.950 880.050 661.050 ;
        RECT 887.400 658.050 888.450 683.400 ;
        RECT 890.400 676.050 891.450 718.950 ;
        RECT 889.950 673.950 892.050 676.050 ;
        RECT 893.400 664.050 894.450 721.950 ;
        RECT 898.950 721.800 901.050 723.900 ;
        RECT 901.950 718.950 904.050 721.050 ;
        RECT 902.400 703.050 903.450 718.950 ;
        RECT 908.400 712.050 909.450 733.950 ;
        RECT 911.400 715.050 912.450 742.950 ;
        RECT 910.950 712.950 913.050 715.050 ;
        RECT 907.950 709.950 910.050 712.050 ;
        RECT 907.950 706.800 910.050 708.900 ;
        RECT 908.400 703.050 909.450 706.800 ;
        RECT 910.950 703.950 913.050 706.050 ;
        RECT 901.950 700.950 904.050 703.050 ;
        RECT 907.950 700.950 910.050 703.050 ;
        RECT 895.950 697.950 898.050 700.050 ;
        RECT 896.400 691.050 897.450 697.950 ;
        RECT 911.400 691.050 912.450 703.950 ;
        RECT 895.950 688.950 898.050 691.050 ;
        RECT 907.800 690.000 909.900 691.050 ;
        RECT 907.800 688.950 910.050 690.000 ;
        RECT 910.950 688.950 913.050 691.050 ;
        RECT 907.950 685.950 910.050 688.950 ;
        RECT 914.400 688.050 915.450 755.400 ;
        RECT 920.400 753.450 921.450 763.800 ;
        RECT 923.400 756.450 924.450 796.950 ;
        RECT 926.400 763.050 927.450 808.950 ;
        RECT 929.400 790.050 930.450 817.950 ;
        RECT 943.950 814.950 946.050 817.050 ;
        RECT 937.950 806.100 940.050 808.200 ;
        RECT 944.400 807.600 945.450 814.950 ;
        RECT 947.400 811.050 948.450 853.950 ;
        RECT 946.950 808.950 949.050 811.050 ;
        RECT 938.400 805.350 939.600 806.100 ;
        RECT 944.400 805.350 945.600 807.600 ;
        RECT 934.950 802.950 937.050 805.050 ;
        RECT 937.950 802.950 940.050 805.050 ;
        RECT 940.950 802.950 943.050 805.050 ;
        RECT 943.950 802.950 946.050 805.050 ;
        RECT 935.400 801.900 936.600 802.650 ;
        RECT 934.950 799.800 937.050 801.900 ;
        RECT 941.400 801.000 942.600 802.650 ;
        RECT 940.950 796.950 943.050 801.000 ;
        RECT 946.950 799.950 949.050 802.050 ;
        RECT 943.950 793.950 946.050 796.050 ;
        RECT 928.950 787.950 931.050 790.050 ;
        RECT 929.400 766.050 930.450 787.950 ;
        RECT 944.400 784.050 945.450 793.950 ;
        RECT 943.950 781.950 946.050 784.050 ;
        RECT 937.950 775.950 940.050 778.050 ;
        RECT 931.950 769.950 934.050 772.050 ;
        RECT 928.950 763.950 931.050 766.050 ;
        RECT 925.950 760.950 928.050 763.050 ;
        RECT 932.400 762.600 933.450 769.950 ;
        RECT 938.400 769.050 939.450 775.950 ;
        RECT 943.950 772.950 946.050 775.050 ;
        RECT 937.950 766.950 940.050 769.050 ;
        RECT 938.400 762.600 939.450 766.950 ;
        RECT 932.400 760.350 933.600 762.600 ;
        RECT 938.400 760.350 939.600 762.600 ;
        RECT 928.950 757.950 931.050 760.050 ;
        RECT 931.950 757.950 934.050 760.050 ;
        RECT 934.950 757.950 937.050 760.050 ;
        RECT 937.950 757.950 940.050 760.050 ;
        RECT 923.400 755.400 927.450 756.450 ;
        RECT 917.400 752.400 921.450 753.450 ;
        RECT 917.400 730.050 918.450 752.400 ;
        RECT 926.400 751.050 927.450 755.400 ;
        RECT 929.400 755.400 930.600 757.650 ;
        RECT 935.400 755.400 936.600 757.650 ;
        RECT 919.950 748.950 922.050 751.050 ;
        RECT 925.950 748.950 928.050 751.050 ;
        RECT 920.400 733.050 921.450 748.950 ;
        RECT 929.400 748.050 930.450 755.400 ;
        RECT 931.950 748.950 934.050 751.050 ;
        RECT 928.950 745.950 931.050 748.050 ;
        RECT 925.950 742.950 928.050 745.050 ;
        RECT 926.400 739.050 927.450 742.950 ;
        RECT 925.950 736.950 928.050 739.050 ;
        RECT 916.950 727.950 919.050 730.050 ;
        RECT 919.950 729.000 922.050 733.050 ;
        RECT 926.400 729.600 927.450 736.950 ;
        RECT 920.400 727.350 921.600 729.000 ;
        RECT 926.400 727.350 927.600 729.600 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 922.950 724.950 925.050 727.050 ;
        RECT 925.950 724.950 928.050 727.050 ;
        RECT 923.400 722.400 924.600 724.650 ;
        RECT 923.400 721.050 924.450 722.400 ;
        RECT 919.950 718.950 922.050 721.050 ;
        RECT 923.400 719.400 928.050 721.050 ;
        RECT 924.000 718.950 928.050 719.400 ;
        RECT 928.950 718.950 931.050 724.050 ;
        RECT 916.950 715.950 919.050 718.050 ;
        RECT 917.400 706.050 918.450 715.950 ;
        RECT 928.950 715.800 931.050 717.900 ;
        RECT 919.950 712.950 922.050 715.050 ;
        RECT 916.950 703.950 919.050 706.050 ;
        RECT 913.950 685.950 916.050 688.050 ;
        RECT 898.950 683.100 901.050 685.200 ;
        RECT 904.950 683.100 907.050 685.200 ;
        RECT 899.400 682.350 900.600 683.100 ;
        RECT 905.400 682.350 906.600 683.100 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 902.400 678.000 903.600 679.650 ;
        RECT 908.400 679.050 909.600 679.650 ;
        RECT 908.400 678.900 913.050 679.050 ;
        RECT 901.950 676.050 904.050 678.000 ;
        RECT 907.950 676.950 913.050 678.900 ;
        RECT 907.950 676.800 910.050 676.950 ;
        RECT 914.400 676.050 915.450 685.950 ;
        RECT 916.950 679.950 919.050 682.050 ;
        RECT 901.800 675.000 904.050 676.050 ;
        RECT 901.800 673.950 903.900 675.000 ;
        RECT 904.950 673.950 907.050 676.050 ;
        RECT 913.950 673.950 916.050 676.050 ;
        RECT 893.400 661.950 898.050 664.050 ;
        RECT 880.950 655.950 883.050 658.050 ;
        RECT 886.950 655.950 889.050 658.050 ;
        RECT 866.400 651.450 867.600 651.600 ;
        RECT 863.400 650.400 867.600 651.450 ;
        RECT 866.400 649.350 867.600 650.400 ;
        RECT 872.400 649.350 873.600 651.600 ;
        RECT 881.400 649.050 882.450 655.950 ;
        RECT 893.400 655.050 894.450 661.950 ;
        RECT 886.950 652.800 889.050 654.900 ;
        RECT 892.950 652.950 895.050 655.050 ;
        RECT 883.950 649.950 886.050 652.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 874.950 646.950 877.050 649.050 ;
        RECT 880.950 646.950 883.050 649.050 ;
        RECT 869.400 645.000 870.600 646.650 ;
        RECT 875.400 645.450 876.600 646.650 ;
        RECT 868.950 640.950 871.050 645.000 ;
        RECT 875.400 644.400 879.450 645.450 ;
        RECT 862.950 634.950 865.050 637.050 ;
        RECT 863.400 619.050 864.450 634.950 ;
        RECT 878.400 634.050 879.450 644.400 ;
        RECT 877.950 631.950 880.050 634.050 ;
        RECT 874.950 625.950 877.050 628.050 ;
        RECT 862.950 616.950 865.050 619.050 ;
        RECT 848.400 611.400 852.450 612.450 ;
        RECT 844.950 592.950 847.050 595.050 ;
        RECT 844.950 589.800 847.050 591.900 ;
        RECT 841.950 580.950 844.050 583.050 ;
        RECT 833.400 572.400 837.450 573.450 ;
        RECT 833.400 571.350 834.600 572.400 ;
        RECT 825.000 569.700 831.900 570.900 ;
        RECT 825.000 567.300 825.900 569.700 ;
        RECT 823.800 565.200 825.900 567.300 ;
        RECT 826.800 565.950 828.900 568.050 ;
        RECT 814.950 559.950 817.050 562.050 ;
        RECT 820.500 561.600 822.600 563.700 ;
        RECT 827.400 563.400 828.600 565.650 ;
        RECT 830.700 562.500 831.900 569.700 ;
        RECT 832.800 568.950 834.900 571.050 ;
        RECT 830.100 560.400 832.200 562.500 ;
        RECT 836.400 559.050 837.450 572.400 ;
        RECT 838.950 571.950 841.050 574.050 ;
        RECT 832.800 556.950 834.900 559.050 ;
        RECT 835.950 556.950 838.050 559.050 ;
        RECT 833.400 547.050 834.450 556.950 ;
        RECT 832.950 544.950 835.050 547.050 ;
        RECT 835.950 538.950 838.050 541.050 ;
        RECT 811.950 535.950 814.050 538.050 ;
        RECT 829.950 535.950 832.050 538.050 ;
        RECT 811.950 526.950 814.050 529.050 ;
        RECT 823.950 528.000 826.050 532.050 ;
        RECT 830.400 528.600 831.450 535.950 ;
        RECT 832.950 532.950 835.050 535.050 ;
        RECT 833.400 529.050 834.450 532.950 ;
        RECT 836.400 532.050 837.450 538.950 ;
        RECT 835.950 529.950 838.050 532.050 ;
        RECT 796.950 517.950 799.050 522.000 ;
        RECT 802.950 520.800 805.050 522.900 ;
        RECT 808.950 520.950 811.050 523.050 ;
        RECT 808.950 514.950 811.050 517.050 ;
        RECT 799.950 511.950 802.050 514.050 ;
        RECT 790.950 508.950 793.050 511.050 ;
        RECT 767.700 501.300 769.800 503.400 ;
        RECT 770.700 501.300 772.800 503.400 ;
        RECT 773.700 501.300 775.800 503.400 ;
        RECT 763.950 496.950 766.050 499.050 ;
        RECT 768.300 497.700 769.500 501.300 ;
        RECT 746.100 490.950 748.200 493.050 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 764.400 492.900 765.450 496.950 ;
        RECT 767.400 495.600 769.500 497.700 ;
        RECT 763.950 490.800 766.050 492.900 ;
        RECT 754.800 487.950 756.900 490.050 ;
        RECT 760.800 487.950 762.900 490.050 ;
        RECT 755.400 485.400 756.600 487.650 ;
        RECT 755.400 469.050 756.450 485.400 ;
        RECT 757.950 484.950 760.050 487.050 ;
        RECT 763.950 484.950 766.050 487.050 ;
        RECT 758.400 475.050 759.450 484.950 ;
        RECT 757.950 472.950 760.050 475.050 ;
        RECT 754.950 466.950 757.050 469.050 ;
        RECT 764.400 466.050 765.450 484.950 ;
        RECT 767.400 476.700 768.900 495.600 ;
        RECT 771.300 484.800 772.500 501.300 ;
        RECT 770.400 482.700 772.500 484.800 ;
        RECT 771.300 476.700 772.500 482.700 ;
        RECT 773.700 479.700 774.900 501.300 ;
        RECT 781.800 500.400 783.900 502.500 ;
        RECT 787.200 501.300 789.300 503.400 ;
        RECT 790.200 501.300 792.300 503.400 ;
        RECT 793.200 501.300 795.300 503.400 ;
        RECT 778.800 493.950 780.900 496.050 ;
        RECT 779.400 492.900 780.600 493.650 ;
        RECT 778.950 490.800 781.050 492.900 ;
        RECT 782.400 489.900 783.300 500.400 ;
        RECT 785.100 494.400 787.200 496.500 ;
        RECT 782.400 487.800 784.500 489.900 ;
        RECT 788.100 489.000 789.300 501.300 ;
        RECT 778.950 481.950 781.050 484.050 ;
        RECT 773.700 477.600 775.800 479.700 ;
        RECT 767.400 474.600 770.400 476.700 ;
        RECT 771.300 474.600 773.400 476.700 ;
        RECT 779.400 472.050 780.450 481.950 ;
        RECT 782.400 481.200 783.300 487.800 ;
        RECT 787.800 486.900 789.900 489.000 ;
        RECT 782.400 479.100 784.500 481.200 ;
        RECT 788.100 479.700 789.300 486.900 ;
        RECT 790.800 483.600 792.300 501.300 ;
        RECT 790.800 481.500 792.900 483.600 ;
        RECT 787.800 477.600 789.900 479.700 ;
        RECT 790.800 476.700 792.300 481.500 ;
        RECT 794.100 479.700 795.300 501.300 ;
        RECT 790.200 474.600 792.300 476.700 ;
        RECT 793.200 474.600 795.300 479.700 ;
        RECT 796.200 501.300 798.300 503.400 ;
        RECT 796.200 483.600 797.700 501.300 ;
        RECT 800.400 487.050 801.450 511.950 ;
        RECT 809.400 511.050 810.450 514.950 ;
        RECT 808.950 508.950 811.050 511.050 ;
        RECT 805.950 491.100 808.050 493.200 ;
        RECT 806.400 490.350 807.600 491.100 ;
        RECT 805.800 487.950 807.900 490.050 ;
        RECT 799.950 484.950 802.050 487.050 ;
        RECT 809.400 484.050 810.450 508.950 ;
        RECT 812.400 505.050 813.450 526.950 ;
        RECT 824.400 526.350 825.600 528.000 ;
        RECT 830.400 526.350 831.600 528.600 ;
        RECT 832.800 526.950 834.900 529.050 ;
        RECT 835.950 526.800 838.050 528.900 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 826.950 523.950 829.050 526.050 ;
        RECT 829.950 523.950 832.050 526.050 ;
        RECT 811.950 502.950 814.050 505.050 ;
        RECT 811.950 496.950 814.050 499.050 ;
        RECT 812.400 492.450 813.450 496.950 ;
        RECT 815.400 496.050 816.450 523.950 ;
        RECT 817.950 520.950 820.050 523.050 ;
        RECT 821.400 522.000 822.600 523.650 ;
        RECT 827.400 522.900 828.600 523.650 ;
        RECT 818.400 496.050 819.450 520.950 ;
        RECT 820.950 517.950 823.050 522.000 ;
        RECT 826.950 520.800 829.050 522.900 ;
        RECT 832.950 520.950 835.050 523.050 ;
        RECT 829.950 517.950 832.050 520.050 ;
        RECT 830.400 513.450 831.450 517.950 ;
        RECT 833.400 517.050 834.450 520.950 ;
        RECT 832.950 514.950 835.050 517.050 ;
        RECT 830.400 512.400 834.450 513.450 ;
        RECT 823.950 505.950 826.050 508.050 ;
        RECT 820.950 496.950 823.050 499.050 ;
        RECT 814.950 493.950 817.050 496.050 ;
        RECT 817.800 493.950 819.900 496.050 ;
        RECT 820.950 493.800 823.050 495.900 ;
        RECT 815.400 492.450 816.600 492.600 ;
        RECT 812.400 491.400 816.600 492.450 ;
        RECT 815.400 490.350 816.600 491.400 ;
        RECT 817.950 490.800 820.050 492.900 ;
        RECT 814.800 487.950 816.900 490.050 ;
        RECT 796.200 481.500 798.300 483.600 ;
        RECT 799.950 481.800 802.050 483.900 ;
        RECT 808.800 481.950 810.900 484.050 ;
        RECT 811.950 481.950 814.050 484.050 ;
        RECT 796.200 476.700 797.700 481.500 ;
        RECT 796.200 474.600 798.300 476.700 ;
        RECT 778.950 469.950 781.050 472.050 ;
        RECT 784.950 466.950 787.050 469.050 ;
        RECT 743.700 462.300 745.800 464.400 ;
        RECT 744.300 457.500 745.800 462.300 ;
        RECT 743.700 455.400 745.800 457.500 ;
        RECT 739.950 439.950 742.050 442.050 ;
        RECT 744.300 437.700 745.800 455.400 ;
        RECT 743.700 435.600 745.800 437.700 ;
        RECT 746.700 459.300 748.800 464.400 ;
        RECT 749.700 462.300 751.800 464.400 ;
        RECT 763.950 463.950 766.050 466.050 ;
        RECT 768.600 462.300 770.700 464.400 ;
        RECT 771.600 462.300 774.600 464.400 ;
        RECT 775.950 463.950 778.050 466.050 ;
        RECT 746.700 437.700 747.900 459.300 ;
        RECT 749.700 457.500 751.200 462.300 ;
        RECT 752.100 459.300 754.200 461.400 ;
        RECT 749.100 455.400 751.200 457.500 ;
        RECT 749.700 437.700 751.200 455.400 ;
        RECT 752.700 452.100 753.900 459.300 ;
        RECT 757.500 457.800 759.600 459.900 ;
        RECT 766.200 459.300 768.300 461.400 ;
        RECT 752.100 450.000 754.200 452.100 ;
        RECT 758.700 451.200 759.600 457.800 ;
        RECT 752.700 437.700 753.900 450.000 ;
        RECT 757.500 449.100 759.600 451.200 ;
        RECT 754.800 442.500 756.900 444.600 ;
        RECT 758.700 438.600 759.600 449.100 ;
        RECT 760.950 446.100 763.050 448.200 ;
        RECT 761.400 445.350 762.600 446.100 ;
        RECT 761.100 442.950 763.200 445.050 ;
        RECT 746.700 435.600 748.800 437.700 ;
        RECT 749.700 435.600 751.800 437.700 ;
        RECT 752.700 435.600 754.800 437.700 ;
        RECT 758.100 436.500 760.200 438.600 ;
        RECT 767.100 437.700 768.300 459.300 ;
        RECT 769.500 456.300 770.700 462.300 ;
        RECT 769.500 454.200 771.600 456.300 ;
        RECT 769.500 437.700 770.700 454.200 ;
        RECT 773.100 443.400 774.600 462.300 ;
        RECT 772.500 441.300 774.600 443.400 ;
        RECT 772.500 437.700 773.700 441.300 ;
        RECT 766.200 435.600 768.300 437.700 ;
        RECT 769.200 435.600 771.300 437.700 ;
        RECT 772.200 435.600 774.300 437.700 ;
        RECT 763.950 430.950 766.050 433.050 ;
        RECT 751.950 427.950 754.050 430.050 ;
        RECT 752.400 417.600 753.450 427.950 ;
        RECT 764.400 424.050 765.450 430.950 ;
        RECT 776.400 427.050 777.450 463.950 ;
        RECT 785.400 463.050 786.450 466.950 ;
        RECT 793.950 463.950 796.050 466.050 ;
        RECT 784.950 460.950 787.050 463.050 ;
        RECT 785.400 453.600 786.450 460.950 ;
        RECT 785.400 451.350 786.600 453.600 ;
        RECT 779.100 448.950 781.200 451.050 ;
        RECT 785.100 448.950 787.200 451.050 ;
        RECT 784.950 442.950 787.050 445.050 ;
        RECT 781.950 439.950 784.050 442.050 ;
        RECT 766.950 424.950 769.050 427.050 ;
        RECT 775.950 424.950 778.050 427.050 ;
        RECT 763.950 421.950 766.050 424.050 ;
        RECT 752.400 415.350 753.600 417.600 ;
        RECT 757.950 416.100 760.050 421.050 ;
        RECT 767.400 420.450 768.450 424.950 ;
        RECT 764.400 419.400 768.450 420.450 ;
        RECT 758.400 415.350 759.600 416.100 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 757.950 412.950 760.050 415.050 ;
        RECT 748.950 409.950 751.050 412.050 ;
        RECT 755.400 410.400 756.600 412.650 ;
        RECT 764.400 411.900 765.450 419.400 ;
        RECT 769.950 418.950 772.050 421.050 ;
        RECT 766.950 415.950 769.050 418.050 ;
        RECT 718.950 397.950 721.050 400.050 ;
        RECT 736.950 397.950 739.050 400.050 ;
        RECT 719.400 361.050 720.450 397.950 ;
        RECT 739.950 394.950 742.050 397.050 ;
        RECT 727.950 388.950 730.050 391.050 ;
        RECT 721.950 376.950 724.050 379.050 ;
        RECT 718.950 358.950 721.050 361.050 ;
        RECT 722.400 349.050 723.450 376.950 ;
        RECT 728.400 373.050 729.450 388.950 ;
        RECT 724.950 370.950 727.050 373.050 ;
        RECT 727.950 370.950 730.050 373.050 ;
        RECT 733.950 371.100 736.050 373.200 ;
        RECT 740.400 373.050 741.450 394.950 ;
        RECT 749.400 394.050 750.450 409.950 ;
        RECT 748.950 391.950 751.050 394.050 ;
        RECT 745.950 379.950 748.050 382.050 ;
        RECT 725.400 361.050 726.450 370.950 ;
        RECT 734.400 370.350 735.600 371.100 ;
        RECT 739.950 370.950 742.050 373.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 731.400 366.900 732.600 367.650 ;
        RECT 730.950 364.800 733.050 366.900 ;
        RECT 737.400 365.400 738.600 367.650 ;
        RECT 724.950 358.950 727.050 361.050 ;
        RECT 730.950 360.450 735.000 361.050 ;
        RECT 730.950 358.950 735.450 360.450 ;
        RECT 727.950 355.950 730.050 358.050 ;
        RECT 734.400 352.050 735.450 358.950 ;
        RECT 737.400 358.050 738.450 365.400 ;
        RECT 739.950 364.950 742.050 367.050 ;
        RECT 736.950 355.950 739.050 358.050 ;
        RECT 733.950 349.950 736.050 352.050 ;
        RECT 706.950 345.000 709.050 349.050 ;
        RECT 715.950 346.950 718.050 349.050 ;
        RECT 721.950 346.950 724.050 349.050 ;
        RECT 724.950 346.950 727.050 349.050 ;
        RECT 730.950 346.950 733.050 349.050 ;
        RECT 707.400 343.200 708.600 345.000 ;
        RECT 703.500 341.100 705.600 343.200 ;
        RECT 701.400 339.450 702.600 339.600 ;
        RECT 698.400 338.400 702.600 339.450 ;
        RECT 701.400 337.350 702.600 338.400 ;
        RECT 701.100 334.950 703.200 337.050 ;
        RECT 704.100 336.000 705.000 341.100 ;
        RECT 706.800 340.800 708.900 342.900 ;
        RECT 713.400 341.400 715.500 343.500 ;
        RECT 711.000 339.000 713.100 339.900 ;
        RECT 705.900 337.800 713.100 339.000 ;
        RECT 705.900 336.900 708.000 337.800 ;
        RECT 711.000 336.000 713.100 336.900 ;
        RECT 704.100 335.100 713.100 336.000 ;
        RECT 704.100 328.500 705.000 335.100 ;
        RECT 711.000 334.800 713.100 335.100 ;
        RECT 706.800 331.950 708.900 334.050 ;
        RECT 707.400 329.400 708.600 331.650 ;
        RECT 714.000 328.800 714.900 341.400 ;
        RECT 718.950 340.950 721.050 343.050 ;
        RECT 715.800 334.950 717.900 337.050 ;
        RECT 716.400 333.450 717.600 334.650 ;
        RECT 716.400 333.000 720.450 333.450 ;
        RECT 716.400 332.400 721.050 333.000 ;
        RECT 718.950 328.950 721.050 332.400 ;
        RECT 704.100 326.400 706.200 328.500 ;
        RECT 709.950 325.950 712.050 328.050 ;
        RECT 713.100 326.700 715.200 328.800 ;
        RECT 694.950 310.950 697.050 313.050 ;
        RECT 691.950 298.950 694.050 301.050 ;
        RECT 683.400 296.400 687.450 297.450 ;
        RECT 683.400 294.600 684.450 296.400 ;
        RECT 688.950 296.100 691.050 298.200 ;
        RECT 710.400 298.050 711.450 325.950 ;
        RECT 697.950 295.950 700.050 298.050 ;
        RECT 703.950 295.950 706.050 298.050 ;
        RECT 709.950 295.950 712.050 298.050 ;
        RECT 683.400 292.350 684.600 294.600 ;
        RECT 688.950 292.950 691.050 295.050 ;
        RECT 689.400 292.350 690.600 292.950 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 686.400 287.400 687.600 289.650 ;
        RECT 692.400 287.400 693.600 289.650 ;
        RECT 686.400 283.050 687.450 287.400 ;
        RECT 685.950 280.950 688.050 283.050 ;
        RECT 692.400 280.050 693.450 287.400 ;
        RECT 691.950 277.950 694.050 280.050 ;
        RECT 685.950 274.950 688.050 277.050 ;
        RECT 676.950 265.950 679.050 268.050 ;
        RECT 682.950 265.950 685.050 268.050 ;
        RECT 674.400 260.400 678.450 261.450 ;
        RECT 662.400 259.350 663.600 260.100 ;
        RECT 668.400 259.350 669.600 260.100 ;
        RECT 661.950 256.950 664.050 259.050 ;
        RECT 664.950 256.950 667.050 259.050 ;
        RECT 667.950 256.950 670.050 259.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 677.400 258.600 678.450 260.400 ;
        RECT 665.400 255.900 666.600 256.650 ;
        RECT 655.950 253.800 658.050 255.900 ;
        RECT 664.950 253.800 667.050 255.900 ;
        RECT 671.400 254.400 672.600 256.650 ;
        RECT 677.400 256.350 678.600 258.600 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 646.950 226.950 649.050 229.050 ;
        RECT 634.950 223.950 637.050 226.050 ;
        RECT 629.400 214.350 630.600 216.600 ;
        RECT 634.950 215.100 637.050 217.200 ;
        RECT 643.950 215.100 646.050 217.200 ;
        RECT 635.400 214.350 636.600 215.100 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 632.400 210.900 633.600 211.650 ;
        RECT 631.950 208.800 634.050 210.900 ;
        RECT 638.400 209.400 639.600 211.650 ;
        RECT 638.400 196.050 639.450 209.400 ;
        RECT 634.800 193.950 636.900 196.050 ;
        RECT 637.950 193.950 640.050 196.050 ;
        RECT 628.950 182.100 631.050 184.200 ;
        RECT 635.400 183.600 636.450 193.950 ;
        RECT 644.400 190.050 645.450 215.100 ;
        RECT 643.950 187.950 646.050 190.050 ;
        RECT 629.400 178.050 630.450 182.100 ;
        RECT 635.400 181.350 636.600 183.600 ;
        RECT 640.950 182.100 643.050 184.200 ;
        RECT 647.400 183.450 648.450 226.950 ;
        RECT 650.400 196.050 651.450 241.950 ;
        RECT 655.950 229.950 658.050 232.050 ;
        RECT 656.400 216.600 657.450 229.950 ;
        RECT 671.400 223.050 672.450 254.400 ;
        RECT 673.950 253.950 676.050 256.050 ;
        RECT 677.100 253.950 679.200 256.050 ;
        RECT 670.950 220.950 673.050 223.050 ;
        RECT 656.400 214.350 657.600 216.600 ;
        RECT 661.950 215.100 664.050 217.200 ;
        RECT 667.950 215.100 670.050 217.200 ;
        RECT 662.400 214.350 663.600 215.100 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 659.400 210.900 660.600 211.650 ;
        RECT 658.950 208.800 661.050 210.900 ;
        RECT 668.400 202.050 669.450 215.100 ;
        RECT 667.950 199.950 670.050 202.050 ;
        RECT 649.950 193.950 652.050 196.050 ;
        RECT 664.950 193.950 667.050 196.050 ;
        RECT 665.400 183.600 666.450 193.950 ;
        RECT 647.400 182.400 651.450 183.450 ;
        RECT 641.400 181.350 642.600 182.100 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 628.950 175.950 631.050 178.050 ;
        RECT 638.400 177.000 639.600 178.650 ;
        RECT 637.950 172.950 640.050 177.000 ;
        RECT 644.400 176.400 645.600 178.650 ;
        RECT 650.400 177.900 651.450 182.400 ;
        RECT 665.400 181.350 666.600 183.600 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 662.400 177.900 663.600 178.650 ;
        RECT 644.400 172.050 645.450 176.400 ;
        RECT 649.950 175.800 652.050 177.900 ;
        RECT 661.950 175.800 664.050 177.900 ;
        RECT 643.950 169.950 646.050 172.050 ;
        RECT 644.400 157.050 645.450 169.950 ;
        RECT 655.950 163.950 658.050 166.050 ;
        RECT 631.950 154.950 634.050 157.050 ;
        RECT 643.950 154.950 646.050 157.050 ;
        RECT 632.400 151.050 633.450 154.950 ;
        RECT 631.950 148.950 634.050 151.050 ;
        RECT 628.950 145.950 631.050 148.050 ;
        RECT 628.950 142.800 631.050 144.900 ;
        RECT 614.400 136.350 615.600 138.600 ;
        RECT 620.400 136.350 621.600 138.600 ;
        RECT 622.950 137.100 625.050 139.200 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 611.400 131.400 612.600 133.650 ;
        RECT 617.400 132.000 618.600 133.650 ;
        RECT 611.400 112.050 612.450 131.400 ;
        RECT 616.950 127.950 619.050 132.000 ;
        RECT 629.400 130.050 630.450 142.800 ;
        RECT 628.950 127.950 631.050 130.050 ;
        RECT 632.400 112.050 633.450 148.950 ;
        RECT 634.950 145.950 637.050 148.050 ;
        RECT 640.500 141.300 642.600 143.400 ;
        RECT 650.100 142.500 652.200 144.600 ;
        RECT 637.950 137.100 640.050 139.200 ;
        RECT 638.400 136.350 639.600 137.100 ;
        RECT 638.100 133.950 640.200 136.050 ;
        RECT 634.950 130.800 637.050 132.900 ;
        RECT 641.400 132.300 642.300 141.300 ;
        RECT 643.800 137.700 645.900 139.800 ;
        RECT 647.400 139.350 648.600 141.600 ;
        RECT 645.000 135.300 645.900 137.700 ;
        RECT 646.800 136.950 648.900 139.050 ;
        RECT 650.700 135.300 651.900 142.500 ;
        RECT 645.000 134.100 651.900 135.300 ;
        RECT 648.000 132.300 650.100 133.200 ;
        RECT 641.400 131.100 650.100 132.300 ;
        RECT 635.400 118.050 636.450 130.800 ;
        RECT 642.900 129.300 645.000 131.100 ;
        RECT 646.800 128.100 648.900 130.200 ;
        RECT 651.000 128.700 651.900 134.100 ;
        RECT 652.800 133.950 654.900 136.050 ;
        RECT 653.400 132.900 654.600 133.650 ;
        RECT 652.950 130.800 655.050 132.900 ;
        RECT 647.400 125.550 648.600 127.800 ;
        RECT 650.100 126.600 652.200 128.700 ;
        RECT 634.950 115.950 637.050 118.050 ;
        RECT 647.400 115.050 648.450 125.550 ;
        RECT 646.950 112.950 649.050 115.050 ;
        RECT 610.950 109.950 613.050 112.050 ;
        RECT 625.950 109.950 628.050 112.050 ;
        RECT 631.950 109.950 634.050 112.050 ;
        RECT 604.950 103.950 607.050 106.050 ;
        RECT 616.950 104.100 619.050 106.200 ;
        RECT 601.950 94.950 604.050 97.050 ;
        RECT 605.400 94.050 606.450 103.950 ;
        RECT 617.400 103.350 618.600 104.100 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 614.400 99.000 615.600 100.650 ;
        RECT 620.400 99.900 621.600 100.650 ;
        RECT 626.400 99.900 627.450 109.950 ;
        RECT 646.950 109.800 649.050 111.900 ;
        RECT 647.400 109.200 648.600 109.800 ;
        RECT 642.900 105.900 645.000 107.700 ;
        RECT 646.800 106.800 648.900 108.900 ;
        RECT 650.100 108.300 652.200 110.400 ;
        RECT 641.400 104.700 650.100 105.900 ;
        RECT 638.100 100.950 640.200 103.050 ;
        RECT 638.400 99.900 639.600 100.650 ;
        RECT 613.950 94.950 616.050 99.000 ;
        RECT 619.950 97.800 622.050 99.900 ;
        RECT 625.950 97.800 628.050 99.900 ;
        RECT 631.950 97.800 634.050 99.900 ;
        RECT 637.950 97.800 640.050 99.900 ;
        RECT 604.950 91.950 607.050 94.050 ;
        RECT 616.950 85.950 619.050 88.050 ;
        RECT 595.950 82.950 598.050 85.050 ;
        RECT 580.950 79.950 583.050 82.050 ;
        RECT 607.950 67.950 610.050 70.050 ;
        RECT 550.800 64.200 552.900 66.300 ;
        RECT 559.800 64.500 561.900 66.600 ;
        RECT 577.950 64.950 580.050 67.050 ;
        RECT 547.950 59.100 550.050 61.200 ;
        RECT 548.400 58.350 549.600 59.100 ;
        RECT 548.100 55.950 550.200 58.050 ;
        RECT 544.950 52.800 547.050 54.900 ;
        RECT 551.100 51.600 552.000 64.200 ;
        RECT 557.400 61.350 558.600 63.600 ;
        RECT 557.100 58.950 559.200 61.050 ;
        RECT 552.900 57.900 555.000 58.200 ;
        RECT 561.000 57.900 561.900 64.500 ;
        RECT 568.950 59.100 571.050 61.200 ;
        RECT 552.900 57.000 561.900 57.900 ;
        RECT 552.900 56.100 555.000 57.000 ;
        RECT 558.000 55.200 560.100 56.100 ;
        RECT 552.900 54.000 560.100 55.200 ;
        RECT 552.900 53.100 555.000 54.000 ;
        RECT 550.500 49.500 552.600 51.600 ;
        RECT 557.100 50.100 559.200 52.200 ;
        RECT 561.000 51.900 561.900 57.000 ;
        RECT 562.800 55.950 564.900 58.050 ;
        RECT 563.400 54.450 564.600 55.650 ;
        RECT 563.400 53.400 567.450 54.450 ;
        RECT 560.400 49.800 562.500 51.900 ;
        RECT 557.400 48.000 558.600 49.800 ;
        RECT 566.400 49.050 567.450 53.400 ;
        RECT 556.950 43.950 559.050 48.000 ;
        RECT 565.950 46.950 568.050 49.050 ;
        RECT 547.950 26.100 550.050 28.200 ;
        RECT 553.950 26.100 556.050 28.200 ;
        RECT 569.400 28.050 570.450 59.100 ;
        RECT 578.400 54.450 579.450 64.950 ;
        RECT 583.800 64.500 585.900 66.600 ;
        RECT 581.100 55.950 583.200 58.050 ;
        RECT 584.100 57.300 585.300 64.500 ;
        RECT 587.400 61.350 588.600 63.600 ;
        RECT 593.400 63.300 595.500 65.400 ;
        RECT 587.100 58.950 589.200 61.050 ;
        RECT 590.100 59.700 592.200 61.800 ;
        RECT 590.100 57.300 591.000 59.700 ;
        RECT 584.100 56.100 591.000 57.300 ;
        RECT 581.400 54.450 582.600 55.650 ;
        RECT 578.400 53.400 582.600 54.450 ;
        RECT 584.100 50.700 585.000 56.100 ;
        RECT 585.900 54.300 588.000 55.200 ;
        RECT 593.700 54.300 594.600 63.300 ;
        RECT 595.950 59.100 598.050 61.200 ;
        RECT 604.950 59.100 607.050 61.200 ;
        RECT 596.400 58.350 597.600 59.100 ;
        RECT 595.800 55.950 597.900 58.050 ;
        RECT 585.900 53.100 594.600 54.300 ;
        RECT 583.800 48.600 585.900 50.700 ;
        RECT 587.100 50.100 589.200 52.200 ;
        RECT 591.000 51.300 593.100 53.100 ;
        RECT 587.400 49.050 588.600 49.800 ;
        RECT 586.950 46.950 589.050 49.050 ;
        RECT 577.950 43.950 580.050 46.050 ;
        RECT 548.400 25.350 549.600 26.100 ;
        RECT 554.400 25.350 555.600 26.100 ;
        RECT 568.950 25.950 571.050 28.050 ;
        RECT 578.400 27.600 579.450 43.950 ;
        RECT 587.400 34.050 588.450 46.950 ;
        RECT 605.400 46.050 606.450 59.100 ;
        RECT 608.400 54.900 609.450 67.950 ;
        RECT 617.400 60.600 618.450 85.950 ;
        RECT 617.400 58.350 618.600 60.600 ;
        RECT 622.950 59.100 625.050 61.200 ;
        RECT 623.400 58.350 624.600 59.100 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 614.400 54.900 615.600 55.650 ;
        RECT 620.400 54.900 621.600 55.650 ;
        RECT 607.950 52.800 610.050 54.900 ;
        RECT 613.950 52.800 616.050 54.900 ;
        RECT 619.950 52.800 622.050 54.900 ;
        RECT 604.950 43.950 607.050 46.050 ;
        RECT 605.400 40.050 606.450 43.950 ;
        RECT 604.950 37.950 607.050 40.050 ;
        RECT 586.950 31.950 589.050 34.050 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 551.400 21.000 552.600 22.650 ;
        RECT 557.400 21.000 558.600 22.650 ;
        RECT 569.400 21.900 570.450 25.950 ;
        RECT 578.400 25.350 579.600 27.600 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 575.400 21.900 576.600 22.650 ;
        RECT 550.950 16.950 553.050 21.000 ;
        RECT 556.950 16.950 559.050 21.000 ;
        RECT 568.950 19.800 571.050 21.900 ;
        RECT 574.950 19.800 577.050 21.900 ;
        RECT 581.400 21.450 582.600 22.650 ;
        RECT 587.400 21.450 588.450 31.950 ;
        RECT 598.950 26.100 601.050 28.200 ;
        RECT 604.950 26.100 607.050 28.200 ;
        RECT 610.950 26.100 613.050 28.200 ;
        RECT 625.950 26.100 628.050 28.200 ;
        RECT 632.400 27.600 633.450 97.800 ;
        RECT 641.400 95.700 642.300 104.700 ;
        RECT 648.000 103.800 650.100 104.700 ;
        RECT 651.000 102.900 651.900 108.300 ;
        RECT 652.950 104.100 655.050 106.200 ;
        RECT 653.400 103.350 654.600 104.100 ;
        RECT 645.000 101.700 651.900 102.900 ;
        RECT 645.000 99.300 645.900 101.700 ;
        RECT 643.800 97.200 645.900 99.300 ;
        RECT 646.800 97.950 648.900 100.050 ;
        RECT 640.500 93.600 642.600 95.700 ;
        RECT 647.400 95.400 648.600 97.650 ;
        RECT 650.700 94.500 651.900 101.700 ;
        RECT 652.800 100.950 654.900 103.050 ;
        RECT 650.100 92.400 652.200 94.500 ;
        RECT 656.400 70.050 657.450 163.950 ;
        RECT 658.950 160.950 661.050 163.050 ;
        RECT 659.400 130.050 660.450 160.950 ;
        RECT 671.400 145.050 672.450 220.950 ;
        RECT 674.400 157.050 675.450 253.950 ;
        RECT 679.950 229.950 682.050 232.050 ;
        RECT 680.400 216.600 681.450 229.950 ;
        RECT 683.400 220.050 684.450 265.950 ;
        RECT 686.400 258.600 687.450 274.950 ;
        RECT 698.400 274.050 699.450 295.950 ;
        RECT 700.950 289.950 703.050 295.050 ;
        RECT 704.400 283.050 705.450 295.950 ;
        RECT 706.950 294.600 711.000 295.050 ;
        RECT 706.950 292.950 711.600 294.600 ;
        RECT 715.950 294.000 718.050 298.050 ;
        RECT 710.400 292.350 711.600 292.950 ;
        RECT 716.400 292.350 717.600 294.000 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 713.400 287.400 714.600 289.650 ;
        RECT 719.400 287.400 720.600 289.650 ;
        RECT 703.950 280.950 706.050 283.050 ;
        RECT 713.400 274.050 714.450 287.400 ;
        RECT 719.400 283.050 720.450 287.400 ;
        RECT 718.950 280.950 721.050 283.050 ;
        RECT 725.400 274.050 726.450 346.950 ;
        RECT 737.400 343.050 738.450 355.950 ;
        RECT 740.400 355.050 741.450 364.950 ;
        RECT 746.400 355.050 747.450 379.950 ;
        RECT 755.400 376.050 756.450 410.400 ;
        RECT 763.950 409.800 766.050 411.900 ;
        RECT 767.400 409.050 768.450 415.950 ;
        RECT 757.950 406.950 760.050 409.050 ;
        RECT 766.950 406.950 769.050 409.050 ;
        RECT 758.400 403.050 759.450 406.950 ;
        RECT 757.950 400.950 760.050 403.050 ;
        RECT 763.950 400.950 766.050 403.050 ;
        RECT 748.950 373.950 751.050 376.050 ;
        RECT 749.400 366.900 750.450 373.950 ;
        RECT 751.950 370.950 754.050 376.050 ;
        RECT 754.950 373.950 757.050 376.050 ;
        RECT 757.950 372.000 760.050 376.050 ;
        RECT 764.400 373.050 765.450 400.950 ;
        RECT 770.400 382.050 771.450 418.950 ;
        RECT 772.950 417.450 775.050 421.050 ;
        RECT 782.400 417.600 783.450 439.950 ;
        RECT 785.400 421.050 786.450 442.950 ;
        RECT 790.950 441.450 793.050 444.900 ;
        RECT 788.400 441.000 793.050 441.450 ;
        RECT 788.400 440.400 792.450 441.000 ;
        RECT 788.400 436.050 789.450 440.400 ;
        RECT 794.400 438.450 795.450 463.950 ;
        RECT 796.950 457.950 799.050 460.050 ;
        RECT 791.400 437.400 795.450 438.450 ;
        RECT 787.950 433.950 790.050 436.050 ;
        RECT 784.950 418.950 787.050 421.050 ;
        RECT 776.400 417.450 777.600 417.600 ;
        RECT 772.950 417.000 777.600 417.450 ;
        RECT 773.400 416.400 777.600 417.000 ;
        RECT 776.400 415.350 777.600 416.400 ;
        RECT 782.400 415.350 783.600 417.600 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 772.950 409.950 775.050 412.050 ;
        RECT 779.400 411.900 780.600 412.650 ;
        RECT 769.950 379.950 772.050 382.050 ;
        RECT 758.400 370.350 759.600 372.000 ;
        RECT 763.950 370.950 766.050 373.050 ;
        RECT 767.100 370.950 769.200 373.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 767.400 368.400 768.600 370.650 ;
        RECT 755.400 366.900 756.600 367.650 ;
        RECT 748.950 364.800 751.050 366.900 ;
        RECT 754.950 364.800 757.050 366.900 ;
        RECT 761.400 365.400 762.600 367.650 ;
        RECT 739.950 352.950 742.050 355.050 ;
        RECT 745.950 352.950 748.050 355.050 ;
        RECT 727.950 340.950 730.050 343.050 ;
        RECT 730.950 342.450 735.000 343.050 ;
        RECT 730.950 340.950 735.450 342.450 ;
        RECT 736.950 340.950 739.050 343.050 ;
        RECT 728.400 319.050 729.450 340.950 ;
        RECT 734.400 339.600 735.450 340.950 ;
        RECT 740.400 339.600 741.450 352.950 ;
        RECT 749.400 343.050 750.450 364.800 ;
        RECT 761.400 361.050 762.450 365.400 ;
        RECT 763.950 364.950 766.050 367.050 ;
        RECT 760.950 358.950 763.050 361.050 ;
        RECT 751.950 352.950 754.050 355.050 ;
        RECT 748.950 340.950 751.050 343.050 ;
        RECT 734.400 337.350 735.600 339.600 ;
        RECT 740.400 337.350 741.600 339.600 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 737.400 333.900 738.600 334.650 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 743.400 333.000 744.600 334.650 ;
        RECT 742.950 328.950 745.050 333.000 ;
        RECT 752.400 325.050 753.450 352.950 ;
        RECT 764.400 342.450 765.450 364.950 ;
        RECT 767.400 349.050 768.450 368.400 ;
        RECT 769.950 367.950 772.050 370.050 ;
        RECT 766.950 346.950 769.050 349.050 ;
        RECT 770.400 346.050 771.450 367.950 ;
        RECT 769.950 343.950 772.050 346.050 ;
        RECT 764.400 341.400 771.450 342.450 ;
        RECT 754.950 337.950 757.050 340.050 ;
        RECT 763.950 338.100 766.050 340.200 ;
        RECT 770.400 339.600 771.450 341.400 ;
        RECT 773.400 340.050 774.450 409.950 ;
        RECT 778.950 409.800 781.050 411.900 ;
        RECT 785.400 410.400 786.600 412.650 ;
        RECT 785.400 403.050 786.450 410.400 ;
        RECT 784.950 400.950 787.050 403.050 ;
        RECT 791.400 394.050 792.450 437.400 ;
        RECT 793.950 433.950 796.050 436.050 ;
        RECT 794.400 397.050 795.450 433.950 ;
        RECT 797.400 433.050 798.450 457.950 ;
        RECT 796.950 430.950 799.050 433.050 ;
        RECT 800.400 418.050 801.450 481.800 ;
        RECT 812.400 478.050 813.450 481.950 ;
        RECT 818.400 481.050 819.450 490.800 ;
        RECT 817.950 478.950 820.050 481.050 ;
        RECT 802.950 475.950 805.050 478.050 ;
        RECT 808.950 476.400 813.450 478.050 ;
        RECT 808.950 475.950 813.000 476.400 ;
        RECT 814.950 475.950 817.050 478.050 ;
        RECT 803.400 451.050 804.450 475.950 ;
        RECT 811.950 472.950 814.050 475.050 ;
        RECT 812.400 469.050 813.450 472.950 ;
        RECT 811.950 466.950 814.050 469.050 ;
        RECT 808.950 463.950 811.050 466.050 ;
        RECT 809.400 460.050 810.450 463.950 ;
        RECT 808.950 457.950 811.050 460.050 ;
        RECT 802.950 448.950 805.050 451.050 ;
        RECT 805.950 450.000 808.050 454.050 ;
        RECT 812.400 451.050 813.450 466.950 ;
        RECT 806.400 448.350 807.600 450.000 ;
        RECT 811.950 448.950 814.050 451.050 ;
        RECT 805.950 445.950 808.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 809.400 444.900 810.600 445.650 ;
        RECT 815.400 445.050 816.450 475.950 ;
        RECT 818.400 469.050 819.450 478.950 ;
        RECT 817.950 466.950 820.050 469.050 ;
        RECT 817.950 463.800 820.050 465.900 ;
        RECT 808.950 442.800 811.050 444.900 ;
        RECT 814.950 442.950 817.050 445.050 ;
        RECT 814.950 439.800 817.050 441.900 ;
        RECT 811.950 436.950 814.050 439.050 ;
        RECT 802.950 430.950 805.050 433.050 ;
        RECT 799.950 415.950 802.050 418.050 ;
        RECT 803.400 417.600 804.450 430.950 ;
        RECT 803.400 415.350 804.600 417.600 ;
        RECT 802.950 412.950 805.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 806.400 411.900 807.600 412.650 ;
        RECT 805.950 409.800 808.050 411.900 ;
        RECT 793.950 394.950 796.050 397.050 ;
        RECT 802.950 394.950 805.050 397.050 ;
        RECT 790.950 391.950 793.050 394.050 ;
        RECT 781.950 385.950 784.050 388.050 ;
        RECT 776.100 370.950 778.200 373.050 ;
        RECT 776.400 369.900 777.600 370.650 ;
        RECT 775.950 367.800 778.050 369.900 ;
        RECT 776.400 361.050 777.450 367.800 ;
        RECT 782.400 367.050 783.450 385.950 ;
        RECT 785.700 384.300 787.800 386.400 ;
        RECT 786.300 379.500 787.800 384.300 ;
        RECT 785.700 377.400 787.800 379.500 ;
        RECT 781.950 364.950 784.050 367.050 ;
        RECT 775.950 358.950 778.050 361.050 ;
        RECT 781.950 358.950 784.050 361.050 ;
        RECT 786.300 359.700 787.800 377.400 ;
        RECT 782.400 355.050 783.450 358.950 ;
        RECT 785.700 357.600 787.800 359.700 ;
        RECT 788.700 381.300 790.800 386.400 ;
        RECT 791.700 384.300 793.800 386.400 ;
        RECT 788.700 359.700 789.900 381.300 ;
        RECT 791.700 379.500 793.200 384.300 ;
        RECT 794.100 381.300 796.200 383.400 ;
        RECT 791.100 377.400 793.200 379.500 ;
        RECT 791.700 359.700 793.200 377.400 ;
        RECT 794.700 374.100 795.900 381.300 ;
        RECT 799.500 379.800 801.600 381.900 ;
        RECT 794.100 372.000 796.200 374.100 ;
        RECT 800.700 373.200 801.600 379.800 ;
        RECT 803.400 376.050 804.450 394.950 ;
        RECT 806.400 388.050 807.450 409.800 ;
        RECT 812.400 391.050 813.450 436.950 ;
        RECT 815.400 397.050 816.450 439.800 ;
        RECT 818.400 433.050 819.450 463.800 ;
        RECT 821.400 460.050 822.450 493.800 ;
        RECT 820.950 457.950 823.050 460.050 ;
        RECT 820.950 454.800 823.050 456.900 ;
        RECT 817.950 430.950 820.050 433.050 ;
        RECT 821.400 427.050 822.450 454.800 ;
        RECT 824.400 451.050 825.450 505.950 ;
        RECT 829.950 499.950 832.050 502.050 ;
        RECT 826.950 493.950 829.050 496.050 ;
        RECT 827.400 466.050 828.450 493.950 ;
        RECT 826.950 463.950 829.050 466.050 ;
        RECT 826.950 457.950 829.050 460.050 ;
        RECT 823.950 448.950 826.050 451.050 ;
        RECT 827.400 450.600 828.450 457.950 ;
        RECT 830.400 453.450 831.450 499.950 ;
        RECT 833.400 496.050 834.450 512.400 ;
        RECT 836.400 502.050 837.450 526.800 ;
        RECT 839.400 514.050 840.450 571.950 ;
        RECT 842.400 534.450 843.450 580.950 ;
        RECT 845.400 541.050 846.450 589.800 ;
        RECT 848.400 574.050 849.450 611.400 ;
        RECT 859.950 610.950 862.050 613.050 ;
        RECT 868.950 610.950 871.050 613.050 ;
        RECT 850.950 607.950 853.050 610.050 ;
        RECT 851.400 598.050 852.450 607.950 ;
        RECT 856.950 605.100 859.050 607.200 ;
        RECT 862.950 605.100 865.050 607.200 ;
        RECT 857.400 604.350 858.600 605.100 ;
        RECT 863.400 604.350 864.600 605.100 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 853.950 598.950 856.050 601.050 ;
        RECT 860.400 599.400 861.600 601.650 ;
        RECT 850.950 595.950 853.050 598.050 ;
        RECT 854.400 592.050 855.450 598.950 ;
        RECT 860.400 595.050 861.450 599.400 ;
        RECT 862.950 595.050 865.050 598.050 ;
        RECT 859.950 592.950 862.050 595.050 ;
        RECT 862.950 594.000 868.050 595.050 ;
        RECT 863.400 593.400 868.050 594.000 ;
        RECT 864.000 592.950 868.050 593.400 ;
        RECT 853.950 589.950 856.050 592.050 ;
        RECT 850.950 586.950 853.050 589.050 ;
        RECT 847.950 571.950 850.050 574.050 ;
        RECT 851.400 573.600 852.450 586.950 ;
        RECT 856.950 583.950 859.050 586.050 ;
        RECT 857.400 573.600 858.450 583.950 ;
        RECT 869.400 583.050 870.450 610.950 ;
        RECT 871.950 604.950 874.050 607.050 ;
        RECT 872.400 586.050 873.450 604.950 ;
        RECT 871.950 583.950 874.050 586.050 ;
        RECT 868.950 580.950 871.050 583.050 ;
        RECT 865.950 577.950 868.050 580.050 ;
        RECT 851.400 571.350 852.600 573.600 ;
        RECT 857.400 571.350 858.600 573.600 ;
        RECT 866.400 571.050 867.450 577.950 ;
        RECT 871.950 574.950 874.050 577.050 ;
        RECT 868.950 571.950 871.050 574.050 ;
        RECT 850.950 568.950 853.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 854.400 567.000 855.600 568.650 ;
        RECT 860.400 567.000 861.600 568.650 ;
        RECT 853.950 562.950 856.050 567.000 ;
        RECT 859.950 562.950 862.050 567.000 ;
        RECT 865.950 559.950 868.050 562.050 ;
        RECT 850.950 556.950 853.050 559.050 ;
        RECT 862.950 556.950 865.050 559.050 ;
        RECT 847.950 550.950 850.050 553.050 ;
        RECT 844.950 538.950 847.050 541.050 ;
        RECT 842.400 533.400 846.450 534.450 ;
        RECT 841.950 529.950 844.050 532.050 ;
        RECT 842.400 514.050 843.450 529.950 ;
        RECT 845.400 529.050 846.450 533.400 ;
        RECT 848.400 532.050 849.450 550.950 ;
        RECT 851.400 535.050 852.450 556.950 ;
        RECT 859.950 547.950 862.050 550.050 ;
        RECT 853.950 544.950 856.050 547.050 ;
        RECT 850.950 532.950 853.050 535.050 ;
        RECT 847.950 529.950 850.050 532.050 ;
        RECT 854.400 531.450 855.450 544.950 ;
        RECT 851.400 530.400 855.450 531.450 ;
        RECT 844.950 526.950 847.050 529.050 ;
        RECT 851.400 528.600 852.450 530.400 ;
        RECT 851.400 526.350 852.600 528.600 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 850.950 523.950 853.050 526.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 848.400 523.050 849.600 523.650 ;
        RECT 844.950 521.400 849.600 523.050 ;
        RECT 854.400 523.050 855.600 523.650 ;
        RECT 854.400 521.400 859.050 523.050 ;
        RECT 844.950 520.950 849.000 521.400 ;
        RECT 855.000 520.950 859.050 521.400 ;
        RECT 838.950 511.950 841.050 514.050 ;
        RECT 841.950 511.950 844.050 514.050 ;
        RECT 844.950 511.950 847.050 514.050 ;
        RECT 850.950 511.950 853.050 514.050 ;
        RECT 841.950 508.800 844.050 510.900 ;
        RECT 838.950 502.950 841.050 505.050 ;
        RECT 835.950 499.950 838.050 502.050 ;
        RECT 839.400 499.050 840.450 502.950 ;
        RECT 837.000 498.900 840.450 499.050 ;
        RECT 835.950 497.400 840.450 498.900 ;
        RECT 835.950 496.950 840.000 497.400 ;
        RECT 835.950 496.800 838.050 496.950 ;
        RECT 842.400 496.050 843.450 508.800 ;
        RECT 832.950 495.450 835.050 496.050 ;
        RECT 836.400 495.450 837.600 495.600 ;
        RECT 832.950 494.400 837.600 495.450 ;
        RECT 832.950 493.950 835.050 494.400 ;
        RECT 836.400 493.350 837.600 494.400 ;
        RECT 841.950 493.950 844.050 496.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 832.950 487.950 835.050 490.050 ;
        RECT 839.400 488.400 840.600 490.650 ;
        RECT 833.400 484.050 834.450 487.950 ;
        RECT 839.400 484.050 840.450 488.400 ;
        RECT 841.950 487.950 844.050 490.050 ;
        RECT 832.950 481.950 835.050 484.050 ;
        RECT 838.950 481.950 841.050 484.050 ;
        RECT 838.950 469.950 841.050 472.050 ;
        RECT 839.400 460.050 840.450 469.950 ;
        RECT 838.950 457.950 841.050 460.050 ;
        RECT 842.400 456.450 843.450 487.950 ;
        RECT 845.400 472.050 846.450 511.950 ;
        RECT 851.400 507.450 852.450 511.950 ;
        RECT 848.400 506.400 852.450 507.450 ;
        RECT 844.950 469.950 847.050 472.050 ;
        RECT 844.950 463.950 847.050 466.050 ;
        RECT 839.400 455.400 843.450 456.450 ;
        RECT 830.400 452.400 834.450 453.450 ;
        RECT 833.400 450.600 834.450 452.400 ;
        RECT 839.400 451.050 840.450 455.400 ;
        RECT 841.950 451.950 844.050 454.050 ;
        RECT 827.400 448.350 828.600 450.600 ;
        RECT 833.400 448.350 834.600 450.600 ;
        RECT 838.950 448.950 841.050 451.050 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 830.400 443.400 831.600 445.650 ;
        RECT 836.400 444.900 837.600 445.650 ;
        RECT 823.950 433.950 826.050 436.050 ;
        RECT 824.400 430.050 825.450 433.950 ;
        RECT 830.400 433.050 831.450 443.400 ;
        RECT 835.950 442.800 838.050 444.900 ;
        RECT 838.950 442.950 841.050 445.050 ;
        RECT 839.400 435.450 840.450 442.950 ;
        RECT 836.400 434.400 840.450 435.450 ;
        RECT 829.950 430.950 832.050 433.050 ;
        RECT 823.950 427.950 826.050 430.050 ;
        RECT 820.950 424.950 823.050 427.050 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 817.950 415.950 820.050 418.050 ;
        RECT 823.950 416.100 826.050 418.200 ;
        RECT 830.400 417.600 831.450 424.950 ;
        RECT 836.400 418.050 837.450 434.400 ;
        RECT 838.950 430.950 841.050 433.050 ;
        RECT 814.950 394.950 817.050 397.050 ;
        RECT 818.400 393.450 819.450 415.950 ;
        RECT 824.400 415.350 825.600 416.100 ;
        RECT 830.400 415.350 831.600 417.600 ;
        RECT 835.950 415.950 838.050 418.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 827.400 410.400 828.600 412.650 ;
        RECT 833.400 411.900 834.600 412.650 ;
        RECT 827.400 394.050 828.450 410.400 ;
        RECT 832.950 409.800 835.050 411.900 ;
        RECT 829.950 406.950 832.050 409.050 ;
        RECT 830.400 403.050 831.450 406.950 ;
        RECT 829.950 400.950 832.050 403.050 ;
        RECT 818.400 392.400 822.450 393.450 ;
        RECT 811.950 388.950 814.050 391.050 ;
        RECT 817.950 388.950 820.050 391.050 ;
        RECT 805.950 385.950 808.050 388.050 ;
        RECT 810.600 384.300 812.700 386.400 ;
        RECT 813.600 384.300 816.600 386.400 ;
        RECT 808.200 381.300 810.300 383.400 ;
        RECT 805.950 376.950 808.050 379.050 ;
        RECT 802.950 373.950 805.050 376.050 ;
        RECT 794.700 359.700 795.900 372.000 ;
        RECT 799.500 371.100 801.600 373.200 ;
        RECT 796.800 364.500 798.900 366.600 ;
        RECT 800.700 360.600 801.600 371.100 ;
        RECT 802.800 368.100 804.900 370.200 ;
        RECT 806.400 370.050 807.450 376.950 ;
        RECT 803.400 367.350 804.600 368.100 ;
        RECT 805.950 367.950 808.050 370.050 ;
        RECT 803.100 364.950 805.200 367.050 ;
        RECT 788.700 357.600 790.800 359.700 ;
        RECT 791.700 357.600 793.800 359.700 ;
        RECT 794.700 357.600 796.800 359.700 ;
        RECT 800.100 358.500 802.200 360.600 ;
        RECT 809.100 359.700 810.300 381.300 ;
        RECT 811.500 378.300 812.700 384.300 ;
        RECT 811.500 376.200 813.600 378.300 ;
        RECT 811.500 359.700 812.700 376.200 ;
        RECT 815.100 365.400 816.600 384.300 ;
        RECT 814.500 363.300 816.600 365.400 ;
        RECT 814.500 359.700 815.700 363.300 ;
        RECT 808.200 357.600 810.300 359.700 ;
        RECT 811.200 357.600 813.300 359.700 ;
        RECT 814.200 357.600 816.300 359.700 ;
        RECT 775.950 352.950 778.050 355.050 ;
        RECT 781.950 352.950 784.050 355.050 ;
        RECT 755.400 331.050 756.450 337.950 ;
        RECT 764.400 337.350 765.600 338.100 ;
        RECT 770.400 337.350 771.600 339.600 ;
        RECT 772.950 337.950 775.050 340.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 757.950 331.950 760.050 334.050 ;
        RECT 761.400 332.400 762.600 334.650 ;
        RECT 767.400 332.400 768.600 334.650 ;
        RECT 754.950 328.950 757.050 331.050 ;
        RECT 745.950 322.950 748.050 325.050 ;
        RECT 751.950 322.950 754.050 325.050 ;
        RECT 727.950 316.950 730.050 319.050 ;
        RECT 730.950 310.950 733.050 313.050 ;
        RECT 727.950 286.800 730.050 288.900 ;
        RECT 691.950 271.950 694.050 274.050 ;
        RECT 697.950 271.950 700.050 274.050 ;
        RECT 712.950 271.950 715.050 274.050 ;
        RECT 724.950 271.950 727.050 274.050 ;
        RECT 686.400 256.350 687.600 258.600 ;
        RECT 686.100 253.950 688.200 256.050 ;
        RECT 692.400 229.050 693.450 271.950 ;
        RECT 695.700 267.300 697.800 269.400 ;
        RECT 696.300 249.600 697.800 267.300 ;
        RECT 695.700 247.500 697.800 249.600 ;
        RECT 696.300 242.700 697.800 247.500 ;
        RECT 695.700 240.600 697.800 242.700 ;
        RECT 698.700 267.300 700.800 269.400 ;
        RECT 701.700 267.300 703.800 269.400 ;
        RECT 704.700 267.300 706.800 269.400 ;
        RECT 698.700 245.700 699.900 267.300 ;
        RECT 701.700 249.600 703.200 267.300 ;
        RECT 704.700 255.000 705.900 267.300 ;
        RECT 710.100 266.400 712.200 268.500 ;
        RECT 718.200 267.300 720.300 269.400 ;
        RECT 721.200 267.300 723.300 269.400 ;
        RECT 724.200 267.300 726.300 269.400 ;
        RECT 706.800 260.400 708.900 262.500 ;
        RECT 710.700 255.900 711.600 266.400 ;
        RECT 713.100 259.950 715.200 262.050 ;
        RECT 713.400 258.900 714.600 259.650 ;
        RECT 712.950 256.800 715.050 258.900 ;
        RECT 704.100 252.900 706.200 255.000 ;
        RECT 709.500 253.800 711.600 255.900 ;
        RECT 701.100 247.500 703.200 249.600 ;
        RECT 698.700 240.600 700.800 245.700 ;
        RECT 701.700 242.700 703.200 247.500 ;
        RECT 704.700 245.700 705.900 252.900 ;
        RECT 710.700 247.200 711.600 253.800 ;
        RECT 704.100 243.600 706.200 245.700 ;
        RECT 709.500 245.100 711.600 247.200 ;
        RECT 719.100 245.700 720.300 267.300 ;
        RECT 718.200 243.600 720.300 245.700 ;
        RECT 721.500 250.800 722.700 267.300 ;
        RECT 724.500 263.700 725.700 267.300 ;
        RECT 724.500 261.600 726.600 263.700 ;
        RECT 721.500 248.700 723.600 250.800 ;
        RECT 721.500 242.700 722.700 248.700 ;
        RECT 725.100 242.700 726.600 261.600 ;
        RECT 728.400 250.050 729.450 286.800 ;
        RECT 731.400 283.050 732.450 310.950 ;
        RECT 741.000 297.450 745.050 298.050 ;
        RECT 740.400 295.950 745.050 297.450 ;
        RECT 740.400 294.600 741.450 295.950 ;
        RECT 746.400 295.050 747.450 322.950 ;
        RECT 758.400 322.050 759.450 331.950 ;
        RECT 751.950 319.800 754.050 321.900 ;
        RECT 757.950 319.950 760.050 322.050 ;
        RECT 740.400 292.350 741.600 294.600 ;
        RECT 745.950 292.950 748.050 295.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 737.400 288.900 738.600 289.650 ;
        RECT 736.950 286.800 739.050 288.900 ;
        RECT 743.400 287.400 744.600 289.650 ;
        RECT 743.400 283.050 744.450 287.400 ;
        RECT 730.950 280.950 733.050 283.050 ;
        RECT 742.950 280.950 745.050 283.050 ;
        RECT 745.950 271.950 748.050 274.050 ;
        RECT 731.100 253.950 733.200 256.050 ;
        RECT 737.100 253.950 739.200 256.050 ;
        RECT 737.400 252.000 738.600 253.650 ;
        RECT 727.950 247.950 730.050 250.050 ;
        RECT 736.950 247.950 739.050 252.000 ;
        RECT 701.700 240.600 703.800 242.700 ;
        RECT 720.600 240.600 722.700 242.700 ;
        RECT 723.600 240.600 726.600 242.700 ;
        RECT 724.950 235.950 727.050 238.050 ;
        RECT 691.950 226.950 694.050 229.050 ;
        RECT 712.950 226.950 715.050 229.050 ;
        RECT 682.950 217.950 685.050 220.050 ;
        RECT 680.400 214.350 681.600 216.600 ;
        RECT 685.950 215.100 688.050 217.200 ;
        RECT 691.950 216.000 694.050 220.050 ;
        RECT 686.400 214.350 687.600 215.100 ;
        RECT 692.400 214.350 693.600 216.000 ;
        RECT 697.950 214.950 700.050 217.050 ;
        RECT 703.950 215.100 706.050 217.200 ;
        RECT 713.400 216.600 714.450 226.950 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 683.400 209.400 684.600 211.650 ;
        RECT 689.400 210.000 690.600 211.650 ;
        RECT 683.400 202.050 684.450 209.400 ;
        RECT 688.950 205.950 691.050 210.000 ;
        RECT 682.950 199.950 685.050 202.050 ;
        RECT 682.950 187.950 685.050 190.050 ;
        RECT 676.950 182.100 679.050 184.200 ;
        RECT 683.400 183.600 684.450 187.950 ;
        RECT 677.400 172.050 678.450 182.100 ;
        RECT 683.400 181.350 684.600 183.600 ;
        RECT 688.950 182.100 691.050 184.200 ;
        RECT 689.400 181.350 690.600 182.100 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 685.950 178.950 688.050 181.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 691.950 178.950 694.050 181.050 ;
        RECT 686.400 176.400 687.600 178.650 ;
        RECT 692.400 177.900 693.600 178.650 ;
        RECT 686.400 175.050 687.450 176.400 ;
        RECT 691.950 175.800 694.050 177.900 ;
        RECT 685.950 172.950 688.050 175.050 ;
        RECT 676.950 169.950 679.050 172.050 ;
        RECT 673.950 154.950 676.050 157.050 ;
        RECT 677.400 145.050 678.450 169.950 ;
        RECT 664.950 142.950 667.050 145.050 ;
        RECT 670.950 142.950 673.050 145.050 ;
        RECT 676.950 142.950 679.050 145.050 ;
        RECT 661.950 137.100 664.050 139.200 ;
        RECT 658.950 127.950 661.050 130.050 ;
        RECT 662.400 124.050 663.450 137.100 ;
        RECT 665.400 130.050 666.450 142.950 ;
        RECT 679.950 139.950 682.050 145.050 ;
        RECT 670.950 137.100 673.050 139.200 ;
        RECT 676.950 137.100 679.050 139.200 ;
        RECT 671.400 136.350 672.600 137.100 ;
        RECT 677.400 136.350 678.600 137.100 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 674.400 131.400 675.600 133.650 ;
        RECT 674.400 130.050 675.450 131.400 ;
        RECT 682.950 130.800 685.050 132.900 ;
        RECT 664.950 127.950 667.050 130.050 ;
        RECT 670.950 128.400 675.450 130.050 ;
        RECT 670.950 127.950 675.000 128.400 ;
        RECT 676.950 127.950 679.050 130.050 ;
        RECT 661.950 121.950 664.050 124.050 ;
        RECT 677.400 118.050 678.450 127.950 ;
        RECT 683.400 124.050 684.450 130.800 ;
        RECT 682.950 121.950 685.050 124.050 ;
        RECT 664.950 115.950 667.050 118.050 ;
        RECT 676.950 115.950 679.050 118.050 ;
        RECT 658.950 112.950 661.050 115.050 ;
        RECT 659.400 106.200 660.450 112.950 ;
        RECT 658.950 104.100 661.050 106.200 ;
        RECT 665.400 99.900 666.450 115.950 ;
        RECT 679.950 109.950 682.050 112.050 ;
        RECT 673.950 104.100 676.050 106.200 ;
        RECT 680.400 105.600 681.450 109.950 ;
        RECT 686.400 106.050 687.450 172.950 ;
        RECT 698.400 166.050 699.450 214.950 ;
        RECT 704.400 211.050 705.450 215.100 ;
        RECT 713.400 214.350 714.600 216.600 ;
        RECT 718.950 215.100 721.050 217.200 ;
        RECT 725.400 217.050 726.450 235.950 ;
        RECT 727.950 223.950 730.050 226.050 ;
        RECT 719.400 214.350 720.600 215.100 ;
        RECT 724.950 214.950 727.050 217.050 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 703.950 208.950 706.050 211.050 ;
        RECT 710.400 209.400 711.600 211.650 ;
        RECT 716.400 210.900 717.600 211.650 ;
        RECT 725.400 210.900 726.450 214.950 ;
        RECT 703.950 193.950 706.050 196.050 ;
        RECT 700.950 181.950 703.050 184.050 ;
        RECT 701.400 177.900 702.450 181.950 ;
        RECT 700.950 175.800 703.050 177.900 ;
        RECT 700.950 166.950 703.050 169.050 ;
        RECT 697.950 163.950 700.050 166.050 ;
        RECT 701.400 148.050 702.450 166.950 ;
        RECT 704.400 151.050 705.450 193.950 ;
        RECT 710.400 190.050 711.450 209.400 ;
        RECT 715.950 208.800 718.050 210.900 ;
        RECT 724.950 208.800 727.050 210.900 ;
        RECT 712.950 193.950 715.050 196.050 ;
        RECT 709.950 187.950 712.050 190.050 ;
        RECT 713.400 184.200 714.450 193.950 ;
        RECT 718.950 187.950 721.050 190.050 ;
        RECT 712.950 182.100 715.050 184.200 ;
        RECT 713.400 181.350 714.600 182.100 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 710.400 176.400 711.600 178.650 ;
        RECT 710.400 160.050 711.450 176.400 ;
        RECT 709.950 157.950 712.050 160.050 ;
        RECT 703.950 148.950 706.050 151.050 ;
        RECT 715.950 148.950 718.050 151.050 ;
        RECT 700.950 145.950 703.050 148.050 ;
        RECT 688.950 142.950 691.050 145.050 ;
        RECT 689.400 123.450 690.450 142.950 ;
        RECT 698.100 142.500 700.200 144.600 ;
        RECT 691.950 139.950 694.050 142.050 ;
        RECT 692.400 127.050 693.450 139.950 ;
        RECT 695.100 133.950 697.200 136.050 ;
        RECT 698.100 135.900 699.000 142.500 ;
        RECT 707.100 142.200 709.200 144.300 ;
        RECT 712.950 142.950 715.050 145.050 ;
        RECT 701.400 139.350 702.600 141.600 ;
        RECT 700.800 136.950 702.900 139.050 ;
        RECT 705.000 135.900 707.100 136.200 ;
        RECT 698.100 135.000 707.100 135.900 ;
        RECT 695.400 132.900 696.600 133.650 ;
        RECT 694.950 130.800 697.050 132.900 ;
        RECT 698.100 129.900 699.000 135.000 ;
        RECT 705.000 134.100 707.100 135.000 ;
        RECT 699.900 133.200 702.000 134.100 ;
        RECT 699.900 132.000 707.100 133.200 ;
        RECT 705.000 131.100 707.100 132.000 ;
        RECT 697.500 127.800 699.600 129.900 ;
        RECT 700.800 128.100 702.900 130.200 ;
        RECT 708.000 129.600 708.900 142.200 ;
        RECT 709.950 138.450 712.050 139.200 ;
        RECT 713.400 138.450 714.450 142.950 ;
        RECT 709.950 137.400 714.450 138.450 ;
        RECT 709.950 137.100 712.050 137.400 ;
        RECT 710.400 136.350 711.600 137.100 ;
        RECT 709.800 133.950 711.900 136.050 ;
        RECT 716.400 132.900 717.450 148.950 ;
        RECT 715.950 130.800 718.050 132.900 ;
        RECT 701.400 127.050 702.600 127.800 ;
        RECT 707.400 127.500 709.500 129.600 ;
        RECT 691.950 124.950 694.050 127.050 ;
        RECT 700.950 124.950 703.050 127.050 ;
        RECT 689.400 122.400 696.450 123.450 ;
        RECT 695.400 120.450 696.450 122.400 ;
        RECT 706.950 121.950 709.050 124.050 ;
        RECT 695.400 119.400 699.450 120.450 ;
        RECT 694.950 115.950 697.050 118.050 ;
        RECT 691.950 109.950 694.050 112.050 ;
        RECT 674.400 103.350 675.600 104.100 ;
        RECT 680.400 103.350 681.600 105.600 ;
        RECT 685.950 103.950 688.050 106.050 ;
        RECT 688.950 103.950 691.050 106.050 ;
        RECT 670.950 100.950 673.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 664.950 97.800 667.050 99.900 ;
        RECT 671.400 98.400 672.600 100.650 ;
        RECT 677.400 99.900 678.600 100.650 ;
        RECT 671.400 96.450 672.450 98.400 ;
        RECT 676.950 97.800 679.050 99.900 ;
        RECT 689.400 97.050 690.450 103.950 ;
        RECT 692.400 99.900 693.450 109.950 ;
        RECT 695.400 106.050 696.450 115.950 ;
        RECT 698.400 108.450 699.450 119.400 ;
        RECT 698.400 107.400 702.450 108.450 ;
        RECT 694.950 103.950 697.050 106.050 ;
        RECT 701.400 105.600 702.450 107.400 ;
        RECT 707.400 105.600 708.450 121.950 ;
        RECT 701.400 103.350 702.600 105.600 ;
        RECT 707.400 103.350 708.600 105.600 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 712.950 102.000 715.050 106.050 ;
        RECT 698.400 99.900 699.600 100.650 ;
        RECT 691.950 97.800 694.050 99.900 ;
        RECT 697.950 97.800 700.050 99.900 ;
        RECT 704.400 99.000 705.600 100.650 ;
        RECT 713.400 100.350 714.600 102.000 ;
        RECT 671.400 95.400 675.450 96.450 ;
        RECT 674.400 85.050 675.450 95.400 ;
        RECT 688.950 94.950 691.050 97.050 ;
        RECT 703.950 94.950 706.050 99.000 ;
        RECT 713.100 97.950 715.200 100.050 ;
        RECT 703.950 85.950 706.050 88.050 ;
        RECT 673.950 82.950 676.050 85.050 ;
        RECT 655.950 67.950 658.050 70.050 ;
        RECT 634.950 59.100 637.050 61.200 ;
        RECT 640.950 59.100 643.050 61.200 ;
        RECT 646.950 59.100 649.050 61.200 ;
        RECT 652.950 59.100 655.050 61.200 ;
        RECT 658.950 59.100 661.050 61.200 ;
        RECT 664.950 59.100 667.050 61.200 ;
        RECT 670.950 60.000 673.050 64.050 ;
        RECT 674.400 61.050 675.450 82.950 ;
        RECT 697.950 64.950 700.050 67.050 ;
        RECT 676.950 61.950 679.050 64.050 ;
        RECT 635.400 55.050 636.450 59.100 ;
        RECT 641.400 58.350 642.600 59.100 ;
        RECT 647.400 58.350 648.600 59.100 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 634.950 52.950 637.050 55.050 ;
        RECT 644.400 54.900 645.600 55.650 ;
        RECT 643.950 52.800 646.050 54.900 ;
        RECT 653.400 49.050 654.450 59.100 ;
        RECT 659.400 55.050 660.450 59.100 ;
        RECT 665.400 58.350 666.600 59.100 ;
        RECT 671.400 58.350 672.600 60.000 ;
        RECT 673.950 58.950 676.050 61.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 668.400 54.900 669.600 55.650 ;
        RECT 667.950 52.800 670.050 54.900 ;
        RECT 652.950 46.950 655.050 49.050 ;
        RECT 677.400 34.050 678.450 61.950 ;
        RECT 691.950 59.100 694.050 61.200 ;
        RECT 692.400 58.350 693.600 59.100 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 689.400 53.400 690.600 55.650 ;
        RECT 689.400 49.050 690.450 53.400 ;
        RECT 688.950 46.950 691.050 49.050 ;
        RECT 698.400 46.050 699.450 64.950 ;
        RECT 700.950 58.950 703.050 61.050 ;
        RECT 697.950 43.950 700.050 46.050 ;
        RECT 691.950 37.950 694.050 40.050 ;
        RECT 670.950 31.950 673.050 34.050 ;
        RECT 676.950 31.950 679.050 34.050 ;
        RECT 637.950 28.950 640.050 31.050 ;
        RECT 599.400 25.350 600.600 26.100 ;
        RECT 605.400 25.350 606.600 26.100 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 602.400 21.900 603.600 22.650 ;
        RECT 611.400 22.050 612.450 26.100 ;
        RECT 626.400 25.350 627.600 26.100 ;
        RECT 632.400 25.350 633.600 27.600 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 581.400 20.400 588.450 21.450 ;
        RECT 601.950 19.800 604.050 21.900 ;
        RECT 610.950 19.950 613.050 22.050 ;
        RECT 623.400 20.400 624.600 22.650 ;
        RECT 629.400 21.900 630.600 22.650 ;
        RECT 638.400 21.900 639.450 28.950 ;
        RECT 643.950 26.100 646.050 28.200 ;
        RECT 649.950 26.100 652.050 28.200 ;
        RECT 655.950 27.000 658.050 31.050 ;
        RECT 623.400 16.050 624.450 20.400 ;
        RECT 628.950 19.800 631.050 21.900 ;
        RECT 637.950 19.800 640.050 21.900 ;
        RECT 553.950 15.450 556.050 16.050 ;
        RECT 559.950 15.450 562.050 16.050 ;
        RECT 553.950 14.400 562.050 15.450 ;
        RECT 553.950 13.950 556.050 14.400 ;
        RECT 559.950 13.950 562.050 14.400 ;
        RECT 622.950 13.950 625.050 16.050 ;
        RECT 644.400 13.050 645.450 26.100 ;
        RECT 650.400 25.350 651.600 26.100 ;
        RECT 656.400 25.350 657.600 27.000 ;
        RECT 664.950 25.950 667.050 28.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 653.400 21.900 654.600 22.650 ;
        RECT 652.950 19.800 655.050 21.900 ;
        RECT 659.400 20.400 660.600 22.650 ;
        RECT 665.400 21.900 666.450 25.950 ;
        RECT 671.400 21.900 672.450 31.950 ;
        RECT 679.950 26.100 682.050 28.200 ;
        RECT 692.400 28.050 693.450 37.950 ;
        RECT 697.950 31.950 700.050 34.050 ;
        RECT 694.950 28.950 697.050 31.050 ;
        RECT 680.400 25.350 681.600 26.100 ;
        RECT 691.950 25.950 694.050 28.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 677.400 21.900 678.600 22.650 ;
        RECT 683.400 21.900 684.600 22.650 ;
        RECT 695.400 21.900 696.450 28.950 ;
        RECT 698.400 27.450 699.450 31.950 ;
        RECT 701.400 31.050 702.450 58.950 ;
        RECT 704.400 54.900 705.450 85.950 ;
        RECT 719.400 64.050 720.450 187.950 ;
        RECT 728.400 177.450 729.450 223.950 ;
        RECT 746.400 223.050 747.450 271.950 ;
        RECT 730.950 220.950 733.050 223.050 ;
        RECT 745.950 220.950 748.050 223.050 ;
        RECT 731.400 208.050 732.450 220.950 ;
        RECT 736.950 215.100 739.050 217.200 ;
        RECT 752.400 217.050 753.450 319.800 ;
        RECT 761.400 318.450 762.450 332.400 ;
        RECT 758.400 317.400 762.450 318.450 ;
        RECT 754.950 304.950 757.050 307.050 ;
        RECT 755.400 255.450 756.450 304.950 ;
        RECT 758.400 295.050 759.450 317.400 ;
        RECT 763.950 316.950 766.050 319.050 ;
        RECT 760.950 313.950 763.050 316.050 ;
        RECT 761.400 304.050 762.450 313.950 ;
        RECT 764.400 307.050 765.450 316.950 ;
        RECT 763.950 304.950 766.050 307.050 ;
        RECT 767.400 304.050 768.450 332.400 ;
        RECT 776.400 313.050 777.450 352.950 ;
        RECT 818.400 349.050 819.450 388.950 ;
        RECT 821.400 379.050 822.450 392.400 ;
        RECT 826.950 391.950 829.050 394.050 ;
        RECT 839.400 382.050 840.450 430.950 ;
        RECT 842.400 411.900 843.450 451.950 ;
        RECT 841.950 409.800 844.050 411.900 ;
        RECT 823.950 379.950 826.050 382.050 ;
        RECT 838.950 379.950 841.050 382.050 ;
        RECT 820.950 376.950 823.050 379.050 ;
        RECT 824.400 376.050 825.450 379.950 ;
        RECT 845.400 379.050 846.450 463.950 ;
        RECT 848.400 424.050 849.450 506.400 ;
        RECT 850.950 502.950 853.050 505.050 ;
        RECT 851.400 487.050 852.450 502.950 ;
        RECT 860.400 498.450 861.450 547.950 ;
        RECT 863.400 508.050 864.450 556.950 ;
        RECT 866.400 556.050 867.450 559.950 ;
        RECT 865.950 553.950 868.050 556.050 ;
        RECT 866.400 511.050 867.450 553.950 ;
        RECT 869.400 532.050 870.450 571.950 ;
        RECT 872.400 565.050 873.450 574.950 ;
        RECT 875.400 574.050 876.450 625.950 ;
        RECT 881.400 609.450 882.450 646.950 ;
        RECT 884.400 643.050 885.450 649.950 ;
        RECT 887.400 643.050 888.450 652.800 ;
        RECT 895.950 650.100 898.050 652.200 ;
        RECT 896.400 649.350 897.600 650.100 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 898.950 646.950 901.050 649.050 ;
        RECT 889.950 643.950 892.050 646.050 ;
        RECT 893.400 644.400 894.600 646.650 ;
        RECT 899.400 645.000 900.600 646.650 ;
        RECT 883.950 640.950 886.050 643.050 ;
        RECT 886.950 640.950 889.050 643.050 ;
        RECT 890.400 640.050 891.450 643.950 ;
        RECT 889.950 637.950 892.050 640.050 ;
        RECT 889.950 634.800 892.050 636.900 ;
        RECT 883.950 631.950 886.050 634.050 ;
        RECT 884.400 625.050 885.450 631.950 ;
        RECT 883.950 622.950 886.050 625.050 ;
        RECT 878.400 609.000 882.450 609.450 ;
        RECT 877.950 608.400 882.450 609.000 ;
        RECT 877.950 604.950 880.050 608.400 ;
        RECT 884.400 606.600 885.450 622.950 ;
        RECT 890.400 606.600 891.450 634.800 ;
        RECT 893.400 628.050 894.450 644.400 ;
        RECT 898.950 640.950 901.050 645.000 ;
        RECT 901.950 643.950 904.050 646.050 ;
        RECT 902.400 640.050 903.450 643.950 ;
        RECT 895.950 637.950 898.050 640.050 ;
        RECT 901.950 637.950 904.050 640.050 ;
        RECT 892.950 625.950 895.050 628.050 ;
        RECT 893.400 607.050 894.450 625.950 ;
        RECT 884.400 604.350 885.600 606.600 ;
        RECT 890.400 604.350 891.600 606.600 ;
        RECT 892.950 604.950 895.050 607.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 881.400 600.900 882.600 601.650 ;
        RECT 887.400 600.900 888.600 601.650 ;
        RECT 880.950 598.800 883.050 600.900 ;
        RECT 886.950 598.800 889.050 600.900 ;
        RECT 874.950 571.950 877.050 574.050 ;
        RECT 881.400 573.600 882.450 598.800 ;
        RECT 896.400 598.050 897.450 637.950 ;
        RECT 905.400 637.050 906.450 673.950 ;
        RECT 917.400 667.050 918.450 679.950 ;
        RECT 920.400 673.050 921.450 712.950 ;
        RECT 925.950 688.950 928.050 691.050 ;
        RECT 926.400 685.200 927.450 688.950 ;
        RECT 925.950 683.100 928.050 685.200 ;
        RECT 929.400 684.600 930.450 715.800 ;
        RECT 932.400 715.050 933.450 748.950 ;
        RECT 931.950 712.950 934.050 715.050 ;
        RECT 935.400 709.050 936.450 755.400 ;
        RECT 940.950 748.950 943.050 751.050 ;
        RECT 941.400 730.050 942.450 748.950 ;
        RECT 937.950 727.950 940.050 730.050 ;
        RECT 940.950 727.950 943.050 730.050 ;
        RECT 944.400 729.600 945.450 772.950 ;
        RECT 947.400 739.050 948.450 799.950 ;
        RECT 950.400 799.050 951.450 868.800 ;
        RECT 955.950 847.950 958.050 850.050 ;
        RECT 956.400 841.200 957.450 847.950 ;
        RECT 955.950 839.100 958.050 841.200 ;
        RECT 961.950 839.100 964.050 841.200 ;
        RECT 968.400 841.050 969.450 871.950 ;
        RECT 970.950 862.950 973.050 865.050 ;
        RECT 956.400 838.350 957.600 839.100 ;
        RECT 962.400 838.350 963.600 839.100 ;
        RECT 967.950 838.950 970.050 841.050 ;
        RECT 955.950 835.950 958.050 838.050 ;
        RECT 958.950 835.950 961.050 838.050 ;
        RECT 961.950 835.950 964.050 838.050 ;
        RECT 964.950 835.950 967.050 838.050 ;
        RECT 952.950 832.950 955.050 835.050 ;
        RECT 959.400 834.000 960.600 835.650 ;
        RECT 965.400 834.900 966.600 835.650 ;
        RECT 953.400 820.050 954.450 832.950 ;
        RECT 958.950 832.050 961.050 834.000 ;
        RECT 964.950 832.800 967.050 834.900 ;
        RECT 967.950 832.950 970.050 835.050 ;
        RECT 958.800 831.000 961.050 832.050 ;
        RECT 958.800 829.950 960.900 831.000 ;
        RECT 961.950 829.950 964.050 832.050 ;
        RECT 952.950 817.950 955.050 820.050 ;
        RECT 955.950 814.950 958.050 817.050 ;
        RECT 949.950 796.950 952.050 799.050 ;
        RECT 952.950 796.950 955.050 799.050 ;
        RECT 953.400 778.050 954.450 796.950 ;
        RECT 956.400 790.050 957.450 814.950 ;
        RECT 959.400 814.050 960.450 829.950 ;
        RECT 962.400 826.050 963.450 829.950 ;
        RECT 961.950 823.950 964.050 826.050 ;
        RECT 958.950 811.950 961.050 814.050 ;
        RECT 962.400 810.450 963.450 823.950 ;
        RECT 968.400 817.050 969.450 832.950 ;
        RECT 971.400 829.050 972.450 862.950 ;
        RECT 973.950 838.950 976.050 841.050 ;
        RECT 980.400 840.450 981.450 964.950 ;
        RECT 988.950 961.950 991.050 964.200 ;
        RECT 997.950 962.100 1000.050 964.200 ;
        RECT 1006.950 962.100 1009.050 964.200 ;
        RECT 1012.950 962.100 1015.050 964.200 ;
        RECT 1030.950 963.000 1033.050 967.050 ;
        RECT 998.400 961.350 999.600 962.100 ;
        RECT 1007.400 961.350 1008.600 962.100 ;
        RECT 992.400 958.950 994.500 961.050 ;
        RECT 997.950 958.950 1000.050 961.050 ;
        RECT 1000.950 958.950 1003.050 961.050 ;
        RECT 1007.100 958.950 1009.200 961.050 ;
        RECT 992.400 956.400 993.600 958.650 ;
        RECT 1001.400 957.900 1002.600 958.650 ;
        RECT 992.400 928.050 993.450 956.400 ;
        RECT 1000.950 955.800 1003.050 957.900 ;
        RECT 1009.950 955.800 1012.050 957.900 ;
        RECT 991.950 925.950 994.050 928.050 ;
        RECT 1006.950 922.950 1009.050 925.050 ;
        RECT 991.950 918.000 994.050 922.050 ;
        RECT 992.400 916.350 993.600 918.000 ;
        RECT 997.950 917.100 1000.050 919.200 ;
        RECT 998.400 916.350 999.600 917.100 ;
        RECT 991.950 913.950 994.050 916.050 ;
        RECT 994.950 913.950 997.050 916.050 ;
        RECT 997.950 913.950 1000.050 916.050 ;
        RECT 1000.950 913.950 1003.050 916.050 ;
        RECT 995.400 912.000 996.600 913.650 ;
        RECT 1001.400 912.450 1002.600 913.650 ;
        RECT 994.950 907.950 997.050 912.000 ;
        RECT 1001.400 911.400 1005.450 912.450 ;
        RECT 1000.950 907.950 1003.050 910.050 ;
        RECT 985.950 889.950 988.050 892.050 ;
        RECT 982.950 877.800 985.050 879.900 ;
        RECT 983.400 844.200 984.450 877.800 ;
        RECT 986.400 874.050 987.450 889.950 ;
        RECT 994.950 884.100 997.050 886.200 ;
        RECT 995.400 883.350 996.600 884.100 ;
        RECT 989.100 880.950 991.200 883.050 ;
        RECT 994.500 880.950 996.600 883.050 ;
        RECT 997.800 880.950 999.900 883.050 ;
        RECT 989.400 879.000 990.600 880.650 ;
        RECT 988.950 874.950 991.050 879.000 ;
        RECT 998.400 878.400 999.600 880.650 ;
        RECT 998.400 874.050 999.450 878.400 ;
        RECT 985.950 871.950 988.050 874.050 ;
        RECT 997.950 871.950 1000.050 874.050 ;
        RECT 997.950 868.800 1000.050 870.900 ;
        RECT 994.950 850.950 997.050 853.050 ;
        RECT 985.950 847.950 988.050 850.050 ;
        RECT 982.950 842.100 985.050 844.200 ;
        RECT 986.400 844.050 987.450 847.950 ;
        RECT 985.950 841.950 988.050 844.050 ;
        RECT 977.400 839.400 981.450 840.450 ;
        RECT 974.400 835.050 975.450 838.950 ;
        RECT 973.950 832.950 976.050 835.050 ;
        RECT 970.950 826.950 973.050 829.050 ;
        RECT 967.950 814.950 970.050 817.050 ;
        RECT 967.950 811.800 970.050 813.900 ;
        RECT 959.400 810.000 963.450 810.450 ;
        RECT 958.950 809.400 963.450 810.000 ;
        RECT 958.950 805.950 961.050 809.400 ;
        RECT 961.950 806.100 964.050 808.200 ;
        RECT 968.400 807.600 969.450 811.800 ;
        RECT 962.400 805.350 963.600 806.100 ;
        RECT 968.400 805.350 969.600 807.600 ;
        RECT 961.950 802.950 964.050 805.050 ;
        RECT 964.950 802.950 967.050 805.050 ;
        RECT 967.950 802.950 970.050 805.050 ;
        RECT 970.950 802.950 973.050 805.050 ;
        RECT 958.950 799.800 961.050 802.050 ;
        RECT 965.400 801.900 966.600 802.650 ;
        RECT 964.950 799.800 967.050 801.900 ;
        RECT 971.400 800.400 972.600 802.650 ;
        RECT 971.400 799.050 972.450 800.400 ;
        RECT 970.950 796.950 973.050 799.050 ;
        RECT 964.950 793.950 967.050 796.050 ;
        RECT 955.950 787.950 958.050 790.050 ;
        RECT 961.950 781.950 964.050 784.050 ;
        RECT 952.950 775.950 955.050 778.050 ;
        RECT 955.950 761.100 958.050 763.200 ;
        RECT 962.400 763.050 963.450 781.950 ;
        RECT 965.400 772.050 966.450 793.950 ;
        RECT 971.400 781.050 972.450 796.950 ;
        RECT 977.400 784.050 978.450 839.400 ;
        RECT 982.950 838.950 985.050 841.050 ;
        RECT 988.950 839.100 991.050 841.200 ;
        RECT 983.400 838.350 984.600 838.950 ;
        RECT 989.400 838.350 990.600 839.100 ;
        RECT 982.950 835.950 985.050 838.050 ;
        RECT 985.950 835.950 988.050 838.050 ;
        RECT 988.950 835.950 991.050 838.050 ;
        RECT 979.950 832.950 982.050 835.050 ;
        RECT 986.400 833.400 987.600 835.650 ;
        RECT 980.400 808.050 981.450 832.950 ;
        RECT 986.400 829.050 987.450 833.400 ;
        RECT 991.950 832.950 994.050 835.050 ;
        RECT 985.950 826.950 988.050 829.050 ;
        RECT 982.950 808.950 985.050 811.050 ;
        RECT 979.950 805.950 982.050 808.050 ;
        RECT 983.400 801.900 984.450 808.950 ;
        RECT 992.400 807.600 993.450 832.950 ;
        RECT 995.400 811.050 996.450 850.950 ;
        RECT 998.400 823.050 999.450 868.800 ;
        RECT 997.950 820.950 1000.050 823.050 ;
        RECT 994.950 808.950 997.050 811.050 ;
        RECT 998.400 808.050 999.450 820.950 ;
        RECT 992.400 805.350 993.600 807.600 ;
        RECT 997.950 805.950 1000.050 808.050 ;
        RECT 988.950 802.950 991.050 805.050 ;
        RECT 991.950 802.950 994.050 805.050 ;
        RECT 994.950 802.950 997.050 805.050 ;
        RECT 989.400 801.900 990.600 802.650 ;
        RECT 982.950 799.800 985.050 801.900 ;
        RECT 988.950 799.800 991.050 801.900 ;
        RECT 995.400 801.000 996.600 802.650 ;
        RECT 994.950 796.950 997.050 801.000 ;
        RECT 997.950 799.950 1000.050 802.050 ;
        RECT 979.950 790.950 982.050 796.050 ;
        RECT 991.950 784.950 994.050 787.050 ;
        RECT 976.950 781.950 979.050 784.050 ;
        RECT 988.950 781.950 991.050 784.050 ;
        RECT 970.950 778.950 973.050 781.050 ;
        RECT 967.950 775.950 970.050 778.050 ;
        RECT 968.400 772.050 969.450 775.950 ;
        RECT 964.800 769.950 966.900 772.050 ;
        RECT 967.950 769.950 970.050 772.050 ;
        RECT 967.950 763.950 970.050 766.050 ;
        RECT 956.400 760.350 957.600 761.100 ;
        RECT 961.950 760.950 964.050 763.050 ;
        RECT 964.950 760.950 967.050 763.050 ;
        RECT 952.950 757.950 955.050 760.050 ;
        RECT 955.950 757.950 958.050 760.050 ;
        RECT 958.950 757.950 961.050 760.050 ;
        RECT 953.400 756.900 954.600 757.650 ;
        RECT 952.950 754.800 955.050 756.900 ;
        RECT 959.400 755.400 960.600 757.650 ;
        RECT 959.400 751.050 960.450 755.400 ;
        RECT 961.950 754.950 964.050 757.050 ;
        RECT 958.950 748.950 961.050 751.050 ;
        RECT 946.950 736.950 949.050 739.050 ;
        RECT 949.950 733.950 952.050 736.050 ;
        RECT 950.400 729.600 951.450 733.950 ;
        RECT 958.950 730.950 961.050 733.050 ;
        RECT 938.400 718.050 939.450 727.950 ;
        RECT 944.400 727.350 945.600 729.600 ;
        RECT 950.400 727.350 951.600 729.600 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 946.950 724.950 949.050 727.050 ;
        RECT 949.950 724.950 952.050 727.050 ;
        RECT 952.950 724.950 955.050 727.050 ;
        RECT 947.400 723.900 948.600 724.650 ;
        RECT 953.400 723.900 954.600 724.650 ;
        RECT 940.950 718.950 943.050 723.900 ;
        RECT 946.950 721.800 949.050 723.900 ;
        RECT 952.950 721.800 955.050 723.900 ;
        RECT 937.950 715.950 940.050 718.050 ;
        RECT 934.950 706.950 937.050 709.050 ;
        RECT 949.950 703.950 952.050 706.050 ;
        RECT 934.950 697.950 937.050 700.050 ;
        RECT 935.400 688.050 936.450 697.950 ;
        RECT 946.950 694.950 949.050 697.050 ;
        RECT 934.950 685.950 937.050 688.050 ;
        RECT 929.400 682.350 930.600 684.600 ;
        RECT 937.950 683.100 940.050 685.200 ;
        RECT 947.400 685.050 948.450 694.950 ;
        RECT 938.400 682.350 939.600 683.100 ;
        RECT 946.950 682.950 949.050 685.050 ;
        RECT 929.400 679.950 931.500 682.050 ;
        RECT 934.950 679.950 937.050 682.050 ;
        RECT 937.950 679.950 940.050 682.050 ;
        RECT 944.100 679.950 946.200 682.050 ;
        RECT 925.950 676.950 928.050 679.050 ;
        RECT 935.400 677.400 936.600 679.650 ;
        RECT 944.400 678.900 945.600 679.650 ;
        RECT 931.950 673.950 934.050 676.050 ;
        RECT 919.950 670.950 922.050 673.050 ;
        RECT 928.950 670.950 931.050 673.050 ;
        RECT 916.950 664.950 919.050 667.050 ;
        RECT 916.950 658.950 919.050 661.050 ;
        RECT 910.950 655.950 913.050 658.050 ;
        RECT 907.950 649.950 910.050 652.050 ;
        RECT 898.950 634.950 901.050 637.050 ;
        RECT 904.950 634.950 907.050 637.050 ;
        RECT 889.950 595.950 892.050 598.050 ;
        RECT 895.950 595.950 898.050 598.050 ;
        RECT 881.400 571.350 882.600 573.600 ;
        RECT 886.950 573.000 889.050 577.050 ;
        RECT 890.400 574.050 891.450 595.950 ;
        RECT 892.950 592.950 895.050 595.050 ;
        RECT 893.400 574.050 894.450 592.950 ;
        RECT 899.400 589.050 900.450 634.950 ;
        RECT 908.400 621.450 909.450 649.950 ;
        RECT 911.400 637.050 912.450 655.950 ;
        RECT 917.400 655.050 918.450 658.950 ;
        RECT 916.950 652.950 919.050 655.050 ;
        RECT 913.950 651.600 918.000 652.050 ;
        RECT 913.950 649.950 918.600 651.600 ;
        RECT 922.950 651.000 925.050 655.050 ;
        RECT 917.400 649.350 918.600 649.950 ;
        RECT 923.400 649.350 924.600 651.000 ;
        RECT 916.950 646.950 919.050 649.050 ;
        RECT 919.950 646.950 922.050 649.050 ;
        RECT 922.950 646.950 925.050 649.050 ;
        RECT 913.950 643.950 916.050 646.050 ;
        RECT 920.400 644.400 921.600 646.650 ;
        RECT 910.950 634.950 913.050 637.050 ;
        RECT 911.400 631.050 912.450 634.950 ;
        RECT 910.950 628.950 913.050 631.050 ;
        RECT 910.950 621.450 913.050 622.050 ;
        RECT 908.400 620.400 913.050 621.450 ;
        RECT 910.950 619.950 913.050 620.400 ;
        RECT 901.950 616.950 904.050 619.050 ;
        RECT 902.400 601.050 903.450 616.950 ;
        RECT 911.400 606.600 912.450 619.950 ;
        RECT 914.400 610.050 915.450 643.950 ;
        RECT 920.400 643.050 921.450 644.400 ;
        RECT 925.950 643.950 928.050 646.050 ;
        RECT 920.400 640.950 925.050 643.050 ;
        RECT 916.950 628.950 919.050 631.050 ;
        RECT 917.400 613.050 918.450 628.950 ;
        RECT 920.400 625.050 921.450 640.950 ;
        RECT 925.950 637.950 928.050 640.050 ;
        RECT 922.950 634.950 925.050 637.050 ;
        RECT 919.950 622.950 922.050 625.050 ;
        RECT 916.950 610.950 919.050 613.050 ;
        RECT 913.950 607.950 916.050 610.050 ;
        RECT 911.400 604.350 912.600 606.600 ;
        RECT 916.950 605.100 919.050 607.200 ;
        RECT 917.400 604.350 918.600 605.100 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 916.950 601.950 919.050 604.050 ;
        RECT 901.950 598.950 904.050 601.050 ;
        RECT 908.400 600.900 909.600 601.650 ;
        RECT 907.950 598.800 910.050 600.900 ;
        RECT 914.400 599.400 915.600 601.650 ;
        RECT 898.950 586.950 901.050 589.050 ;
        RECT 895.950 583.950 898.050 586.050 ;
        RECT 887.400 571.350 888.600 573.000 ;
        RECT 889.950 571.950 892.050 574.050 ;
        RECT 892.950 571.950 895.050 574.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 892.950 568.800 895.050 570.900 ;
        RECT 878.400 567.450 879.600 568.650 ;
        RECT 884.400 567.900 885.600 568.650 ;
        RECT 875.400 566.400 879.600 567.450 ;
        RECT 871.950 562.950 874.050 565.050 ;
        RECT 871.950 553.950 874.050 556.050 ;
        RECT 872.400 541.050 873.450 553.950 ;
        RECT 871.950 538.950 874.050 541.050 ;
        RECT 871.950 532.950 874.050 535.050 ;
        RECT 868.950 529.950 871.050 532.050 ;
        RECT 872.400 528.600 873.450 532.950 ;
        RECT 875.400 532.050 876.450 566.400 ;
        RECT 883.950 565.800 886.050 567.900 ;
        RECT 893.400 565.050 894.450 568.800 ;
        RECT 877.950 562.950 880.050 565.050 ;
        RECT 892.950 562.950 895.050 565.050 ;
        RECT 878.400 550.050 879.450 562.950 ;
        RECT 893.400 559.050 894.450 562.950 ;
        RECT 892.950 556.950 895.050 559.050 ;
        RECT 877.950 547.950 880.050 550.050 ;
        RECT 886.950 541.950 889.050 544.050 ;
        RECT 877.950 535.950 880.050 538.050 ;
        RECT 874.950 529.950 877.050 532.050 ;
        RECT 878.400 528.600 879.450 535.950 ;
        RECT 887.400 535.050 888.450 541.950 ;
        RECT 886.950 532.950 889.050 535.050 ;
        RECT 889.950 532.950 892.050 535.050 ;
        RECT 872.400 526.350 873.600 528.600 ;
        RECT 878.400 526.350 879.600 528.600 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 875.400 522.900 876.600 523.650 ;
        RECT 874.950 520.800 877.050 522.900 ;
        RECT 880.950 519.450 883.050 522.900 ;
        RECT 878.400 519.000 883.050 519.450 ;
        RECT 878.400 518.400 882.450 519.000 ;
        RECT 865.950 508.950 868.050 511.050 ;
        RECT 862.950 505.950 865.050 508.050 ;
        RECT 857.400 497.400 861.450 498.450 ;
        RECT 857.400 495.600 858.450 497.400 ;
        RECT 857.400 493.350 858.600 495.600 ;
        RECT 862.950 494.100 865.050 496.200 ;
        RECT 863.400 493.350 864.600 494.100 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 853.950 487.950 856.050 490.050 ;
        RECT 860.400 488.400 861.600 490.650 ;
        RECT 850.950 484.950 853.050 487.050 ;
        RECT 854.400 481.050 855.450 487.950 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 853.800 478.950 855.900 481.050 ;
        RECT 856.950 478.950 859.050 481.050 ;
        RECT 850.950 469.950 853.050 472.050 ;
        RECT 847.950 421.950 850.050 424.050 ;
        RECT 851.400 420.450 852.450 469.950 ;
        RECT 853.950 466.950 856.050 469.050 ;
        RECT 854.400 454.050 855.450 466.950 ;
        RECT 857.400 460.050 858.450 478.950 ;
        RECT 860.400 469.050 861.450 488.400 ;
        RECT 868.800 487.950 870.900 490.050 ;
        RECT 874.800 487.950 876.900 490.050 ;
        RECT 869.400 485.400 870.600 487.650 ;
        RECT 865.950 475.950 868.050 478.050 ;
        RECT 866.400 469.050 867.450 475.950 ;
        RECT 859.950 466.950 862.050 469.050 ;
        RECT 865.950 466.950 868.050 469.050 ;
        RECT 859.950 460.950 862.050 463.050 ;
        RECT 856.950 457.950 859.050 460.050 ;
        RECT 860.400 457.050 861.450 460.950 ;
        RECT 859.950 454.950 862.050 457.050 ;
        RECT 865.950 456.450 868.050 457.050 ;
        RECT 869.400 456.450 870.450 485.400 ;
        RECT 878.400 484.050 879.450 518.400 ;
        RECT 890.400 517.050 891.450 532.950 ;
        RECT 896.400 532.050 897.450 583.950 ;
        RECT 908.400 580.050 909.450 598.800 ;
        RECT 914.400 597.450 915.450 599.400 ;
        RECT 919.950 597.450 922.050 598.050 ;
        RECT 914.400 596.400 922.050 597.450 ;
        RECT 919.950 595.950 922.050 596.400 ;
        RECT 916.950 592.950 919.050 595.050 ;
        RECT 917.400 583.050 918.450 592.950 ;
        RECT 919.950 586.950 922.050 589.050 ;
        RECT 916.950 580.950 919.050 583.050 ;
        RECT 898.950 577.950 901.050 580.050 ;
        RECT 907.950 577.950 910.050 580.050 ;
        RECT 899.400 562.050 900.450 577.950 ;
        RECT 907.950 572.100 910.050 574.200 ;
        RECT 913.950 573.000 916.050 577.050 ;
        RECT 908.400 571.350 909.600 572.100 ;
        RECT 914.400 571.350 915.600 573.000 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 913.950 568.950 916.050 571.050 ;
        RECT 905.400 567.000 906.600 568.650 ;
        RECT 911.400 567.000 912.600 568.650 ;
        RECT 920.400 568.050 921.450 586.950 ;
        RECT 904.950 562.950 907.050 567.000 ;
        RECT 910.950 562.950 913.050 567.000 ;
        RECT 916.950 565.950 919.050 568.050 ;
        RECT 919.950 565.950 922.050 568.050 ;
        RECT 913.950 562.950 916.050 565.050 ;
        RECT 898.950 559.950 901.050 562.050 ;
        RECT 898.950 556.800 901.050 558.900 ;
        RECT 899.400 550.050 900.450 556.800 ;
        RECT 914.400 556.050 915.450 562.950 ;
        RECT 917.400 559.050 918.450 565.950 ;
        RECT 923.400 565.050 924.450 634.950 ;
        RECT 926.400 607.050 927.450 637.950 ;
        RECT 929.400 628.050 930.450 670.950 ;
        RECT 932.400 670.050 933.450 673.950 ;
        RECT 931.950 667.950 934.050 670.050 ;
        RECT 935.400 667.050 936.450 677.400 ;
        RECT 943.950 676.800 946.050 678.900 ;
        RECT 946.950 676.950 949.050 679.050 ;
        RECT 940.950 667.950 943.050 670.050 ;
        RECT 944.400 669.450 945.450 676.800 ;
        RECT 947.400 673.050 948.450 676.950 ;
        RECT 946.950 670.950 949.050 673.050 ;
        RECT 944.400 668.400 948.450 669.450 ;
        RECT 934.950 664.950 937.050 667.050 ;
        RECT 941.400 661.050 942.450 667.950 ;
        RECT 947.400 661.050 948.450 668.400 ;
        RECT 934.950 658.950 937.050 661.050 ;
        RECT 940.950 658.950 943.050 661.050 ;
        RECT 946.950 658.950 949.050 661.050 ;
        RECT 931.950 649.950 934.050 655.050 ;
        RECT 932.400 646.050 933.450 649.950 ;
        RECT 931.950 643.950 934.050 646.050 ;
        RECT 931.950 640.800 934.050 642.900 ;
        RECT 928.950 625.950 931.050 628.050 ;
        RECT 932.400 619.050 933.450 640.800 ;
        RECT 935.400 631.050 936.450 658.950 ;
        RECT 943.950 655.950 946.050 658.050 ;
        RECT 944.400 651.600 945.450 655.950 ;
        RECT 950.400 652.050 951.450 703.950 ;
        RECT 953.400 691.050 954.450 721.800 ;
        RECT 955.950 700.950 958.050 703.050 ;
        RECT 952.950 688.950 955.050 691.050 ;
        RECT 952.950 683.100 955.050 685.200 ;
        RECT 953.400 676.050 954.450 683.100 ;
        RECT 956.400 678.900 957.450 700.950 ;
        RECT 955.950 676.800 958.050 678.900 ;
        RECT 952.950 673.950 955.050 676.050 ;
        RECT 952.950 670.800 955.050 672.900 ;
        RECT 944.400 649.350 945.600 651.600 ;
        RECT 949.950 649.950 952.050 652.050 ;
        RECT 940.950 646.950 943.050 649.050 ;
        RECT 943.950 646.950 946.050 649.050 ;
        RECT 946.950 646.950 949.050 649.050 ;
        RECT 941.400 645.000 942.600 646.650 ;
        RECT 947.400 645.900 948.600 646.650 ;
        RECT 953.400 646.050 954.450 670.800 ;
        RECT 940.950 640.950 943.050 645.000 ;
        RECT 946.950 640.950 949.050 645.900 ;
        RECT 952.950 643.950 955.050 646.050 ;
        RECT 952.950 640.800 955.050 642.900 ;
        RECT 940.950 637.800 943.050 639.900 ;
        RECT 946.950 637.800 949.050 639.900 ;
        RECT 934.950 628.950 937.050 631.050 ;
        RECT 931.950 618.450 934.050 619.050 ;
        RECT 929.400 617.400 934.050 618.450 ;
        RECT 925.950 604.950 928.050 607.050 ;
        RECT 925.950 601.800 928.050 603.900 ;
        RECT 926.400 598.050 927.450 601.800 ;
        RECT 925.950 595.950 928.050 598.050 ;
        RECT 926.400 589.050 927.450 595.950 ;
        RECT 925.950 586.950 928.050 589.050 ;
        RECT 925.950 580.950 928.050 583.050 ;
        RECT 926.400 577.050 927.450 580.950 ;
        RECT 925.950 574.950 928.050 577.050 ;
        RECT 929.400 574.050 930.450 617.400 ;
        RECT 931.950 616.950 934.050 617.400 ;
        RECT 947.400 615.450 948.450 637.800 ;
        RECT 949.950 625.950 952.050 628.050 ;
        RECT 944.400 614.400 948.450 615.450 ;
        RECT 934.950 609.450 937.050 613.050 ;
        RECT 934.950 609.000 942.450 609.450 ;
        RECT 935.400 608.400 942.450 609.000 ;
        RECT 934.950 605.100 937.050 607.200 ;
        RECT 941.400 606.600 942.450 608.400 ;
        RECT 944.400 607.050 945.450 614.400 ;
        RECT 946.950 610.950 949.050 613.050 ;
        RECT 935.400 604.350 936.600 605.100 ;
        RECT 941.400 604.350 942.600 606.600 ;
        RECT 943.950 604.950 946.050 607.050 ;
        RECT 934.950 601.950 937.050 604.050 ;
        RECT 937.950 601.950 940.050 604.050 ;
        RECT 940.950 601.950 943.050 604.050 ;
        RECT 931.950 598.950 934.050 601.050 ;
        RECT 938.400 599.400 939.600 601.650 ;
        RECT 932.400 577.050 933.450 598.950 ;
        RECT 938.400 595.050 939.450 599.400 ;
        RECT 943.950 598.950 946.050 601.050 ;
        RECT 937.950 592.950 940.050 595.050 ;
        RECT 940.950 591.450 943.050 592.050 ;
        RECT 935.400 590.400 943.050 591.450 ;
        RECT 935.400 583.050 936.450 590.400 ;
        RECT 940.950 589.950 943.050 590.400 ;
        RECT 937.950 586.950 940.050 589.050 ;
        RECT 934.950 580.950 937.050 583.050 ;
        RECT 938.400 579.450 939.450 586.950 ;
        RECT 940.950 580.950 943.050 583.050 ;
        RECT 935.400 578.400 939.450 579.450 ;
        RECT 931.950 574.950 934.050 577.050 ;
        RECT 925.950 571.800 928.050 573.900 ;
        RECT 928.950 571.950 931.050 574.050 ;
        RECT 935.400 573.600 936.450 578.400 ;
        RECT 941.400 573.600 942.450 580.950 ;
        RECT 944.400 574.050 945.450 598.950 ;
        RECT 922.950 562.950 925.050 565.050 ;
        RECT 916.950 556.950 919.050 559.050 ;
        RECT 913.950 553.950 916.050 556.050 ;
        RECT 926.400 553.050 927.450 571.800 ;
        RECT 935.400 571.350 936.600 573.600 ;
        RECT 941.400 571.350 942.600 573.600 ;
        RECT 943.950 571.950 946.050 574.050 ;
        RECT 931.950 568.950 934.050 571.050 ;
        RECT 934.950 568.950 937.050 571.050 ;
        RECT 937.950 568.950 940.050 571.050 ;
        RECT 940.950 568.950 943.050 571.050 ;
        RECT 928.950 565.950 931.050 568.050 ;
        RECT 932.400 567.000 933.600 568.650 ;
        RECT 938.400 567.900 939.600 568.650 ;
        RECT 929.400 553.050 930.450 565.950 ;
        RECT 931.950 562.950 934.050 567.000 ;
        RECT 937.950 565.800 940.050 567.900 ;
        RECT 934.950 562.950 937.050 565.050 ;
        RECT 931.950 556.950 934.050 561.900 ;
        RECT 919.950 550.950 922.050 553.050 ;
        RECT 925.800 550.950 927.900 553.050 ;
        RECT 928.950 550.950 931.050 553.050 ;
        RECT 898.950 547.950 901.050 550.050 ;
        RECT 913.950 547.950 916.050 550.050 ;
        RECT 910.950 538.950 913.050 541.050 ;
        RECT 911.400 535.050 912.450 538.950 ;
        RECT 901.950 532.950 904.050 535.050 ;
        RECT 910.950 532.950 913.050 535.050 ;
        RECT 895.950 529.950 898.050 532.050 ;
        RECT 901.950 527.100 904.050 529.200 ;
        RECT 910.950 527.100 913.050 529.200 ;
        RECT 902.400 526.350 903.600 527.100 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 899.400 522.900 900.600 523.650 ;
        RECT 898.950 520.800 901.050 522.900 ;
        RECT 905.400 521.400 906.600 523.650 ;
        RECT 911.400 523.050 912.450 527.100 ;
        RECT 889.950 514.950 892.050 517.050 ;
        RECT 905.400 508.050 906.450 521.400 ;
        RECT 910.950 520.950 913.050 523.050 ;
        RECT 914.400 514.050 915.450 547.950 ;
        RECT 916.950 538.950 919.050 541.050 ;
        RECT 920.400 534.450 921.450 550.950 ;
        RECT 922.950 538.950 925.050 541.050 ;
        RECT 917.400 533.400 921.450 534.450 ;
        RECT 913.950 511.950 916.050 514.050 ;
        RECT 904.950 505.950 907.050 508.050 ;
        RECT 913.950 505.950 916.050 508.050 ;
        RECT 881.700 501.300 883.800 503.400 ;
        RECT 884.700 501.300 886.800 503.400 ;
        RECT 887.700 501.300 889.800 503.400 ;
        RECT 882.300 497.700 883.500 501.300 ;
        RECT 881.400 495.600 883.500 497.700 ;
        RECT 877.950 481.950 880.050 484.050 ;
        RECT 874.950 475.950 877.050 478.050 ;
        RECT 881.400 476.700 882.900 495.600 ;
        RECT 885.300 484.800 886.500 501.300 ;
        RECT 884.400 482.700 886.500 484.800 ;
        RECT 885.300 476.700 886.500 482.700 ;
        RECT 887.700 479.700 888.900 501.300 ;
        RECT 895.800 500.400 897.900 502.500 ;
        RECT 901.200 501.300 903.300 503.400 ;
        RECT 904.200 501.300 906.300 503.400 ;
        RECT 907.200 501.300 909.300 503.400 ;
        RECT 892.800 493.950 894.900 496.050 ;
        RECT 893.400 491.400 894.600 493.650 ;
        RECT 887.700 477.600 889.800 479.700 ;
        RECT 893.400 478.050 894.450 491.400 ;
        RECT 896.400 489.900 897.300 500.400 ;
        RECT 899.100 494.400 901.200 496.500 ;
        RECT 896.400 487.800 898.500 489.900 ;
        RECT 902.100 489.000 903.300 501.300 ;
        RECT 896.400 481.200 897.300 487.800 ;
        RECT 901.800 486.900 903.900 489.000 ;
        RECT 896.400 479.100 898.500 481.200 ;
        RECT 902.100 479.700 903.300 486.900 ;
        RECT 904.800 483.600 906.300 501.300 ;
        RECT 904.800 481.500 906.900 483.600 ;
        RECT 865.950 455.400 870.450 456.450 ;
        RECT 853.950 451.950 856.050 454.050 ;
        RECT 860.400 450.600 861.450 454.950 ;
        RECT 865.950 453.000 868.050 455.400 ;
        RECT 866.400 451.350 867.600 453.000 ;
        RECT 860.400 448.350 861.600 450.600 ;
        RECT 865.800 448.950 867.900 451.050 ;
        RECT 871.800 448.950 873.900 451.050 ;
        RECT 854.400 445.950 856.500 448.050 ;
        RECT 859.800 445.950 861.900 448.050 ;
        RECT 868.950 445.950 871.050 448.050 ;
        RECT 854.400 443.400 855.600 445.650 ;
        RECT 854.400 439.050 855.450 443.400 ;
        RECT 853.950 436.950 856.050 439.050 ;
        RECT 869.400 433.050 870.450 445.950 ;
        RECT 868.950 430.950 871.050 433.050 ;
        RECT 871.950 421.800 874.050 423.900 ;
        RECT 848.400 419.400 852.450 420.450 ;
        RECT 848.400 409.050 849.450 419.400 ;
        RECT 853.950 416.100 856.050 418.200 ;
        RECT 862.950 417.000 865.050 421.050 ;
        RECT 854.400 415.350 855.600 416.100 ;
        RECT 863.400 415.350 864.600 417.000 ;
        RECT 851.100 412.950 853.200 415.050 ;
        RECT 854.100 412.950 856.200 415.050 ;
        RECT 859.800 412.950 861.900 415.050 ;
        RECT 862.800 412.950 864.900 415.050 ;
        RECT 851.400 411.000 852.600 412.650 ;
        RECT 847.950 406.950 850.050 409.050 ;
        RECT 850.950 406.950 853.050 411.000 ;
        RECT 860.400 410.400 861.600 412.650 ;
        RECT 860.400 390.450 861.450 410.400 ;
        RECT 872.400 403.050 873.450 421.800 ;
        RECT 871.950 400.950 874.050 403.050 ;
        RECT 875.400 400.050 876.450 475.950 ;
        RECT 881.400 474.600 884.400 476.700 ;
        RECT 885.300 474.600 887.400 476.700 ;
        RECT 892.950 475.950 895.050 478.050 ;
        RECT 901.800 477.600 903.900 479.700 ;
        RECT 904.800 476.700 906.300 481.500 ;
        RECT 908.100 479.700 909.300 501.300 ;
        RECT 904.200 474.600 906.300 476.700 ;
        RECT 907.200 474.600 909.300 479.700 ;
        RECT 910.200 501.300 912.300 503.400 ;
        RECT 910.200 483.600 911.700 501.300 ;
        RECT 914.400 496.050 915.450 505.950 ;
        RECT 917.400 502.050 918.450 533.400 ;
        RECT 919.950 526.950 922.050 532.050 ;
        RECT 923.400 531.450 924.450 538.950 ;
        RECT 935.400 534.450 936.450 562.950 ;
        RECT 938.400 538.050 939.450 565.800 ;
        RECT 940.950 553.950 943.050 556.050 ;
        RECT 937.950 535.950 940.050 538.050 ;
        RECT 935.400 533.400 939.450 534.450 ;
        RECT 923.400 530.400 927.450 531.450 ;
        RECT 926.400 528.600 927.450 530.400 ;
        RECT 926.400 526.350 927.600 528.600 ;
        RECT 931.950 528.000 934.050 532.050 ;
        RECT 932.400 526.350 933.600 528.000 ;
        RECT 922.950 523.950 925.050 526.050 ;
        RECT 925.950 523.950 928.050 526.050 ;
        RECT 928.950 523.950 931.050 526.050 ;
        RECT 931.950 523.950 934.050 526.050 ;
        RECT 919.950 520.950 922.050 523.050 ;
        RECT 923.400 522.900 924.600 523.650 ;
        RECT 929.400 522.900 930.600 523.650 ;
        RECT 916.950 499.950 919.050 502.050 ;
        RECT 920.400 499.050 921.450 520.950 ;
        RECT 922.950 520.800 925.050 522.900 ;
        RECT 928.950 520.800 931.050 522.900 ;
        RECT 934.950 520.800 937.050 523.050 ;
        RECT 922.950 514.950 925.050 517.050 ;
        RECT 919.950 496.950 922.050 499.050 ;
        RECT 913.950 493.950 916.050 496.050 ;
        RECT 913.950 490.800 916.050 492.900 ;
        RECT 919.950 491.100 922.050 493.200 ;
        RECT 910.200 481.500 912.300 483.600 ;
        RECT 914.400 483.450 915.450 490.800 ;
        RECT 920.400 490.350 921.600 491.100 ;
        RECT 919.800 487.950 921.900 490.050 ;
        RECT 914.400 482.400 918.450 483.450 ;
        RECT 910.200 476.700 911.700 481.500 ;
        RECT 913.950 478.950 916.050 481.050 ;
        RECT 910.200 474.600 912.300 476.700 ;
        RECT 914.400 472.050 915.450 478.950 ;
        RECT 913.950 469.950 916.050 472.050 ;
        RECT 878.400 462.300 881.400 464.400 ;
        RECT 882.300 462.300 884.400 464.400 ;
        RECT 889.950 463.950 892.050 466.050 ;
        RECT 878.400 443.400 879.900 462.300 ;
        RECT 882.300 456.300 883.500 462.300 ;
        RECT 881.400 454.200 883.500 456.300 ;
        RECT 878.400 441.300 880.500 443.400 ;
        RECT 879.300 437.700 880.500 441.300 ;
        RECT 882.300 437.700 883.500 454.200 ;
        RECT 884.700 459.300 886.800 461.400 ;
        RECT 884.700 437.700 885.900 459.300 ;
        RECT 890.400 453.450 891.450 463.950 ;
        RECT 901.200 462.300 903.300 464.400 ;
        RECT 887.400 452.400 891.450 453.450 ;
        RECT 893.400 457.800 895.500 459.900 ;
        RECT 898.800 459.300 900.900 461.400 ;
        RECT 887.400 448.050 888.450 452.400 ;
        RECT 893.400 451.200 894.300 457.800 ;
        RECT 899.100 452.100 900.300 459.300 ;
        RECT 901.800 457.500 903.300 462.300 ;
        RECT 904.200 459.300 906.300 464.400 ;
        RECT 901.800 455.400 903.900 457.500 ;
        RECT 893.400 449.100 895.500 451.200 ;
        RECT 898.800 450.000 900.900 452.100 ;
        RECT 886.800 445.950 888.900 448.050 ;
        RECT 889.950 446.100 892.050 448.200 ;
        RECT 890.400 445.350 891.600 446.100 ;
        RECT 889.800 442.950 891.900 445.050 ;
        RECT 893.400 438.600 894.300 449.100 ;
        RECT 896.100 442.500 898.200 444.600 ;
        RECT 878.700 435.600 880.800 437.700 ;
        RECT 881.700 435.600 883.800 437.700 ;
        RECT 884.700 435.600 886.800 437.700 ;
        RECT 892.800 436.500 894.900 438.600 ;
        RECT 899.100 437.700 900.300 450.000 ;
        RECT 901.800 437.700 903.300 455.400 ;
        RECT 905.100 437.700 906.300 459.300 ;
        RECT 898.200 435.600 900.300 437.700 ;
        RECT 901.200 435.600 903.300 437.700 ;
        RECT 904.200 435.600 906.300 437.700 ;
        RECT 907.200 462.300 909.300 464.400 ;
        RECT 917.400 463.050 918.450 482.400 ;
        RECT 919.950 481.950 922.050 484.050 ;
        RECT 920.400 475.050 921.450 481.950 ;
        RECT 919.950 472.950 922.050 475.050 ;
        RECT 923.400 471.450 924.450 514.950 ;
        RECT 931.950 511.950 934.050 514.050 ;
        RECT 925.950 492.600 930.000 493.050 ;
        RECT 925.950 490.950 930.600 492.600 ;
        RECT 929.400 490.350 930.600 490.950 ;
        RECT 928.800 487.950 930.900 490.050 ;
        RECT 925.950 483.450 928.050 487.050 ;
        RECT 925.950 483.000 930.450 483.450 ;
        RECT 926.400 482.400 930.450 483.000 ;
        RECT 929.400 472.050 930.450 482.400 ;
        RECT 923.400 470.400 927.450 471.450 ;
        RECT 919.950 466.950 922.050 469.050 ;
        RECT 920.400 463.050 921.450 466.950 ;
        RECT 907.200 457.500 908.700 462.300 ;
        RECT 910.950 460.950 913.050 463.050 ;
        RECT 916.800 460.950 918.900 463.050 ;
        RECT 919.950 460.950 922.050 463.050 ;
        RECT 907.200 455.400 909.300 457.500 ;
        RECT 907.200 437.700 908.700 455.400 ;
        RECT 911.400 447.900 912.450 460.950 ;
        RECT 919.950 454.950 922.050 457.050 ;
        RECT 926.400 456.450 927.450 470.400 ;
        RECT 928.950 469.950 931.050 472.050 ;
        RECT 926.400 455.400 930.450 456.450 ;
        RECT 916.800 448.950 918.900 451.050 ;
        RECT 917.400 447.900 918.600 448.650 ;
        RECT 910.950 445.800 913.050 447.900 ;
        RECT 916.950 445.800 919.050 447.900 ;
        RECT 907.200 435.600 909.300 437.700 ;
        RECT 910.950 436.950 913.050 439.050 ;
        RECT 883.950 430.950 886.050 433.050 ;
        RECT 895.950 430.950 898.050 433.050 ;
        RECT 884.400 417.600 885.450 430.950 ;
        RECT 892.950 421.950 895.050 424.050 ;
        RECT 893.400 417.600 894.450 421.950 ;
        RECT 884.400 415.350 885.600 417.600 ;
        RECT 893.400 415.350 894.600 417.600 ;
        RECT 881.100 412.950 883.200 415.050 ;
        RECT 884.100 412.950 886.200 415.050 ;
        RECT 889.800 412.950 891.900 415.050 ;
        RECT 892.800 412.950 894.900 415.050 ;
        RECT 881.400 410.400 882.600 412.650 ;
        RECT 890.400 411.900 891.600 412.650 ;
        RECT 896.400 412.050 897.450 430.950 ;
        RECT 911.400 427.050 912.450 436.950 ;
        RECT 920.400 430.050 921.450 454.950 ;
        RECT 925.800 448.950 927.900 451.050 ;
        RECT 926.400 446.400 927.600 448.650 ;
        RECT 926.400 442.050 927.450 446.400 ;
        RECT 925.950 439.950 928.050 442.050 ;
        RECT 922.950 438.450 925.050 439.050 ;
        RECT 929.400 438.450 930.450 455.400 ;
        RECT 922.950 437.400 930.450 438.450 ;
        RECT 922.950 436.950 925.050 437.400 ;
        RECT 928.950 433.950 931.050 436.050 ;
        RECT 919.950 427.950 922.050 430.050 ;
        RECT 904.950 424.950 907.050 427.050 ;
        RECT 910.950 424.950 913.050 427.050 ;
        RECT 929.400 426.450 930.450 433.950 ;
        RECT 926.400 425.400 930.450 426.450 ;
        RECT 881.400 409.050 882.450 410.400 ;
        RECT 889.950 409.800 892.050 411.900 ;
        RECT 895.950 409.950 898.050 412.050 ;
        RECT 880.950 406.950 883.050 409.050 ;
        RECT 874.950 397.950 877.050 400.050 ;
        RECT 881.400 391.050 882.450 406.950 ;
        RECT 889.800 397.950 891.900 400.050 ;
        RECT 892.950 397.950 895.050 400.050 ;
        RECT 860.400 389.400 864.450 390.450 ;
        RECT 848.400 384.300 851.400 386.400 ;
        RECT 852.300 384.300 854.400 386.400 ;
        RECT 859.950 385.950 862.050 388.050 ;
        RECT 844.950 376.950 847.050 379.050 ;
        RECT 823.800 373.950 825.900 376.050 ;
        RECT 826.950 374.100 829.050 376.200 ;
        RECT 835.950 374.100 838.050 376.200 ;
        RECT 827.400 373.350 828.600 374.100 ;
        RECT 836.400 373.350 837.600 374.100 ;
        RECT 844.950 373.800 847.050 375.900 ;
        RECT 821.100 370.950 823.200 373.050 ;
        RECT 827.100 370.950 829.200 373.050 ;
        RECT 835.800 370.950 837.900 373.050 ;
        RECT 841.800 370.950 843.900 373.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 820.950 364.950 823.050 367.050 ;
        RECT 817.950 346.950 820.050 349.050 ;
        RECT 799.950 343.950 802.050 346.050 ;
        RECT 778.950 338.100 781.050 340.200 ;
        RECT 775.950 310.950 778.050 313.050 ;
        RECT 779.400 304.050 780.450 338.100 ;
        RECT 781.950 337.950 784.050 340.050 ;
        RECT 787.950 338.100 790.050 340.200 ;
        RECT 793.950 338.100 796.050 340.200 ;
        RECT 800.400 339.450 801.450 343.950 ;
        RECT 821.400 343.050 822.450 364.950 ;
        RECT 826.950 361.950 829.050 364.050 ;
        RECT 823.950 346.950 826.050 349.050 ;
        RECT 811.950 340.950 814.050 343.050 ;
        RECT 820.950 340.950 823.050 343.050 ;
        RECT 800.400 338.400 804.450 339.450 ;
        RECT 782.400 333.900 783.450 337.950 ;
        RECT 788.400 337.350 789.600 338.100 ;
        RECT 794.400 337.350 795.600 338.100 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 791.400 333.900 792.600 334.650 ;
        RECT 797.400 333.900 798.600 334.650 ;
        RECT 803.400 333.900 804.450 338.400 ;
        RECT 805.950 337.950 808.050 340.050 ;
        RECT 781.950 331.800 784.050 333.900 ;
        RECT 790.950 331.800 793.050 333.900 ;
        RECT 796.950 331.800 799.050 333.900 ;
        RECT 802.950 331.800 805.050 333.900 ;
        RECT 802.950 319.950 805.050 322.050 ;
        RECT 760.950 301.950 763.050 304.050 ;
        RECT 766.950 301.950 769.050 304.050 ;
        RECT 778.950 301.950 781.050 304.050 ;
        RECT 772.950 298.950 775.050 301.050 ;
        RECT 757.800 292.950 759.900 295.050 ;
        RECT 760.950 293.100 763.050 298.050 ;
        RECT 766.950 294.000 769.050 298.050 ;
        RECT 761.400 292.350 762.600 293.100 ;
        RECT 767.400 292.350 768.600 294.000 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 757.950 286.950 760.050 289.050 ;
        RECT 764.400 288.900 765.600 289.650 ;
        RECT 758.400 274.050 759.450 286.950 ;
        RECT 763.950 286.800 766.050 288.900 ;
        RECT 766.950 283.950 769.050 286.050 ;
        RECT 757.950 271.950 760.050 274.050 ;
        RECT 767.400 267.450 768.450 283.950 ;
        RECT 773.400 271.050 774.450 298.950 ;
        RECT 775.950 295.950 778.050 298.050 ;
        RECT 776.400 292.050 777.450 295.950 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 776.400 286.050 777.450 289.950 ;
        RECT 775.950 283.950 778.050 286.050 ;
        RECT 779.400 285.450 780.450 301.950 ;
        RECT 788.100 298.500 790.200 300.600 ;
        RECT 781.950 292.950 784.050 295.050 ;
        RECT 782.400 288.450 783.450 292.950 ;
        RECT 785.100 289.950 787.200 292.050 ;
        RECT 788.100 291.900 789.000 298.500 ;
        RECT 797.100 298.200 799.200 300.300 ;
        RECT 791.400 295.350 792.600 297.600 ;
        RECT 790.800 292.950 792.900 295.050 ;
        RECT 795.000 291.900 797.100 292.200 ;
        RECT 788.100 291.000 797.100 291.900 ;
        RECT 785.400 288.450 786.600 289.650 ;
        RECT 782.400 287.400 786.600 288.450 ;
        RECT 788.100 285.900 789.000 291.000 ;
        RECT 795.000 290.100 797.100 291.000 ;
        RECT 789.900 289.200 792.000 290.100 ;
        RECT 789.900 288.000 797.100 289.200 ;
        RECT 795.000 287.100 797.100 288.000 ;
        RECT 779.400 284.400 783.450 285.450 ;
        RECT 778.950 274.950 781.050 277.050 ;
        RECT 775.950 271.950 778.050 274.050 ;
        RECT 772.950 268.950 775.050 271.050 ;
        RECT 767.400 265.200 768.600 267.450 ;
        RECT 762.900 261.900 765.000 263.700 ;
        RECT 766.800 262.800 768.900 264.900 ;
        RECT 770.100 264.300 772.200 266.400 ;
        RECT 761.400 260.700 770.100 261.900 ;
        RECT 758.100 256.950 760.200 259.050 ;
        RECT 758.400 255.450 759.600 256.650 ;
        RECT 755.400 254.400 759.600 255.450 ;
        RECT 761.400 251.700 762.300 260.700 ;
        RECT 768.000 259.800 770.100 260.700 ;
        RECT 771.000 258.900 771.900 264.300 ;
        RECT 772.950 260.100 775.050 262.200 ;
        RECT 773.400 259.350 774.600 260.100 ;
        RECT 765.000 257.700 771.900 258.900 ;
        RECT 765.000 255.300 765.900 257.700 ;
        RECT 763.800 253.200 765.900 255.300 ;
        RECT 766.800 253.950 768.900 256.050 ;
        RECT 760.500 249.600 762.600 251.700 ;
        RECT 767.400 251.400 768.600 253.650 ;
        RECT 770.700 250.500 771.900 257.700 ;
        RECT 772.800 256.950 774.900 259.050 ;
        RECT 770.100 248.400 772.200 250.500 ;
        RECT 766.950 229.950 769.050 232.050 ;
        RECT 737.400 214.350 738.600 215.100 ;
        RECT 745.950 214.950 748.050 217.050 ;
        RECT 751.950 214.950 754.050 217.050 ;
        RECT 760.950 215.100 763.050 217.200 ;
        RECT 767.400 216.600 768.450 229.950 ;
        RECT 776.400 220.050 777.450 271.950 ;
        RECT 775.950 217.950 778.050 220.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 740.400 210.900 741.600 211.650 ;
        RECT 746.400 210.900 747.450 214.950 ;
        RECT 761.400 214.350 762.600 215.100 ;
        RECT 767.400 214.350 768.600 216.600 ;
        RECT 773.100 214.950 775.200 217.050 ;
        RECT 751.950 211.800 754.050 213.900 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 773.400 213.900 774.600 214.650 ;
        RECT 772.950 211.800 775.050 213.900 ;
        RECT 779.400 213.450 780.450 274.950 ;
        RECT 782.400 256.050 783.450 284.400 ;
        RECT 787.500 283.800 789.600 285.900 ;
        RECT 790.800 284.100 792.900 286.200 ;
        RECT 798.000 285.600 798.900 298.200 ;
        RECT 799.950 293.100 802.050 295.200 ;
        RECT 800.400 292.350 801.600 293.100 ;
        RECT 799.800 289.950 801.900 292.050 ;
        RECT 791.400 283.050 792.600 283.800 ;
        RECT 797.400 283.500 799.500 285.600 ;
        RECT 790.950 280.950 793.050 283.050 ;
        RECT 799.950 268.950 802.050 271.050 ;
        RECT 784.950 259.950 787.050 262.050 ;
        RECT 790.950 260.100 793.050 262.200 ;
        RECT 781.950 253.950 784.050 256.050 ;
        RECT 785.400 231.450 786.450 259.950 ;
        RECT 791.400 259.350 792.600 260.100 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 794.400 255.900 795.600 256.650 ;
        RECT 793.950 253.800 796.050 255.900 ;
        RECT 800.400 238.050 801.450 268.950 ;
        RECT 799.950 235.950 802.050 238.050 ;
        RECT 803.400 232.050 804.450 319.950 ;
        RECT 806.400 301.050 807.450 337.950 ;
        RECT 808.950 304.950 811.050 307.050 ;
        RECT 805.950 298.950 808.050 301.050 ;
        RECT 809.400 298.050 810.450 304.950 ;
        RECT 808.950 295.950 811.050 298.050 ;
        RECT 806.100 292.950 808.200 295.050 ;
        RECT 806.400 291.900 807.600 292.650 ;
        RECT 805.950 289.800 808.050 291.900 ;
        RECT 805.950 268.950 808.050 271.050 ;
        RECT 806.400 250.050 807.450 268.950 ;
        RECT 812.400 268.050 813.450 340.950 ;
        RECT 821.400 339.450 822.600 339.600 ;
        RECT 824.400 339.450 825.450 346.950 ;
        RECT 821.400 338.400 825.450 339.450 ;
        RECT 821.400 337.350 822.600 338.400 ;
        RECT 815.100 334.950 817.200 337.050 ;
        RECT 820.500 334.950 822.600 337.050 ;
        RECT 815.400 333.900 816.600 334.650 ;
        RECT 814.950 331.800 817.050 333.900 ;
        RECT 815.400 300.450 816.450 331.800 ;
        RECT 824.400 325.050 825.450 338.400 ;
        RECT 827.400 334.050 828.450 361.950 ;
        RECT 826.950 331.950 829.050 334.050 ;
        RECT 826.950 325.950 829.050 328.050 ;
        RECT 823.950 322.950 826.050 325.050 ;
        RECT 823.950 316.950 826.050 319.050 ;
        RECT 827.400 316.050 828.450 325.950 ;
        RECT 833.400 322.050 834.450 367.950 ;
        RECT 845.400 367.050 846.450 373.800 ;
        RECT 844.950 364.950 847.050 367.050 ;
        RECT 848.400 365.400 849.900 384.300 ;
        RECT 852.300 378.300 853.500 384.300 ;
        RECT 851.400 376.200 853.500 378.300 ;
        RECT 848.400 363.300 850.500 365.400 ;
        RECT 844.950 358.950 847.050 361.050 ;
        RECT 849.300 359.700 850.500 363.300 ;
        RECT 852.300 359.700 853.500 376.200 ;
        RECT 854.700 381.300 856.800 383.400 ;
        RECT 854.700 359.700 855.900 381.300 ;
        RECT 856.950 376.950 859.050 379.050 ;
        RECT 857.400 370.050 858.450 376.950 ;
        RECT 860.400 376.050 861.450 385.950 ;
        RECT 863.400 385.050 864.450 389.400 ;
        RECT 880.950 388.950 883.050 391.050 ;
        RECT 862.950 382.950 865.050 385.050 ;
        RECT 871.200 384.300 873.300 386.400 ;
        RECT 863.400 379.800 865.500 381.900 ;
        RECT 868.800 381.300 870.900 383.400 ;
        RECT 859.950 373.950 862.050 376.050 ;
        RECT 863.400 373.200 864.300 379.800 ;
        RECT 869.100 374.100 870.300 381.300 ;
        RECT 871.800 379.500 873.300 384.300 ;
        RECT 874.200 381.300 876.300 386.400 ;
        RECT 871.800 377.400 873.900 379.500 ;
        RECT 863.400 371.100 865.500 373.200 ;
        RECT 868.800 372.000 870.900 374.100 ;
        RECT 856.800 367.950 858.900 370.050 ;
        RECT 859.950 368.100 862.050 370.200 ;
        RECT 860.400 367.350 861.600 368.100 ;
        RECT 859.800 364.950 861.900 367.050 ;
        RECT 863.400 360.600 864.300 371.100 ;
        RECT 866.100 364.500 868.200 366.600 ;
        RECT 845.400 352.050 846.450 358.950 ;
        RECT 848.700 357.600 850.800 359.700 ;
        RECT 851.700 357.600 853.800 359.700 ;
        RECT 854.700 357.600 856.800 359.700 ;
        RECT 862.800 358.500 864.900 360.600 ;
        RECT 869.100 359.700 870.300 372.000 ;
        RECT 871.800 359.700 873.300 377.400 ;
        RECT 875.100 359.700 876.300 381.300 ;
        RECT 868.200 357.600 870.300 359.700 ;
        RECT 871.200 357.600 873.300 359.700 ;
        RECT 874.200 357.600 876.300 359.700 ;
        RECT 877.200 384.300 879.300 386.400 ;
        RECT 877.200 379.500 878.700 384.300 ;
        RECT 880.950 382.950 883.050 385.050 ;
        RECT 877.200 377.400 879.300 379.500 ;
        RECT 877.200 359.700 878.700 377.400 ;
        RECT 881.400 370.200 882.450 382.950 ;
        RECT 886.800 370.950 888.900 373.050 ;
        RECT 880.950 368.100 883.050 370.200 ;
        RECT 887.400 368.400 888.600 370.650 ;
        RECT 890.400 369.450 891.450 397.950 ;
        RECT 893.400 394.050 894.450 397.950 ;
        RECT 892.950 391.950 895.050 394.050 ;
        RECT 895.800 370.950 897.900 373.050 ;
        RECT 896.400 369.450 897.600 370.650 ;
        RECT 898.950 369.450 901.050 373.050 ;
        RECT 901.950 370.950 904.050 373.050 ;
        RECT 890.400 368.400 894.450 369.450 ;
        RECT 896.400 369.000 901.050 369.450 ;
        RECT 896.400 368.400 900.450 369.000 ;
        RECT 887.400 361.050 888.450 368.400 ;
        RECT 889.950 364.950 892.050 367.050 ;
        RECT 886.950 360.450 889.050 361.050 ;
        RECT 877.200 357.600 879.300 359.700 ;
        RECT 884.400 359.400 889.050 360.450 ;
        RECT 853.950 352.950 856.050 355.050 ;
        RECT 844.950 349.950 847.050 352.050 ;
        RECT 844.950 342.450 847.050 346.050 ;
        RECT 842.400 342.000 847.050 342.450 ;
        RECT 842.400 341.400 846.450 342.000 ;
        RECT 842.400 339.600 843.450 341.400 ;
        RECT 842.400 337.350 843.600 339.600 ;
        RECT 847.950 338.100 850.050 340.200 ;
        RECT 848.400 337.350 849.600 338.100 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 839.400 332.400 840.600 334.650 ;
        RECT 845.400 333.000 846.600 334.650 ;
        RECT 835.950 322.950 838.050 325.050 ;
        RECT 832.950 319.950 835.050 322.050 ;
        RECT 836.400 319.050 837.450 322.950 ;
        RECT 835.950 316.950 838.050 319.050 ;
        RECT 826.800 313.950 828.900 316.050 ;
        RECT 839.400 310.050 840.450 332.400 ;
        RECT 844.950 328.950 847.050 333.000 ;
        RECT 854.400 325.050 855.450 352.950 ;
        RECT 856.950 349.950 859.050 352.050 ;
        RECT 857.400 328.050 858.450 349.950 ;
        RECT 880.950 346.950 883.050 349.050 ;
        RECT 859.950 337.950 862.050 340.050 ;
        RECT 865.950 338.100 868.050 340.200 ;
        RECT 871.950 338.100 874.050 340.200 ;
        RECT 860.400 331.050 861.450 337.950 ;
        RECT 866.400 337.350 867.600 338.100 ;
        RECT 872.400 337.350 873.600 338.100 ;
        RECT 865.950 334.950 868.050 337.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 862.950 331.950 865.050 334.050 ;
        RECT 869.400 333.000 870.600 334.650 ;
        RECT 859.950 328.950 862.050 331.050 ;
        RECT 856.950 325.950 859.050 328.050 ;
        RECT 853.950 322.950 856.050 325.050 ;
        RECT 841.950 316.950 844.050 319.050 ;
        RECT 842.400 313.050 843.450 316.950 ;
        RECT 863.400 313.050 864.450 331.950 ;
        RECT 868.950 328.950 871.050 333.000 ;
        RECT 875.400 332.400 876.600 334.650 ;
        RECT 875.400 325.050 876.450 332.400 ;
        RECT 877.950 331.950 880.050 334.050 ;
        RECT 874.950 322.950 877.050 325.050 ;
        RECT 871.950 313.950 874.050 316.050 ;
        RECT 841.950 310.950 844.050 313.050 ;
        RECT 862.950 310.950 865.050 313.050 ;
        RECT 824.700 306.300 826.800 308.400 ;
        RECT 825.300 301.500 826.800 306.300 ;
        RECT 815.400 300.000 819.450 300.450 ;
        RECT 815.400 299.400 820.050 300.000 ;
        RECT 824.700 299.400 826.800 301.500 ;
        RECT 817.950 297.450 820.050 299.400 ;
        RECT 817.950 296.400 822.450 297.450 ;
        RECT 817.950 296.100 820.050 296.400 ;
        RECT 815.100 292.950 817.200 295.050 ;
        RECT 815.400 290.400 816.600 292.650 ;
        RECT 815.400 277.050 816.450 290.400 ;
        RECT 814.950 274.950 817.050 277.050 ;
        RECT 821.400 271.050 822.450 296.400 ;
        RECT 825.300 281.700 826.800 299.400 ;
        RECT 824.700 279.600 826.800 281.700 ;
        RECT 827.700 303.300 829.800 308.400 ;
        RECT 830.700 306.300 832.800 308.400 ;
        RECT 838.950 307.950 841.050 310.050 ;
        RECT 849.600 306.300 851.700 308.400 ;
        RECT 852.600 306.300 855.600 308.400 ;
        RECT 827.700 281.700 828.900 303.300 ;
        RECT 830.700 301.500 832.200 306.300 ;
        RECT 833.100 303.300 835.200 305.400 ;
        RECT 830.100 299.400 832.200 301.500 ;
        RECT 830.700 281.700 832.200 299.400 ;
        RECT 833.700 296.100 834.900 303.300 ;
        RECT 838.500 301.800 840.600 303.900 ;
        RECT 847.200 303.300 849.300 305.400 ;
        RECT 833.100 294.000 835.200 296.100 ;
        RECT 839.700 295.200 840.600 301.800 ;
        RECT 833.700 281.700 834.900 294.000 ;
        RECT 838.500 293.100 840.600 295.200 ;
        RECT 835.800 286.500 837.900 288.600 ;
        RECT 839.700 282.600 840.600 293.100 ;
        RECT 841.950 291.000 844.050 295.050 ;
        RECT 842.400 289.350 843.600 291.000 ;
        RECT 842.100 286.950 844.200 289.050 ;
        RECT 827.700 279.600 829.800 281.700 ;
        RECT 830.700 279.600 832.800 281.700 ;
        RECT 833.700 279.600 835.800 281.700 ;
        RECT 839.100 280.500 841.200 282.600 ;
        RECT 848.100 281.700 849.300 303.300 ;
        RECT 850.500 300.300 851.700 306.300 ;
        RECT 850.500 298.200 852.600 300.300 ;
        RECT 850.500 281.700 851.700 298.200 ;
        RECT 854.100 287.400 855.600 306.300 ;
        RECT 865.950 296.100 868.050 298.200 ;
        RECT 866.400 295.350 867.600 296.100 ;
        RECT 856.950 292.950 859.050 295.050 ;
        RECT 860.100 292.950 862.200 295.050 ;
        RECT 866.100 292.950 868.200 295.050 ;
        RECT 853.500 285.300 855.600 287.400 ;
        RECT 853.500 281.700 854.700 285.300 ;
        RECT 847.200 279.600 849.300 281.700 ;
        RECT 850.200 279.600 852.300 281.700 ;
        RECT 853.200 279.600 855.300 281.700 ;
        RECT 857.400 280.050 858.450 292.950 ;
        RECT 868.950 283.950 871.050 286.050 ;
        RECT 856.950 277.950 859.050 280.050 ;
        RECT 820.950 268.950 823.050 271.050 ;
        RECT 811.950 265.950 814.050 268.050 ;
        RECT 817.950 265.950 820.050 268.050 ;
        RECT 836.700 267.300 838.800 269.400 ;
        RECT 839.700 267.300 841.800 269.400 ;
        RECT 842.700 267.300 844.800 269.400 ;
        RECT 818.400 262.200 819.450 265.950 ;
        RECT 837.300 263.700 838.500 267.300 ;
        RECT 811.950 260.100 814.050 262.200 ;
        RECT 817.950 260.100 820.050 262.200 ;
        RECT 836.400 261.600 838.500 263.700 ;
        RECT 812.400 259.350 813.600 260.100 ;
        RECT 818.400 259.350 819.600 260.100 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 808.950 253.950 811.050 256.050 ;
        RECT 815.400 254.400 816.600 256.650 ;
        RECT 805.950 247.950 808.050 250.050 ;
        RECT 809.400 244.050 810.450 253.950 ;
        RECT 808.950 241.950 811.050 244.050 ;
        RECT 815.400 241.050 816.450 254.400 ;
        RECT 823.800 253.950 825.900 256.050 ;
        RECT 829.800 253.950 831.900 256.050 ;
        RECT 824.400 252.000 825.600 253.650 ;
        RECT 823.950 247.950 826.050 252.000 ;
        RECT 826.950 250.950 829.050 253.050 ;
        RECT 814.950 238.950 817.050 241.050 ;
        RECT 808.950 235.950 811.050 238.050 ;
        RECT 785.400 230.400 789.450 231.450 ;
        RECT 782.100 214.950 784.200 217.050 ;
        RECT 782.400 213.450 783.600 214.650 ;
        RECT 788.400 213.900 789.450 230.400 ;
        RECT 791.700 228.300 793.800 230.400 ;
        RECT 792.300 223.500 793.800 228.300 ;
        RECT 791.700 221.400 793.800 223.500 ;
        RECT 779.400 212.400 783.600 213.450 ;
        RECT 787.950 211.800 790.050 213.900 ;
        RECT 739.950 208.800 742.050 210.900 ;
        RECT 745.950 208.800 748.050 210.900 ;
        RECT 730.950 205.950 733.050 208.050 ;
        RECT 746.400 205.050 747.450 208.800 ;
        RECT 752.400 208.050 753.450 211.800 ;
        RECT 758.400 209.400 759.600 211.650 ;
        RECT 764.400 210.000 765.600 211.650 ;
        RECT 751.950 205.950 754.050 208.050 ;
        RECT 745.950 202.950 748.050 205.050 ;
        RECT 758.400 199.050 759.450 209.400 ;
        RECT 763.950 205.950 766.050 210.000 ;
        RECT 784.950 208.950 787.050 211.050 ;
        RECT 760.950 202.950 763.050 205.050 ;
        RECT 751.950 196.950 754.050 199.050 ;
        RECT 757.950 196.950 760.050 199.050 ;
        RECT 739.950 193.950 742.050 196.050 ;
        RECT 740.400 189.450 741.450 193.950 ;
        RECT 740.400 187.200 741.600 189.450 ;
        RECT 735.900 183.900 738.000 185.700 ;
        RECT 739.800 184.800 741.900 186.900 ;
        RECT 743.100 186.300 745.200 188.400 ;
        RECT 734.400 182.700 743.100 183.900 ;
        RECT 731.100 178.950 733.200 181.050 ;
        RECT 731.400 177.450 732.600 178.650 ;
        RECT 728.400 176.400 732.600 177.450 ;
        RECT 728.400 148.050 729.450 176.400 ;
        RECT 734.400 173.700 735.300 182.700 ;
        RECT 741.000 181.800 743.100 182.700 ;
        RECT 744.000 180.900 744.900 186.300 ;
        RECT 745.950 182.100 748.050 184.200 ;
        RECT 746.400 181.350 747.600 182.100 ;
        RECT 738.000 179.700 744.900 180.900 ;
        RECT 738.000 177.300 738.900 179.700 ;
        RECT 736.800 175.200 738.900 177.300 ;
        RECT 739.800 175.950 741.900 178.050 ;
        RECT 733.500 171.600 735.600 173.700 ;
        RECT 740.400 173.400 741.600 175.650 ;
        RECT 743.700 172.500 744.900 179.700 ;
        RECT 745.800 178.950 747.900 181.050 ;
        RECT 743.100 170.400 745.200 172.500 ;
        RECT 736.950 154.950 739.050 157.050 ;
        RECT 727.950 145.950 730.050 148.050 ;
        RECT 721.950 137.100 724.050 139.200 ;
        RECT 730.950 137.100 733.050 139.200 ;
        RECT 737.400 138.600 738.450 154.950 ;
        RECT 722.400 127.050 723.450 137.100 ;
        RECT 731.400 136.350 732.600 137.100 ;
        RECT 737.400 136.350 738.600 138.600 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 728.400 132.900 729.600 133.650 ;
        RECT 727.950 130.800 730.050 132.900 ;
        RECT 734.400 131.400 735.600 133.650 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 727.950 121.950 730.050 124.050 ;
        RECT 721.950 118.950 724.050 121.050 ;
        RECT 722.400 102.600 723.450 118.950 ;
        RECT 722.400 100.350 723.600 102.600 ;
        RECT 722.100 97.950 724.200 100.050 ;
        RECT 718.950 61.950 721.050 64.050 ;
        RECT 712.950 59.100 715.050 61.200 ;
        RECT 719.400 60.600 720.450 61.950 ;
        RECT 728.400 61.200 729.450 121.950 ;
        RECT 734.400 118.050 735.450 131.400 ;
        RECT 752.400 124.050 753.450 196.950 ;
        RECT 761.400 183.450 762.450 202.950 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 770.400 183.600 771.450 187.950 ;
        RECT 764.400 183.450 765.600 183.600 ;
        RECT 761.400 182.400 765.600 183.450 ;
        RECT 764.400 181.350 765.600 182.400 ;
        RECT 770.400 181.350 771.600 183.600 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 769.950 178.950 772.050 181.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 767.400 176.400 768.600 178.650 ;
        RECT 773.400 177.900 774.600 178.650 ;
        RECT 767.400 166.050 768.450 176.400 ;
        RECT 772.950 175.800 775.050 177.900 ;
        RECT 766.950 163.950 769.050 166.050 ;
        RECT 778.950 157.950 781.050 160.050 ;
        RECT 776.400 138.450 777.600 138.600 ;
        RECT 779.400 138.450 780.450 157.950 ;
        RECT 776.400 137.400 780.450 138.450 ;
        RECT 776.400 136.350 777.600 137.400 ;
        RECT 757.800 133.950 759.900 136.050 ;
        RECT 775.800 133.950 777.900 136.050 ;
        RECT 751.950 121.950 754.050 124.050 ;
        RECT 779.400 121.050 780.450 137.400 ;
        RECT 785.400 124.050 786.450 208.950 ;
        RECT 792.300 203.700 793.800 221.400 ;
        RECT 791.700 201.600 793.800 203.700 ;
        RECT 794.700 225.300 796.800 230.400 ;
        RECT 797.700 228.300 799.800 230.400 ;
        RECT 802.950 229.950 805.050 232.050 ;
        RECT 794.700 203.700 795.900 225.300 ;
        RECT 797.700 223.500 799.200 228.300 ;
        RECT 800.100 225.300 802.200 227.400 ;
        RECT 797.100 221.400 799.200 223.500 ;
        RECT 797.700 203.700 799.200 221.400 ;
        RECT 800.700 218.100 801.900 225.300 ;
        RECT 805.500 223.800 807.600 225.900 ;
        RECT 800.100 216.000 802.200 218.100 ;
        RECT 806.700 217.200 807.600 223.800 ;
        RECT 800.700 203.700 801.900 216.000 ;
        RECT 805.500 215.100 807.600 217.200 ;
        RECT 802.800 208.500 804.900 210.600 ;
        RECT 806.700 204.600 807.600 215.100 ;
        RECT 809.400 213.600 810.450 235.950 ;
        RECT 816.600 228.300 818.700 230.400 ;
        RECT 819.600 228.300 822.600 230.400 ;
        RECT 814.200 225.300 816.300 227.400 ;
        RECT 809.400 211.350 810.600 213.600 ;
        RECT 809.100 208.950 811.200 211.050 ;
        RECT 794.700 201.600 796.800 203.700 ;
        RECT 797.700 201.600 799.800 203.700 ;
        RECT 800.700 201.600 802.800 203.700 ;
        RECT 806.100 202.500 808.200 204.600 ;
        RECT 815.100 203.700 816.300 225.300 ;
        RECT 817.500 222.300 818.700 228.300 ;
        RECT 817.500 220.200 819.600 222.300 ;
        RECT 817.500 203.700 818.700 220.200 ;
        RECT 821.100 209.400 822.600 228.300 ;
        RECT 824.400 220.200 825.450 247.950 ;
        RECT 827.400 223.050 828.450 250.950 ;
        RECT 836.400 242.700 837.900 261.600 ;
        RECT 840.300 250.800 841.500 267.300 ;
        RECT 839.400 248.700 841.500 250.800 ;
        RECT 840.300 242.700 841.500 248.700 ;
        RECT 842.700 245.700 843.900 267.300 ;
        RECT 850.800 266.400 852.900 268.500 ;
        RECT 856.200 267.300 858.300 269.400 ;
        RECT 859.200 267.300 861.300 269.400 ;
        RECT 862.200 267.300 864.300 269.400 ;
        RECT 847.800 259.950 849.900 262.050 ;
        RECT 848.400 258.900 849.600 259.650 ;
        RECT 847.950 256.800 850.050 258.900 ;
        RECT 851.400 255.900 852.300 266.400 ;
        RECT 854.100 260.400 856.200 262.500 ;
        RECT 851.400 253.800 853.500 255.900 ;
        RECT 857.100 255.000 858.300 267.300 ;
        RECT 847.950 250.950 850.050 253.050 ;
        RECT 842.700 243.600 844.800 245.700 ;
        RECT 836.400 240.600 839.400 242.700 ;
        RECT 840.300 240.600 842.400 242.700 ;
        RECT 848.400 241.050 849.450 250.950 ;
        RECT 851.400 247.200 852.300 253.800 ;
        RECT 856.800 252.900 858.900 255.000 ;
        RECT 851.400 245.100 853.500 247.200 ;
        RECT 857.100 245.700 858.300 252.900 ;
        RECT 859.800 249.600 861.300 267.300 ;
        RECT 859.800 247.500 861.900 249.600 ;
        RECT 856.800 243.600 858.900 245.700 ;
        RECT 859.800 242.700 861.300 247.500 ;
        RECT 863.100 245.700 864.300 267.300 ;
        RECT 847.950 238.950 850.050 241.050 ;
        RECT 859.200 240.600 861.300 242.700 ;
        RECT 862.200 240.600 864.300 245.700 ;
        RECT 865.200 267.300 867.300 269.400 ;
        RECT 865.200 249.600 866.700 267.300 ;
        RECT 869.400 252.450 870.450 283.950 ;
        RECT 872.400 259.200 873.450 313.950 ;
        RECT 874.950 307.950 877.050 310.050 ;
        RECT 871.950 257.100 874.050 259.200 ;
        RECT 875.400 258.600 876.450 307.950 ;
        RECT 878.400 286.050 879.450 331.950 ;
        RECT 881.400 316.050 882.450 346.950 ;
        RECT 880.950 313.950 883.050 316.050 ;
        RECT 884.400 310.050 885.450 359.400 ;
        RECT 886.950 358.950 889.050 359.400 ;
        RECT 890.400 343.050 891.450 364.950 ;
        RECT 889.950 340.950 892.050 343.050 ;
        RECT 886.950 337.950 889.050 340.050 ;
        RECT 893.400 339.600 894.450 368.400 ;
        RECT 897.000 363.450 901.050 364.050 ;
        RECT 896.400 361.950 901.050 363.450 ;
        RECT 896.400 358.050 897.450 361.950 ;
        RECT 898.950 358.800 901.050 360.900 ;
        RECT 895.950 355.950 898.050 358.050 ;
        RECT 899.400 352.050 900.450 358.800 ;
        RECT 898.950 349.950 901.050 352.050 ;
        RECT 902.400 342.450 903.450 370.950 ;
        RECT 905.400 346.050 906.450 424.950 ;
        RECT 913.800 420.300 915.900 422.400 ;
        RECT 916.950 421.950 919.050 424.050 ;
        RECT 917.400 421.200 918.600 421.950 ;
        RECT 926.400 421.050 927.450 425.400 ;
        RECT 928.950 421.950 931.050 424.050 ;
        RECT 910.950 416.100 913.050 418.200 ;
        RECT 911.400 415.350 912.600 416.100 ;
        RECT 907.950 412.950 910.050 415.050 ;
        RECT 911.100 412.950 913.200 415.050 ;
        RECT 914.100 414.900 915.000 420.300 ;
        RECT 917.100 418.800 919.200 420.900 ;
        RECT 921.000 417.900 923.100 419.700 ;
        RECT 925.950 418.950 928.050 421.050 ;
        RECT 915.900 416.700 924.600 417.900 ;
        RECT 915.900 415.800 918.000 416.700 ;
        RECT 914.100 413.700 921.000 414.900 ;
        RECT 908.400 402.450 909.450 412.950 ;
        RECT 914.100 406.500 915.300 413.700 ;
        RECT 917.100 409.950 919.200 412.050 ;
        RECT 920.100 411.300 921.000 413.700 ;
        RECT 917.400 407.400 918.600 409.650 ;
        RECT 920.100 409.200 922.200 411.300 ;
        RECT 923.700 407.700 924.600 416.700 ;
        RECT 929.400 415.050 930.450 421.950 ;
        RECT 925.800 412.950 927.900 415.050 ;
        RECT 928.950 412.950 931.050 415.050 ;
        RECT 926.400 411.450 927.600 412.650 ;
        RECT 926.400 410.400 930.450 411.450 ;
        RECT 913.800 404.400 915.900 406.500 ;
        RECT 923.400 405.600 925.500 407.700 ;
        RECT 929.400 406.050 930.450 410.400 ;
        RECT 928.950 403.950 931.050 406.050 ;
        RECT 908.400 401.400 912.450 402.450 ;
        RECT 907.950 388.950 910.050 391.050 ;
        RECT 908.400 360.450 909.450 388.950 ;
        RECT 911.400 388.050 912.450 401.400 ;
        RECT 919.950 400.950 922.050 403.050 ;
        RECT 913.950 394.950 916.050 397.050 ;
        RECT 910.950 385.950 913.050 388.050 ;
        RECT 910.950 379.950 913.050 382.050 ;
        RECT 911.400 364.050 912.450 379.950 ;
        RECT 914.400 373.050 915.450 394.950 ;
        RECT 920.400 379.050 921.450 400.950 ;
        RECT 922.950 388.950 925.050 391.050 ;
        RECT 919.950 376.950 922.050 379.050 ;
        RECT 923.400 373.200 924.450 388.950 ;
        RECT 932.400 385.050 933.450 511.950 ;
        RECT 934.950 496.950 937.050 499.050 ;
        RECT 935.400 493.050 936.450 496.950 ;
        RECT 938.400 496.050 939.450 533.400 ;
        RECT 937.950 493.950 940.050 496.050 ;
        RECT 934.950 490.950 937.050 493.050 ;
        RECT 934.950 484.950 937.050 487.050 ;
        RECT 935.400 475.050 936.450 484.950 ;
        RECT 934.950 472.950 937.050 475.050 ;
        RECT 934.950 457.950 937.050 460.050 ;
        RECT 931.950 382.950 934.050 385.050 ;
        RECT 931.950 376.950 934.050 379.050 ;
        RECT 913.950 370.950 916.050 373.050 ;
        RECT 916.950 371.100 919.050 373.200 ;
        RECT 922.950 371.100 925.050 373.200 ;
        RECT 917.400 370.350 918.600 371.100 ;
        RECT 925.950 370.950 928.050 373.050 ;
        RECT 928.950 370.950 931.050 373.050 ;
        RECT 916.950 367.950 919.050 370.050 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 920.400 366.900 921.600 367.650 ;
        RECT 919.950 364.800 922.050 366.900 ;
        RECT 910.950 361.950 913.050 364.050 ;
        RECT 908.400 359.400 912.450 360.450 ;
        RECT 904.950 343.950 907.050 346.050 ;
        RECT 902.400 342.000 906.450 342.450 ;
        RECT 902.400 341.400 907.050 342.000 ;
        RECT 887.400 328.050 888.450 337.950 ;
        RECT 893.400 337.350 894.600 339.600 ;
        RECT 898.950 338.100 901.050 340.200 ;
        RECT 899.400 337.350 900.600 338.100 ;
        RECT 904.950 337.950 907.050 341.400 ;
        RECT 907.950 340.950 910.050 343.050 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 896.400 332.400 897.600 334.650 ;
        RECT 902.400 332.400 903.600 334.650 ;
        RECT 892.950 328.950 895.050 331.050 ;
        RECT 886.950 325.950 889.050 328.050 ;
        RECT 883.950 307.950 886.050 310.050 ;
        RECT 889.950 301.950 892.050 304.050 ;
        RECT 890.400 298.050 891.450 301.950 ;
        RECT 893.400 298.050 894.450 328.950 ;
        RECT 896.400 319.050 897.450 332.400 ;
        RECT 898.950 328.950 901.050 331.050 ;
        RECT 895.950 316.950 898.050 319.050 ;
        RECT 880.950 295.950 883.050 298.050 ;
        RECT 877.950 283.950 880.050 286.050 ;
        RECT 881.400 282.450 882.450 295.950 ;
        RECT 889.950 294.000 892.050 298.050 ;
        RECT 892.950 295.950 895.050 298.050 ;
        RECT 895.950 294.000 898.050 298.050 ;
        RECT 899.400 295.050 900.450 328.950 ;
        RECT 902.400 328.050 903.450 332.400 ;
        RECT 901.950 325.950 904.050 328.050 ;
        RECT 908.400 301.050 909.450 340.950 ;
        RECT 911.400 322.050 912.450 359.400 ;
        RECT 920.400 358.050 921.450 364.800 ;
        RECT 919.950 355.950 922.050 358.050 ;
        RECT 926.400 346.050 927.450 370.950 ;
        RECT 916.950 343.950 919.050 346.050 ;
        RECT 925.950 343.950 928.050 346.050 ;
        RECT 917.400 340.050 918.450 343.950 ;
        RECT 929.400 343.050 930.450 370.950 ;
        RECT 928.950 340.950 931.050 343.050 ;
        RECT 913.950 337.950 916.050 340.050 ;
        RECT 916.950 337.950 919.050 340.050 ;
        RECT 919.950 338.100 922.050 340.200 ;
        RECT 925.950 338.100 928.050 340.200 ;
        RECT 932.400 339.450 933.450 376.950 ;
        RECT 935.400 373.050 936.450 457.950 ;
        RECT 938.400 373.200 939.450 493.950 ;
        RECT 941.400 487.050 942.450 553.950 ;
        RECT 943.950 550.950 946.050 553.050 ;
        RECT 944.400 532.050 945.450 550.950 ;
        RECT 947.400 550.050 948.450 610.950 ;
        RECT 946.950 547.950 949.050 550.050 ;
        RECT 950.400 532.200 951.450 625.950 ;
        RECT 953.400 601.050 954.450 640.800 ;
        RECT 956.400 640.050 957.450 676.800 ;
        RECT 955.950 637.950 958.050 640.050 ;
        RECT 955.950 628.950 958.050 631.050 ;
        RECT 956.400 607.050 957.450 628.950 ;
        RECT 959.400 613.050 960.450 730.950 ;
        RECT 962.400 709.050 963.450 754.950 ;
        RECT 961.950 706.950 964.050 709.050 ;
        RECT 965.400 697.050 966.450 760.950 ;
        RECT 968.400 760.050 969.450 763.950 ;
        RECT 967.950 757.950 970.050 760.050 ;
        RECT 967.950 754.800 970.050 756.900 ;
        RECT 968.400 748.050 969.450 754.800 ;
        RECT 967.950 745.950 970.050 748.050 ;
        RECT 971.400 733.200 972.450 778.950 ;
        RECT 973.950 766.950 976.050 769.050 ;
        RECT 974.400 763.200 975.450 766.950 ;
        RECT 973.950 761.100 976.050 763.200 ;
        RECT 976.950 762.000 979.050 766.050 ;
        RECT 977.400 760.350 978.600 762.000 ;
        RECT 982.950 761.100 985.050 763.200 ;
        RECT 983.400 760.350 984.600 761.100 ;
        RECT 976.950 757.950 979.050 760.050 ;
        RECT 979.950 757.950 982.050 760.050 ;
        RECT 982.950 757.950 985.050 760.050 ;
        RECT 973.950 754.950 976.050 757.050 ;
        RECT 980.400 755.400 981.600 757.650 ;
        RECT 970.950 731.100 973.050 733.200 ;
        RECT 974.400 733.050 975.450 754.950 ;
        RECT 976.950 736.950 979.050 739.050 ;
        RECT 973.950 730.950 976.050 733.050 ;
        RECT 977.400 730.050 978.450 736.950 ;
        RECT 980.400 736.050 981.450 755.400 ;
        RECT 985.950 754.950 988.050 757.050 ;
        RECT 986.400 751.050 987.450 754.950 ;
        RECT 985.950 748.950 988.050 751.050 ;
        RECT 982.950 742.950 985.050 745.050 ;
        RECT 979.950 733.950 982.050 736.050 ;
        RECT 983.400 733.050 984.450 742.950 ;
        RECT 985.950 739.950 988.050 742.050 ;
        RECT 979.950 730.800 982.050 732.900 ;
        RECT 982.950 730.950 985.050 733.050 ;
        RECT 970.950 727.950 973.050 730.050 ;
        RECT 976.950 727.950 979.050 730.050 ;
        RECT 971.400 727.350 972.600 727.950 ;
        RECT 970.950 724.950 973.050 727.050 ;
        RECT 973.950 724.950 976.050 727.050 ;
        RECT 974.400 723.900 975.600 724.650 ;
        RECT 973.950 721.800 976.050 723.900 ;
        RECT 976.950 706.950 979.050 709.050 ;
        RECT 964.950 694.950 967.050 697.050 ;
        RECT 967.950 683.100 970.050 685.200 ;
        RECT 968.400 682.350 969.600 683.100 ;
        RECT 964.950 679.950 967.050 682.050 ;
        RECT 967.950 679.950 970.050 682.050 ;
        RECT 970.950 679.950 973.050 682.050 ;
        RECT 961.950 676.950 964.050 679.050 ;
        RECT 965.400 678.900 966.600 679.650 ;
        RECT 962.400 652.050 963.450 676.950 ;
        RECT 964.950 676.800 967.050 678.900 ;
        RECT 971.400 677.400 972.600 679.650 ;
        RECT 971.400 676.050 972.450 677.400 ;
        RECT 977.400 676.050 978.450 706.950 ;
        RECT 970.950 673.950 973.050 676.050 ;
        RECT 976.950 673.950 979.050 676.050 ;
        RECT 964.950 670.950 967.050 673.050 ;
        RECT 965.400 655.050 966.450 670.950 ;
        RECT 971.400 670.050 972.450 673.950 ;
        RECT 976.950 670.800 979.050 672.900 ;
        RECT 970.950 667.950 973.050 670.050 ;
        RECT 973.950 664.950 976.050 667.050 ;
        RECT 964.950 652.950 967.050 655.050 ;
        RECT 961.950 651.600 966.000 652.050 ;
        RECT 961.950 649.950 966.600 651.600 ;
        RECT 970.950 650.100 973.050 652.200 ;
        RECT 974.400 652.050 975.450 664.950 ;
        RECT 977.400 661.050 978.450 670.800 ;
        RECT 976.950 658.950 979.050 661.050 ;
        RECT 965.400 649.350 966.600 649.950 ;
        RECT 971.400 649.350 972.600 650.100 ;
        RECT 973.950 649.950 976.050 652.050 ;
        RECT 964.950 646.950 967.050 649.050 ;
        RECT 967.950 646.950 970.050 649.050 ;
        RECT 970.950 646.950 973.050 649.050 ;
        RECT 968.400 644.400 969.600 646.650 ;
        RECT 968.400 643.050 969.450 644.400 ;
        RECT 973.950 643.950 976.050 646.050 ;
        RECT 961.950 640.950 964.050 643.050 ;
        RECT 964.950 640.950 967.050 643.050 ;
        RECT 968.400 641.400 973.050 643.050 ;
        RECT 969.000 640.950 973.050 641.400 ;
        RECT 962.400 631.050 963.450 640.950 ;
        RECT 965.400 634.050 966.450 640.950 ;
        RECT 974.400 640.050 975.450 643.950 ;
        RECT 967.950 637.950 970.050 640.050 ;
        RECT 973.950 637.950 976.050 640.050 ;
        RECT 964.950 631.950 967.050 634.050 ;
        RECT 961.950 628.950 964.050 631.050 ;
        RECT 958.950 610.950 961.050 613.050 ;
        RECT 964.950 610.950 967.050 613.050 ;
        RECT 955.950 604.950 958.050 607.050 ;
        RECT 961.950 606.000 964.050 610.050 ;
        RECT 965.400 607.050 966.450 610.950 ;
        RECT 962.400 604.350 963.600 606.000 ;
        RECT 964.950 604.950 967.050 607.050 ;
        RECT 958.950 601.950 961.050 604.050 ;
        RECT 961.950 601.950 964.050 604.050 ;
        RECT 952.950 598.950 955.050 601.050 ;
        RECT 955.950 598.950 958.050 601.050 ;
        RECT 959.400 600.900 960.600 601.650 ;
        RECT 956.400 586.050 957.450 598.950 ;
        RECT 958.950 598.800 961.050 600.900 ;
        RECT 964.950 598.950 967.050 601.050 ;
        RECT 958.950 589.950 961.050 592.050 ;
        RECT 955.950 583.950 958.050 586.050 ;
        RECT 952.950 579.450 955.050 583.050 ;
        RECT 952.950 579.000 957.450 579.450 ;
        RECT 953.400 578.400 957.450 579.000 ;
        RECT 952.950 574.950 955.050 577.050 ;
        RECT 953.400 562.050 954.450 574.950 ;
        RECT 956.400 574.050 957.450 578.400 ;
        RECT 955.950 571.950 958.050 574.050 ;
        RECT 959.400 573.600 960.450 589.950 ;
        RECT 965.400 580.050 966.450 598.950 ;
        RECT 964.950 577.950 967.050 580.050 ;
        RECT 968.400 577.050 969.450 637.950 ;
        RECT 973.950 631.950 976.050 634.050 ;
        RECT 974.400 622.050 975.450 631.950 ;
        RECT 973.950 619.950 976.050 622.050 ;
        RECT 970.950 616.950 973.050 619.050 ;
        RECT 971.400 595.050 972.450 616.950 ;
        RECT 973.950 613.950 976.050 616.050 ;
        RECT 974.400 610.050 975.450 613.950 ;
        RECT 977.400 610.050 978.450 658.950 ;
        RECT 980.400 652.050 981.450 730.800 ;
        RECT 982.950 727.800 985.050 729.900 ;
        RECT 983.400 673.050 984.450 727.800 ;
        RECT 986.400 685.050 987.450 739.950 ;
        RECT 989.400 730.050 990.450 781.950 ;
        RECT 992.400 754.050 993.450 784.950 ;
        RECT 994.950 772.950 997.050 775.050 ;
        RECT 991.950 751.950 994.050 754.050 ;
        RECT 995.400 733.050 996.450 772.950 ;
        RECT 998.400 763.050 999.450 799.950 ;
        RECT 1001.400 787.050 1002.450 907.950 ;
        RECT 1004.400 898.050 1005.450 911.400 ;
        RECT 1003.950 895.950 1006.050 898.050 ;
        RECT 1003.950 884.100 1006.050 886.200 ;
        RECT 1004.400 880.050 1005.450 884.100 ;
        RECT 1003.950 877.950 1006.050 880.050 ;
        RECT 1007.400 855.450 1008.450 922.950 ;
        RECT 1010.400 907.050 1011.450 955.800 ;
        RECT 1013.400 949.050 1014.450 962.100 ;
        RECT 1031.400 961.350 1032.600 963.000 ;
        RECT 1027.950 958.950 1030.050 961.050 ;
        RECT 1030.950 958.950 1033.050 961.050 ;
        RECT 1033.950 958.950 1036.050 961.050 ;
        RECT 1028.400 956.400 1029.600 958.650 ;
        RECT 1034.400 956.400 1035.600 958.650 ;
        RECT 1012.950 946.950 1015.050 949.050 ;
        RECT 1013.400 912.900 1014.450 946.950 ;
        RECT 1028.400 925.050 1029.450 956.400 ;
        RECT 1027.950 922.950 1030.050 925.050 ;
        RECT 1021.950 917.100 1024.050 919.200 ;
        RECT 1022.400 916.350 1023.600 917.100 ;
        RECT 1018.950 913.950 1021.050 916.050 ;
        RECT 1021.950 913.950 1024.050 916.050 ;
        RECT 1024.950 913.950 1027.050 916.050 ;
        RECT 1019.400 912.900 1020.600 913.650 ;
        RECT 1012.950 910.800 1015.050 912.900 ;
        RECT 1018.950 910.800 1021.050 912.900 ;
        RECT 1025.400 911.400 1026.600 913.650 ;
        RECT 1025.400 907.050 1026.450 911.400 ;
        RECT 1009.950 904.950 1012.050 907.050 ;
        RECT 1018.950 904.950 1021.050 907.050 ;
        RECT 1024.950 904.950 1027.050 907.050 ;
        RECT 1019.400 885.600 1020.450 904.950 ;
        RECT 1019.400 883.350 1020.600 885.600 ;
        RECT 1015.950 880.950 1018.050 883.050 ;
        RECT 1018.950 880.950 1021.050 883.050 ;
        RECT 1021.950 880.950 1024.050 883.050 ;
        RECT 1016.400 879.900 1017.600 880.650 ;
        RECT 1015.950 877.800 1018.050 879.900 ;
        RECT 1022.400 879.000 1023.600 880.650 ;
        RECT 1004.400 854.400 1008.450 855.450 ;
        RECT 1004.400 841.050 1005.450 854.400 ;
        RECT 1006.950 850.950 1009.050 853.050 ;
        RECT 1003.950 838.950 1006.050 841.050 ;
        RECT 1007.400 840.600 1008.450 850.950 ;
        RECT 1007.400 838.350 1008.600 840.600 ;
        RECT 1012.950 840.000 1015.050 844.050 ;
        RECT 1016.400 841.050 1017.450 877.800 ;
        RECT 1021.950 874.950 1024.050 879.000 ;
        RECT 1021.950 859.950 1024.050 862.050 ;
        RECT 1018.950 844.950 1021.050 847.050 ;
        RECT 1013.400 838.350 1014.600 840.000 ;
        RECT 1015.950 838.950 1018.050 841.050 ;
        RECT 1006.950 835.950 1009.050 838.050 ;
        RECT 1009.950 835.950 1012.050 838.050 ;
        RECT 1012.950 835.950 1015.050 838.050 ;
        RECT 1003.950 832.950 1006.050 835.050 ;
        RECT 1010.400 834.900 1011.600 835.650 ;
        RECT 1004.400 811.050 1005.450 832.950 ;
        RECT 1009.950 832.800 1012.050 834.900 ;
        RECT 1006.950 826.950 1009.050 829.050 ;
        RECT 1003.950 808.950 1006.050 811.050 ;
        RECT 1003.950 805.800 1006.050 807.900 ;
        RECT 1000.950 784.950 1003.050 787.050 ;
        RECT 1004.400 784.050 1005.450 805.800 ;
        RECT 1003.950 781.950 1006.050 784.050 ;
        RECT 1007.400 766.050 1008.450 826.950 ;
        RECT 1019.400 814.050 1020.450 844.950 ;
        RECT 1022.400 826.050 1023.450 859.950 ;
        RECT 1034.400 847.050 1035.450 956.400 ;
        RECT 1033.950 844.950 1036.050 847.050 ;
        RECT 1024.950 839.100 1027.050 841.200 ;
        RECT 1030.950 839.100 1033.050 841.200 ;
        RECT 1036.950 839.100 1039.050 841.200 ;
        RECT 1021.950 823.950 1024.050 826.050 ;
        RECT 1009.950 811.950 1012.050 814.050 ;
        RECT 1018.950 811.950 1021.050 814.050 ;
        RECT 1010.400 808.050 1011.450 811.950 ;
        RECT 1009.950 805.950 1012.050 808.050 ;
        RECT 1015.950 806.100 1018.050 808.200 ;
        RECT 1021.950 806.100 1024.050 808.200 ;
        RECT 1025.400 808.050 1026.450 839.100 ;
        RECT 1031.400 838.350 1032.600 839.100 ;
        RECT 1037.400 838.350 1038.600 839.100 ;
        RECT 1030.950 835.950 1033.050 838.050 ;
        RECT 1033.950 835.950 1036.050 838.050 ;
        RECT 1036.950 835.950 1039.050 838.050 ;
        RECT 1039.950 835.950 1042.050 838.050 ;
        RECT 1034.400 833.400 1035.600 835.650 ;
        RECT 1040.400 833.400 1041.600 835.650 ;
        RECT 1034.400 828.450 1035.450 833.400 ;
        RECT 1040.400 829.050 1041.450 833.400 ;
        RECT 1042.950 832.950 1045.050 835.050 ;
        RECT 1031.400 827.400 1035.450 828.450 ;
        RECT 1016.400 805.350 1017.600 806.100 ;
        RECT 1022.400 805.350 1023.600 806.100 ;
        RECT 1024.950 805.950 1027.050 808.050 ;
        RECT 1027.950 806.100 1030.050 808.200 ;
        RECT 1012.950 802.950 1015.050 805.050 ;
        RECT 1015.950 802.950 1018.050 805.050 ;
        RECT 1018.950 802.950 1021.050 805.050 ;
        RECT 1021.950 802.950 1024.050 805.050 ;
        RECT 1013.400 802.050 1014.600 802.650 ;
        RECT 1009.950 800.400 1014.600 802.050 ;
        RECT 1019.400 800.400 1020.600 802.650 ;
        RECT 1028.400 801.450 1029.450 806.100 ;
        RECT 1025.400 800.400 1029.450 801.450 ;
        RECT 1009.950 799.950 1014.000 800.400 ;
        RECT 1010.400 793.050 1011.450 799.950 ;
        RECT 1012.950 798.450 1017.000 799.050 ;
        RECT 1012.950 796.950 1017.450 798.450 ;
        RECT 1009.950 790.950 1012.050 793.050 ;
        RECT 1006.950 763.950 1009.050 766.050 ;
        RECT 997.950 760.950 1000.050 763.050 ;
        RECT 1003.950 761.100 1006.050 763.200 ;
        RECT 1009.950 761.100 1012.050 763.200 ;
        RECT 1004.400 760.350 1005.600 761.100 ;
        RECT 1010.400 760.350 1011.600 761.100 ;
        RECT 1000.950 757.950 1003.050 760.050 ;
        RECT 1003.950 757.950 1006.050 760.050 ;
        RECT 1006.950 757.950 1009.050 760.050 ;
        RECT 1009.950 757.950 1012.050 760.050 ;
        RECT 1001.400 756.450 1002.600 757.650 ;
        RECT 998.400 755.400 1002.600 756.450 ;
        RECT 1007.400 756.000 1008.600 757.650 ;
        RECT 988.950 727.950 991.050 730.050 ;
        RECT 991.950 729.000 994.050 733.050 ;
        RECT 994.950 730.950 997.050 733.050 ;
        RECT 998.400 730.200 999.450 755.400 ;
        RECT 1006.950 754.050 1009.050 756.000 ;
        RECT 1012.950 754.950 1015.050 757.050 ;
        RECT 1006.800 753.000 1009.050 754.050 ;
        RECT 1006.800 751.950 1008.900 753.000 ;
        RECT 1009.950 751.950 1012.050 754.050 ;
        RECT 1006.950 745.950 1009.050 748.050 ;
        RECT 992.400 727.350 993.600 729.000 ;
        RECT 997.950 728.100 1000.050 730.200 ;
        RECT 998.400 727.350 999.600 728.100 ;
        RECT 1003.950 727.950 1006.050 730.050 ;
        RECT 991.950 724.950 994.050 727.050 ;
        RECT 994.950 724.950 997.050 727.050 ;
        RECT 997.950 724.950 1000.050 727.050 ;
        RECT 988.950 721.950 991.050 724.050 ;
        RECT 995.400 723.000 996.600 724.650 ;
        RECT 989.400 691.050 990.450 721.950 ;
        RECT 994.950 718.950 997.050 723.000 ;
        RECT 988.950 688.950 991.050 691.050 ;
        RECT 1000.950 688.950 1003.050 691.050 ;
        RECT 985.950 682.950 988.050 685.050 ;
        RECT 991.950 683.100 994.050 685.200 ;
        RECT 992.400 682.350 993.600 683.100 ;
        RECT 988.950 679.950 991.050 682.050 ;
        RECT 991.950 679.950 994.050 682.050 ;
        RECT 994.950 679.950 997.050 682.050 ;
        RECT 985.950 676.950 988.050 679.050 ;
        RECT 989.400 677.400 990.600 679.650 ;
        RECT 995.400 677.400 996.600 679.650 ;
        RECT 982.950 670.950 985.050 673.050 ;
        RECT 982.950 661.950 985.050 664.050 ;
        RECT 979.950 649.950 982.050 652.050 ;
        RECT 979.950 646.800 982.050 648.900 ;
        RECT 980.400 616.050 981.450 646.800 ;
        RECT 979.950 613.950 982.050 616.050 ;
        RECT 983.400 613.050 984.450 661.950 ;
        RECT 986.400 651.450 987.450 676.950 ;
        RECT 989.400 673.050 990.450 677.400 ;
        RECT 988.950 670.950 991.050 673.050 ;
        RECT 995.400 667.050 996.450 677.400 ;
        RECT 994.950 664.950 997.050 667.050 ;
        RECT 994.950 658.950 997.050 661.050 ;
        RECT 995.400 652.200 996.450 658.950 ;
        RECT 989.400 651.450 990.600 651.600 ;
        RECT 986.400 650.400 990.600 651.450 ;
        RECT 989.400 649.350 990.600 650.400 ;
        RECT 994.950 650.100 997.050 652.200 ;
        RECT 995.400 649.350 996.600 650.100 ;
        RECT 988.950 646.950 991.050 649.050 ;
        RECT 991.950 646.950 994.050 649.050 ;
        RECT 994.950 646.950 997.050 649.050 ;
        RECT 985.950 643.950 988.050 646.050 ;
        RECT 992.400 644.400 993.600 646.650 ;
        RECT 982.950 610.950 985.050 613.050 ;
        RECT 986.400 610.050 987.450 643.950 ;
        RECT 988.950 640.950 991.050 643.050 ;
        RECT 992.400 637.050 993.450 644.400 ;
        RECT 997.950 643.950 1000.050 646.050 ;
        RECT 991.950 634.950 994.050 637.050 ;
        RECT 973.950 607.950 976.050 610.050 ;
        RECT 976.950 607.950 979.050 610.050 ;
        RECT 985.950 607.950 988.050 610.050 ;
        RECT 994.950 607.950 997.050 610.050 ;
        RECT 977.400 606.450 978.450 607.950 ;
        RECT 974.400 605.400 978.450 606.450 ;
        RECT 970.950 592.950 973.050 595.050 ;
        RECT 959.400 571.350 960.600 573.600 ;
        RECT 964.950 573.000 967.050 576.900 ;
        RECT 968.400 575.400 973.050 577.050 ;
        RECT 969.000 574.950 973.050 575.400 ;
        RECT 965.400 571.350 966.600 573.000 ;
        RECT 958.950 568.950 961.050 571.050 ;
        RECT 961.950 568.950 964.050 571.050 ;
        RECT 964.950 568.950 967.050 571.050 ;
        RECT 967.950 568.950 970.050 571.050 ;
        RECT 955.950 565.950 958.050 568.050 ;
        RECT 962.400 567.900 963.600 568.650 ;
        RECT 968.400 567.900 969.600 568.650 ;
        RECT 952.950 559.950 955.050 562.050 ;
        RECT 956.400 550.050 957.450 565.950 ;
        RECT 961.950 565.800 964.050 567.900 ;
        RECT 967.950 565.800 970.050 567.900 ;
        RECT 970.950 565.950 973.050 568.050 ;
        RECT 974.400 567.900 975.450 605.400 ;
        RECT 982.950 605.100 985.050 607.200 ;
        RECT 983.400 604.350 984.600 605.100 ;
        RECT 988.950 604.950 991.050 607.050 ;
        RECT 979.950 601.950 982.050 604.050 ;
        RECT 982.950 601.950 985.050 604.050 ;
        RECT 985.950 601.950 988.050 604.050 ;
        RECT 980.400 600.900 981.600 601.650 ;
        RECT 979.950 600.450 982.050 600.900 ;
        RECT 977.400 599.400 982.050 600.450 ;
        RECT 977.400 592.050 978.450 599.400 ;
        RECT 979.950 598.800 982.050 599.400 ;
        RECT 986.400 599.400 987.600 601.650 ;
        RECT 986.400 595.050 987.450 599.400 ;
        RECT 985.950 592.950 988.050 595.050 ;
        RECT 976.950 589.950 979.050 592.050 ;
        RECT 982.950 589.950 985.050 592.050 ;
        RECT 976.950 583.950 979.050 586.050 ;
        RECT 967.950 562.650 970.050 564.750 ;
        RECT 961.950 556.950 964.050 562.050 ;
        RECT 964.950 559.950 967.050 562.050 ;
        RECT 955.950 547.950 958.050 550.050 ;
        RECT 961.950 547.950 964.050 550.050 ;
        RECT 955.950 535.950 958.050 538.050 ;
        RECT 943.950 529.950 946.050 532.050 ;
        RECT 949.950 530.100 952.050 532.200 ;
        RECT 943.950 526.800 946.050 528.900 ;
        RECT 949.950 526.950 952.050 529.050 ;
        RECT 956.400 528.600 957.450 535.950 ;
        RECT 962.400 529.050 963.450 547.950 ;
        RECT 944.400 514.050 945.450 526.800 ;
        RECT 950.400 526.350 951.600 526.950 ;
        RECT 956.400 526.350 957.600 528.600 ;
        RECT 961.950 526.950 964.050 529.050 ;
        RECT 949.950 523.950 952.050 526.050 ;
        RECT 952.950 523.950 955.050 526.050 ;
        RECT 955.950 523.950 958.050 526.050 ;
        RECT 958.950 523.950 961.050 526.050 ;
        RECT 946.950 520.950 949.050 523.050 ;
        RECT 953.400 522.900 954.600 523.650 ;
        RECT 959.400 522.900 960.600 523.650 ;
        RECT 952.950 520.800 955.050 522.900 ;
        RECT 958.950 522.450 961.050 522.900 ;
        RECT 958.950 521.400 963.450 522.450 ;
        RECT 958.950 520.800 961.050 521.400 ;
        RECT 955.950 517.950 958.050 520.050 ;
        RECT 943.950 511.950 946.050 514.050 ;
        RECT 943.950 505.950 946.050 508.050 ;
        RECT 940.950 484.950 943.050 487.050 ;
        RECT 940.950 478.950 943.050 481.050 ;
        RECT 941.400 418.050 942.450 478.950 ;
        RECT 944.400 442.050 945.450 505.950 ;
        RECT 952.950 494.100 955.050 496.200 ;
        RECT 956.400 496.050 957.450 517.950 ;
        RECT 958.950 508.950 961.050 511.050 ;
        RECT 953.400 493.350 954.600 494.100 ;
        RECT 955.950 493.950 958.050 496.050 ;
        RECT 949.950 490.950 952.050 493.050 ;
        RECT 952.950 490.950 955.050 493.050 ;
        RECT 946.950 487.950 949.050 490.050 ;
        RECT 950.400 488.400 951.600 490.650 ;
        RECT 947.400 478.050 948.450 487.950 ;
        RECT 946.950 475.950 949.050 478.050 ;
        RECT 947.400 466.050 948.450 475.950 ;
        RECT 950.400 469.050 951.450 488.400 ;
        RECT 949.950 466.950 952.050 469.050 ;
        RECT 946.950 463.950 949.050 466.050 ;
        RECT 959.400 463.050 960.450 508.950 ;
        RECT 962.400 502.050 963.450 521.400 ;
        RECT 965.400 517.050 966.450 559.950 ;
        RECT 968.400 535.050 969.450 562.650 ;
        RECT 971.400 556.050 972.450 565.950 ;
        RECT 973.950 565.800 976.050 567.900 ;
        RECT 977.400 562.050 978.450 583.950 ;
        RECT 979.950 577.950 982.050 580.050 ;
        RECT 980.400 565.050 981.450 577.950 ;
        RECT 983.400 574.050 984.450 589.950 ;
        RECT 986.400 580.050 987.450 592.950 ;
        RECT 995.400 583.050 996.450 607.950 ;
        RECT 998.400 607.050 999.450 643.950 ;
        RECT 1001.400 610.050 1002.450 688.950 ;
        RECT 1004.400 679.050 1005.450 727.950 ;
        RECT 1003.950 676.950 1006.050 679.050 ;
        RECT 1003.950 667.950 1006.050 670.050 ;
        RECT 1004.400 642.450 1005.450 667.950 ;
        RECT 1007.400 646.050 1008.450 745.950 ;
        RECT 1010.400 685.050 1011.450 751.950 ;
        RECT 1013.400 748.050 1014.450 754.950 ;
        RECT 1016.400 751.050 1017.450 796.950 ;
        RECT 1019.400 766.050 1020.450 800.400 ;
        RECT 1021.950 796.950 1024.050 799.050 ;
        RECT 1018.950 763.950 1021.050 766.050 ;
        RECT 1018.950 760.800 1021.050 762.900 ;
        RECT 1015.950 748.950 1018.050 751.050 ;
        RECT 1012.950 745.950 1015.050 748.050 ;
        RECT 1019.400 729.600 1020.450 760.800 ;
        RECT 1022.400 754.050 1023.450 796.950 ;
        RECT 1021.950 751.950 1024.050 754.050 ;
        RECT 1021.950 748.800 1024.050 750.900 ;
        RECT 1022.400 738.450 1023.450 748.800 ;
        RECT 1025.400 742.050 1026.450 800.400 ;
        RECT 1027.950 766.950 1030.050 769.050 ;
        RECT 1028.400 762.600 1029.450 766.950 ;
        RECT 1031.400 766.050 1032.450 827.400 ;
        RECT 1039.950 826.950 1042.050 829.050 ;
        RECT 1033.950 823.950 1036.050 826.050 ;
        RECT 1034.400 808.050 1035.450 823.950 ;
        RECT 1039.950 820.950 1042.050 823.050 ;
        RECT 1033.950 805.950 1036.050 808.050 ;
        RECT 1040.400 807.600 1041.450 820.950 ;
        RECT 1043.400 808.050 1044.450 832.950 ;
        RECT 1040.400 805.350 1041.600 807.600 ;
        RECT 1042.950 805.950 1045.050 808.050 ;
        RECT 1036.950 802.950 1039.050 805.050 ;
        RECT 1039.950 802.950 1042.050 805.050 ;
        RECT 1037.400 802.050 1038.600 802.650 ;
        RECT 1033.950 800.400 1038.600 802.050 ;
        RECT 1033.950 799.950 1038.000 800.400 ;
        RECT 1042.950 799.950 1045.050 802.050 ;
        RECT 1034.400 775.050 1035.450 799.950 ;
        RECT 1039.950 781.950 1042.050 784.050 ;
        RECT 1033.950 772.950 1036.050 775.050 ;
        RECT 1036.950 769.950 1039.050 772.050 ;
        RECT 1030.950 763.950 1033.050 766.050 ;
        RECT 1037.400 762.600 1038.450 769.950 ;
        RECT 1028.400 760.350 1029.600 762.600 ;
        RECT 1037.400 760.350 1038.600 762.600 ;
        RECT 1028.100 757.950 1030.200 760.050 ;
        RECT 1033.500 757.950 1035.600 760.050 ;
        RECT 1036.800 757.950 1038.900 760.050 ;
        RECT 1034.400 755.400 1035.600 757.650 ;
        RECT 1027.950 751.950 1030.050 754.050 ;
        RECT 1024.950 739.950 1027.050 742.050 ;
        RECT 1022.400 737.400 1026.450 738.450 ;
        RECT 1025.400 730.050 1026.450 737.400 ;
        RECT 1019.400 727.350 1020.600 729.600 ;
        RECT 1024.950 727.950 1027.050 730.050 ;
        RECT 1015.950 724.950 1018.050 727.050 ;
        RECT 1018.950 724.950 1021.050 727.050 ;
        RECT 1021.950 724.950 1024.050 727.050 ;
        RECT 1016.400 723.000 1017.600 724.650 ;
        RECT 1022.400 723.000 1023.600 724.650 ;
        RECT 1015.950 718.950 1018.050 723.000 ;
        RECT 1021.950 718.950 1024.050 723.000 ;
        RECT 1024.950 694.950 1027.050 697.050 ;
        RECT 1009.950 682.950 1012.050 685.050 ;
        RECT 1015.950 683.100 1018.050 685.200 ;
        RECT 1021.950 683.100 1024.050 685.200 ;
        RECT 1025.400 685.050 1026.450 694.950 ;
        RECT 1016.400 682.350 1017.600 683.100 ;
        RECT 1022.400 682.350 1023.600 683.100 ;
        RECT 1024.950 682.950 1027.050 685.050 ;
        RECT 1012.950 679.950 1015.050 682.050 ;
        RECT 1015.950 679.950 1018.050 682.050 ;
        RECT 1018.950 679.950 1021.050 682.050 ;
        RECT 1021.950 679.950 1024.050 682.050 ;
        RECT 1013.400 678.900 1014.600 679.650 ;
        RECT 1012.950 676.800 1015.050 678.900 ;
        RECT 1019.400 677.400 1020.600 679.650 ;
        RECT 1015.950 673.950 1018.050 676.050 ;
        RECT 1016.400 651.600 1017.450 673.950 ;
        RECT 1019.400 670.050 1020.450 677.400 ;
        RECT 1024.950 676.950 1027.050 679.050 ;
        RECT 1018.950 667.950 1021.050 670.050 ;
        RECT 1016.400 649.350 1017.600 651.600 ;
        RECT 1012.950 646.950 1015.050 649.050 ;
        RECT 1015.950 646.950 1018.050 649.050 ;
        RECT 1018.950 646.950 1021.050 649.050 ;
        RECT 1006.950 643.950 1009.050 646.050 ;
        RECT 1013.400 644.400 1014.600 646.650 ;
        RECT 1019.400 644.400 1020.600 646.650 ;
        RECT 1004.400 641.400 1008.450 642.450 ;
        RECT 1000.950 607.950 1003.050 610.050 ;
        RECT 997.950 604.950 1000.050 607.050 ;
        RECT 1007.400 606.600 1008.450 641.400 ;
        RECT 1013.400 637.050 1014.450 644.400 ;
        RECT 1012.950 634.950 1015.050 637.050 ;
        RECT 1012.950 628.950 1015.050 631.050 ;
        RECT 1013.400 613.050 1014.450 628.950 ;
        RECT 1019.400 622.050 1020.450 644.400 ;
        RECT 1018.950 621.450 1021.050 622.050 ;
        RECT 1025.400 621.450 1026.450 676.950 ;
        RECT 1016.400 620.400 1021.050 621.450 ;
        RECT 1012.950 610.950 1015.050 613.050 ;
        RECT 998.400 600.900 999.450 604.950 ;
        RECT 1007.400 604.350 1008.600 606.600 ;
        RECT 1003.950 601.950 1006.050 604.050 ;
        RECT 1006.950 601.950 1009.050 604.050 ;
        RECT 1009.950 601.950 1012.050 604.050 ;
        RECT 1004.400 600.900 1005.600 601.650 ;
        RECT 997.950 598.800 1000.050 600.900 ;
        RECT 1003.950 598.800 1006.050 600.900 ;
        RECT 1010.400 599.400 1011.600 601.650 ;
        RECT 1010.400 597.450 1011.450 599.400 ;
        RECT 1016.400 598.050 1017.450 620.400 ;
        RECT 1018.950 619.950 1021.050 620.400 ;
        RECT 1022.400 620.400 1026.450 621.450 ;
        RECT 1018.950 607.950 1021.050 610.050 ;
        RECT 1019.400 601.050 1020.450 607.950 ;
        RECT 1018.950 598.950 1021.050 601.050 ;
        RECT 1004.400 596.400 1011.450 597.450 ;
        RECT 997.950 589.950 1000.050 592.050 ;
        RECT 994.950 580.950 997.050 583.050 ;
        RECT 985.950 577.950 988.050 580.050 ;
        RECT 994.950 577.800 997.050 579.900 ;
        RECT 982.950 571.950 985.050 574.050 ;
        RECT 988.950 572.100 991.050 574.200 ;
        RECT 995.400 574.050 996.450 577.800 ;
        RECT 989.400 571.350 990.600 572.100 ;
        RECT 994.950 571.950 997.050 574.050 ;
        RECT 985.950 568.950 988.050 571.050 ;
        RECT 988.950 568.950 991.050 571.050 ;
        RECT 991.950 568.950 994.050 571.050 ;
        RECT 986.400 567.900 987.600 568.650 ;
        RECT 992.400 567.900 993.600 568.650 ;
        RECT 985.950 565.800 988.050 567.900 ;
        RECT 991.950 565.800 994.050 567.900 ;
        RECT 979.950 562.950 982.050 565.050 ;
        RECT 976.950 556.950 979.050 562.050 ;
        RECT 970.950 553.950 973.050 556.050 ;
        RECT 970.950 550.800 973.050 552.900 ;
        RECT 967.950 532.950 970.050 535.050 ;
        RECT 971.400 531.450 972.450 550.800 ;
        RECT 976.950 547.950 979.050 550.050 ;
        RECT 973.950 532.950 976.050 535.050 ;
        RECT 968.400 530.400 972.450 531.450 ;
        RECT 964.950 514.950 967.050 517.050 ;
        RECT 961.950 499.950 964.050 502.050 ;
        RECT 964.950 499.950 967.050 502.050 ;
        RECT 961.950 493.950 964.050 496.050 ;
        RECT 958.950 460.950 961.050 463.050 ;
        RECT 962.400 460.050 963.450 493.950 ;
        RECT 965.400 493.050 966.450 499.950 ;
        RECT 968.400 496.050 969.450 530.400 ;
        RECT 974.400 529.050 975.450 532.950 ;
        RECT 977.400 532.050 978.450 547.950 ;
        RECT 982.950 544.950 985.050 547.050 ;
        RECT 979.950 532.050 982.050 532.200 ;
        RECT 983.400 532.050 984.450 544.950 ;
        RECT 986.400 538.050 987.450 565.800 ;
        RECT 998.400 553.050 999.450 589.950 ;
        RECT 1000.950 580.950 1003.050 583.050 ;
        RECT 1001.400 553.050 1002.450 580.950 ;
        RECT 1004.400 568.050 1005.450 596.400 ;
        RECT 1015.950 595.950 1018.050 598.050 ;
        RECT 1009.950 592.950 1012.050 595.050 ;
        RECT 1010.400 583.050 1011.450 592.950 ;
        RECT 1012.950 583.950 1015.050 586.050 ;
        RECT 1009.950 580.950 1012.050 583.050 ;
        RECT 1013.400 576.450 1014.450 583.950 ;
        RECT 1010.400 575.400 1014.450 576.450 ;
        RECT 1010.400 573.600 1011.450 575.400 ;
        RECT 1010.400 571.350 1011.600 573.600 ;
        RECT 1015.950 572.100 1018.050 574.200 ;
        RECT 1016.400 571.350 1017.600 572.100 ;
        RECT 1009.950 568.950 1012.050 571.050 ;
        RECT 1012.950 568.950 1015.050 571.050 ;
        RECT 1015.950 568.950 1018.050 571.050 ;
        RECT 1003.950 565.950 1006.050 568.050 ;
        RECT 1006.950 565.950 1009.050 568.050 ;
        RECT 1013.400 567.900 1014.600 568.650 ;
        RECT 994.950 550.950 997.050 553.050 ;
        RECT 997.950 550.950 1000.050 553.050 ;
        RECT 1000.950 550.950 1003.050 553.050 ;
        RECT 985.950 535.950 988.050 538.050 ;
        RECT 991.950 535.950 994.050 538.050 ;
        RECT 977.400 530.700 982.050 532.050 ;
        RECT 978.000 530.100 982.050 530.700 ;
        RECT 978.000 529.950 981.000 530.100 ;
        RECT 982.950 529.950 985.050 532.050 ;
        RECT 970.950 526.950 973.050 529.050 ;
        RECT 973.950 526.950 976.050 529.050 ;
        RECT 979.950 526.950 982.050 529.050 ;
        RECT 985.950 528.000 988.050 532.050 ;
        RECT 971.400 502.050 972.450 526.950 ;
        RECT 980.400 526.350 981.600 526.950 ;
        RECT 986.400 526.350 987.600 528.000 ;
        RECT 976.950 523.950 979.050 526.050 ;
        RECT 979.950 523.950 982.050 526.050 ;
        RECT 982.950 523.950 985.050 526.050 ;
        RECT 985.950 523.950 988.050 526.050 ;
        RECT 973.950 520.950 976.050 523.050 ;
        RECT 977.400 521.400 978.600 523.650 ;
        RECT 983.400 521.400 984.600 523.650 ;
        RECT 974.400 508.050 975.450 520.950 ;
        RECT 977.400 514.050 978.450 521.400 ;
        RECT 976.950 511.950 979.050 514.050 ;
        RECT 973.950 505.950 976.050 508.050 ;
        RECT 970.950 499.950 973.050 502.050 ;
        RECT 967.950 493.950 970.050 496.050 ;
        RECT 970.950 495.000 973.050 498.900 ;
        RECT 974.400 498.450 975.450 505.950 ;
        RECT 983.400 505.050 984.450 521.400 ;
        RECT 988.950 520.950 991.050 523.050 ;
        RECT 989.400 511.050 990.450 520.950 ;
        RECT 988.950 508.950 991.050 511.050 ;
        RECT 992.400 507.450 993.450 535.950 ;
        RECT 989.400 506.400 993.450 507.450 ;
        RECT 982.950 502.950 985.050 505.050 ;
        RECT 982.950 499.800 985.050 501.900 ;
        RECT 974.400 497.400 978.450 498.450 ;
        RECT 977.400 495.600 978.450 497.400 ;
        RECT 971.400 493.350 972.600 495.000 ;
        RECT 977.400 493.350 978.600 495.600 ;
        RECT 964.950 490.950 967.050 493.050 ;
        RECT 970.950 490.950 973.050 493.050 ;
        RECT 973.950 490.950 976.050 493.050 ;
        RECT 976.950 490.950 979.050 493.050 ;
        RECT 967.950 487.950 970.050 490.050 ;
        RECT 974.400 488.400 975.600 490.650 ;
        RECT 964.950 469.950 967.050 472.050 ;
        RECT 961.950 457.950 964.050 460.050 ;
        RECT 965.400 457.050 966.450 469.950 ;
        RECT 968.400 465.450 969.450 487.950 ;
        RECT 974.400 481.050 975.450 488.400 ;
        RECT 983.400 484.050 984.450 499.800 ;
        RECT 985.950 496.950 988.050 499.050 ;
        RECT 976.950 481.950 979.050 484.050 ;
        RECT 982.950 481.950 985.050 484.050 ;
        RECT 973.950 478.950 976.050 481.050 ;
        RECT 970.800 472.950 972.900 475.050 ;
        RECT 973.950 472.950 976.050 475.050 ;
        RECT 971.400 469.050 972.450 472.950 ;
        RECT 970.950 466.950 973.050 469.050 ;
        RECT 968.400 464.400 972.450 465.450 ;
        RECT 967.950 460.950 970.050 463.050 ;
        RECT 949.800 454.500 951.900 456.600 ;
        RECT 947.100 445.950 949.200 448.050 ;
        RECT 950.100 447.300 951.300 454.500 ;
        RECT 953.400 451.350 954.600 453.600 ;
        RECT 959.400 453.300 961.500 455.400 ;
        RECT 964.950 454.950 967.050 457.050 ;
        RECT 953.100 448.950 955.200 451.050 ;
        RECT 956.100 449.700 958.200 451.800 ;
        RECT 956.100 447.300 957.000 449.700 ;
        RECT 950.100 446.100 957.000 447.300 ;
        RECT 947.400 444.900 948.600 445.650 ;
        RECT 946.950 442.800 949.050 444.900 ;
        RECT 943.950 439.950 946.050 442.050 ;
        RECT 950.100 440.700 951.000 446.100 ;
        RECT 951.900 444.300 954.000 445.200 ;
        RECT 959.700 444.300 960.600 453.300 ;
        RECT 968.400 451.200 969.450 460.950 ;
        RECT 961.950 449.100 964.050 451.200 ;
        RECT 967.950 449.100 970.050 451.200 ;
        RECT 962.400 448.350 963.600 449.100 ;
        RECT 961.800 445.950 963.900 448.050 ;
        RECT 951.900 443.100 960.600 444.300 ;
        RECT 944.400 427.050 945.450 439.950 ;
        RECT 949.800 438.600 951.900 440.700 ;
        RECT 953.100 440.100 955.200 442.200 ;
        RECT 957.000 441.300 959.100 443.100 ;
        RECT 964.950 442.800 967.050 444.900 ;
        RECT 961.950 439.950 964.050 442.050 ;
        RECT 953.400 437.550 954.600 439.800 ;
        RECT 943.950 424.950 946.050 427.050 ;
        RECT 953.400 421.050 954.450 437.550 ;
        RECT 962.400 433.050 963.450 439.950 ;
        RECT 961.950 430.950 964.050 433.050 ;
        RECT 958.950 424.950 961.050 427.050 ;
        RECT 952.950 418.950 955.050 421.050 ;
        RECT 940.950 415.950 943.050 418.050 ;
        RECT 946.950 416.100 949.050 418.200 ;
        RECT 947.400 415.350 948.600 416.100 ;
        RECT 943.950 412.950 946.050 415.050 ;
        RECT 946.950 412.950 949.050 415.050 ;
        RECT 949.950 412.950 952.050 415.050 ;
        RECT 940.950 409.950 943.050 412.050 ;
        RECT 944.400 410.400 945.600 412.650 ;
        RECT 950.400 412.050 951.600 412.650 ;
        RECT 959.400 412.050 960.450 424.950 ;
        RECT 965.400 421.050 966.450 442.800 ;
        RECT 967.950 430.950 970.050 436.050 ;
        RECT 971.400 430.050 972.450 464.400 ;
        RECT 970.950 427.950 973.050 430.050 ;
        RECT 970.950 421.950 973.050 424.050 ;
        RECT 964.950 417.000 967.050 421.050 ;
        RECT 971.400 418.200 972.450 421.950 ;
        RECT 965.400 415.350 966.600 417.000 ;
        RECT 970.950 416.100 973.050 418.200 ;
        RECT 974.400 418.050 975.450 472.950 ;
        RECT 977.400 436.050 978.450 481.950 ;
        RECT 982.950 475.950 985.050 478.050 ;
        RECT 983.400 460.050 984.450 475.950 ;
        RECT 986.400 460.050 987.450 496.950 ;
        RECT 989.400 475.050 990.450 506.400 ;
        RECT 991.950 502.950 994.050 505.050 ;
        RECT 992.400 496.050 993.450 502.950 ;
        RECT 995.400 499.050 996.450 550.950 ;
        RECT 1000.950 547.800 1003.050 549.900 ;
        RECT 997.950 529.950 1000.050 532.050 ;
        RECT 998.400 516.450 999.450 529.950 ;
        RECT 1001.400 529.050 1002.450 547.800 ;
        RECT 1007.400 535.050 1008.450 565.950 ;
        RECT 1012.950 565.800 1015.050 567.900 ;
        RECT 1018.950 565.950 1021.050 568.050 ;
        RECT 1012.950 556.950 1015.050 559.050 ;
        RECT 1006.950 532.950 1009.050 535.050 ;
        RECT 1000.950 526.950 1003.050 529.050 ;
        RECT 1006.950 528.000 1009.050 531.900 ;
        RECT 1013.400 528.600 1014.450 556.950 ;
        RECT 1007.400 526.350 1008.600 528.000 ;
        RECT 1013.400 526.350 1014.600 528.600 ;
        RECT 1003.950 523.950 1006.050 526.050 ;
        RECT 1006.950 523.950 1009.050 526.050 ;
        RECT 1009.950 523.950 1012.050 526.050 ;
        RECT 1012.950 523.950 1015.050 526.050 ;
        RECT 1004.400 521.400 1005.600 523.650 ;
        RECT 1010.400 522.900 1011.600 523.650 ;
        RECT 1004.400 517.050 1005.450 521.400 ;
        RECT 1009.950 520.800 1012.050 522.900 ;
        RECT 1015.950 520.950 1018.050 523.050 ;
        RECT 1012.950 517.950 1015.050 520.050 ;
        RECT 998.400 515.400 1002.450 516.450 ;
        RECT 997.950 511.950 1000.050 514.050 ;
        RECT 994.950 496.950 997.050 499.050 ;
        RECT 991.950 493.950 994.050 496.050 ;
        RECT 998.400 495.600 999.450 511.950 ;
        RECT 1001.400 508.050 1002.450 515.400 ;
        RECT 1003.950 514.950 1006.050 517.050 ;
        RECT 1009.950 514.950 1012.050 517.050 ;
        RECT 1000.950 505.950 1003.050 508.050 ;
        RECT 998.400 493.350 999.600 495.600 ;
        RECT 1003.950 494.100 1006.050 496.200 ;
        RECT 1004.400 493.350 1005.600 494.100 ;
        RECT 994.950 490.950 997.050 493.050 ;
        RECT 997.950 490.950 1000.050 493.050 ;
        RECT 1000.950 490.950 1003.050 493.050 ;
        RECT 1003.950 490.950 1006.050 493.050 ;
        RECT 991.950 487.950 994.050 490.050 ;
        RECT 995.400 488.400 996.600 490.650 ;
        RECT 1001.400 489.900 1002.600 490.650 ;
        RECT 1010.400 489.900 1011.450 514.950 ;
        RECT 988.950 472.950 991.050 475.050 ;
        RECT 992.400 466.050 993.450 487.950 ;
        RECT 995.400 481.050 996.450 488.400 ;
        RECT 1000.950 487.800 1003.050 489.900 ;
        RECT 1009.950 487.800 1012.050 489.900 ;
        RECT 994.950 478.950 997.050 481.050 ;
        RECT 1000.950 480.450 1005.000 481.050 ;
        RECT 1000.950 480.000 1005.450 480.450 ;
        RECT 1000.950 478.950 1006.050 480.000 ;
        RECT 995.400 472.050 996.450 478.950 ;
        RECT 1003.950 475.950 1006.050 478.950 ;
        RECT 1013.400 478.050 1014.450 517.950 ;
        RECT 1016.400 514.050 1017.450 520.950 ;
        RECT 1015.950 511.950 1018.050 514.050 ;
        RECT 1015.950 505.950 1018.050 508.050 ;
        RECT 1012.950 475.950 1015.050 478.050 ;
        RECT 1016.400 472.050 1017.450 505.950 ;
        RECT 1019.400 495.450 1020.450 565.950 ;
        RECT 1022.400 508.050 1023.450 620.400 ;
        RECT 1024.950 610.950 1027.050 613.050 ;
        RECT 1028.400 606.600 1029.450 751.950 ;
        RECT 1030.950 730.950 1033.050 733.050 ;
        RECT 1031.400 654.450 1032.450 730.950 ;
        RECT 1034.400 730.050 1035.450 755.400 ;
        RECT 1036.950 745.950 1039.050 748.050 ;
        RECT 1033.950 727.950 1036.050 730.050 ;
        RECT 1033.950 724.800 1036.050 726.900 ;
        RECT 1034.400 661.050 1035.450 724.800 ;
        RECT 1033.950 658.950 1036.050 661.050 ;
        RECT 1031.400 653.400 1035.450 654.450 ;
        RECT 1034.400 607.050 1035.450 653.400 ;
        RECT 1037.400 622.050 1038.450 745.950 ;
        RECT 1040.400 685.200 1041.450 781.950 ;
        RECT 1043.400 769.050 1044.450 799.950 ;
        RECT 1042.950 766.950 1045.050 769.050 ;
        RECT 1042.950 763.800 1045.050 765.900 ;
        RECT 1043.400 721.050 1044.450 763.800 ;
        RECT 1042.950 718.950 1045.050 721.050 ;
        RECT 1039.950 683.100 1042.050 685.200 ;
        RECT 1036.950 619.950 1039.050 622.050 ;
        RECT 1036.950 610.950 1039.050 613.050 ;
        RECT 1028.400 604.350 1029.600 606.600 ;
        RECT 1033.950 604.950 1036.050 607.050 ;
        RECT 1027.950 601.950 1030.050 604.050 ;
        RECT 1030.950 601.950 1033.050 604.050 ;
        RECT 1024.950 598.950 1027.050 601.050 ;
        RECT 1031.400 600.000 1032.600 601.650 ;
        RECT 1025.400 550.050 1026.450 598.950 ;
        RECT 1030.950 595.950 1033.050 600.000 ;
        RECT 1033.950 598.950 1036.050 601.050 ;
        RECT 1034.400 592.050 1035.450 598.950 ;
        RECT 1033.950 589.950 1036.050 592.050 ;
        RECT 1037.400 580.050 1038.450 610.950 ;
        RECT 1040.400 598.050 1041.450 683.100 ;
        RECT 1042.950 619.950 1045.050 622.050 ;
        RECT 1039.950 595.950 1042.050 598.050 ;
        RECT 1043.400 586.050 1044.450 619.950 ;
        RECT 1042.950 583.950 1045.050 586.050 ;
        RECT 1039.950 580.950 1042.050 583.050 ;
        RECT 1036.950 577.950 1039.050 580.050 ;
        RECT 1027.950 571.950 1030.050 574.050 ;
        RECT 1036.800 572.100 1038.900 574.200 ;
        RECT 1040.400 574.050 1041.450 580.950 ;
        RECT 1024.950 547.950 1027.050 550.050 ;
        RECT 1028.400 540.450 1029.450 571.950 ;
        RECT 1037.400 571.350 1038.600 572.100 ;
        RECT 1039.950 571.950 1042.050 574.050 ;
        RECT 1033.950 568.950 1036.050 571.050 ;
        RECT 1036.950 568.950 1039.050 571.050 ;
        RECT 1030.950 565.950 1033.050 568.050 ;
        RECT 1034.400 566.400 1035.600 568.650 ;
        RECT 1025.400 539.400 1029.450 540.450 ;
        RECT 1025.400 520.050 1026.450 539.400 ;
        RECT 1031.400 537.450 1032.450 565.950 ;
        RECT 1034.400 547.050 1035.450 566.400 ;
        RECT 1039.950 565.950 1042.050 568.050 ;
        RECT 1040.400 549.450 1041.450 565.950 ;
        RECT 1037.400 548.400 1041.450 549.450 ;
        RECT 1033.950 544.950 1036.050 547.050 ;
        RECT 1028.400 536.400 1032.450 537.450 ;
        RECT 1028.400 529.050 1029.450 536.400 ;
        RECT 1030.950 532.950 1033.050 535.050 ;
        RECT 1027.950 526.950 1030.050 529.050 ;
        RECT 1031.400 528.600 1032.450 532.950 ;
        RECT 1037.400 528.600 1038.450 548.400 ;
        RECT 1043.400 546.450 1044.450 583.950 ;
        RECT 1040.400 545.400 1044.450 546.450 ;
        RECT 1040.400 529.050 1041.450 545.400 ;
        RECT 1031.400 526.350 1032.600 528.600 ;
        RECT 1037.400 526.350 1038.600 528.600 ;
        RECT 1039.800 526.950 1041.900 529.050 ;
        RECT 1030.950 523.950 1033.050 526.050 ;
        RECT 1033.950 523.950 1036.050 526.050 ;
        RECT 1036.950 523.950 1039.050 526.050 ;
        RECT 1042.950 523.800 1045.050 525.900 ;
        RECT 1027.950 520.950 1030.050 523.050 ;
        RECT 1034.400 522.900 1035.600 523.650 ;
        RECT 1024.950 517.950 1027.050 520.050 ;
        RECT 1021.950 505.950 1024.050 508.050 ;
        RECT 1021.950 495.450 1024.050 496.200 ;
        RECT 1028.400 496.050 1029.450 520.950 ;
        RECT 1033.950 520.800 1036.050 522.900 ;
        RECT 1043.400 517.050 1044.450 523.800 ;
        RECT 1042.950 514.950 1045.050 517.050 ;
        RECT 1030.950 505.950 1033.050 508.050 ;
        RECT 1019.400 494.400 1024.050 495.450 ;
        RECT 1021.950 494.100 1024.050 494.400 ;
        RECT 1022.400 493.350 1023.600 494.100 ;
        RECT 1027.950 493.950 1030.050 496.050 ;
        RECT 1021.950 490.950 1024.050 493.050 ;
        RECT 1024.950 490.950 1027.050 493.050 ;
        RECT 1025.400 488.400 1026.600 490.650 ;
        RECT 994.950 469.950 997.050 472.050 ;
        RECT 1003.950 469.950 1006.050 472.050 ;
        RECT 1015.950 469.950 1018.050 472.050 ;
        RECT 991.950 463.950 994.050 466.050 ;
        RECT 982.800 457.950 984.900 460.050 ;
        RECT 985.950 457.950 988.050 460.050 ;
        RECT 1000.950 457.950 1003.050 460.050 ;
        RECT 982.800 454.500 984.900 456.600 ;
        RECT 980.100 445.950 982.200 448.050 ;
        RECT 983.100 447.300 984.300 454.500 ;
        RECT 986.400 451.350 987.600 453.600 ;
        RECT 992.400 453.300 994.500 455.400 ;
        RECT 986.100 448.950 988.200 451.050 ;
        RECT 989.100 449.700 991.200 451.800 ;
        RECT 989.100 447.300 990.000 449.700 ;
        RECT 983.100 446.100 990.000 447.300 ;
        RECT 980.400 444.900 981.600 445.650 ;
        RECT 979.950 442.800 982.050 444.900 ;
        RECT 983.100 440.700 984.000 446.100 ;
        RECT 984.900 444.300 987.000 445.200 ;
        RECT 992.700 444.300 993.600 453.300 ;
        RECT 995.400 450.450 996.600 450.600 ;
        RECT 995.400 449.400 999.450 450.450 ;
        RECT 995.400 448.350 996.600 449.400 ;
        RECT 994.800 445.950 996.900 448.050 ;
        RECT 984.900 443.100 993.600 444.300 ;
        RECT 982.800 438.600 984.900 440.700 ;
        RECT 986.100 440.100 988.200 442.200 ;
        RECT 990.000 441.300 992.100 443.100 ;
        RECT 986.400 438.000 987.600 439.800 ;
        RECT 976.950 433.950 979.050 436.050 ;
        RECT 985.950 433.950 988.050 438.000 ;
        RECT 998.400 436.050 999.450 449.400 ;
        RECT 997.950 433.950 1000.050 436.050 ;
        RECT 971.400 415.350 972.600 416.100 ;
        RECT 973.950 415.950 976.050 418.050 ;
        RECT 964.950 412.950 967.050 415.050 ;
        RECT 967.950 412.950 970.050 415.050 ;
        RECT 970.950 412.950 973.050 415.050 ;
        RECT 950.400 410.400 955.050 412.050 ;
        RECT 941.400 375.450 942.450 409.950 ;
        RECT 944.400 400.050 945.450 410.400 ;
        RECT 951.000 409.950 955.050 410.400 ;
        RECT 955.950 409.950 958.050 412.050 ;
        RECT 958.950 409.950 961.050 412.050 ;
        RECT 968.400 410.400 969.600 412.650 ;
        RECT 956.400 406.050 957.450 409.950 ;
        RECT 955.950 403.950 958.050 406.050 ;
        RECT 961.950 400.950 964.050 403.050 ;
        RECT 943.950 397.950 946.050 400.050 ;
        RECT 949.950 397.950 952.050 400.050 ;
        RECT 944.400 394.050 945.450 397.950 ;
        RECT 943.950 391.950 946.050 394.050 ;
        RECT 941.400 374.400 945.450 375.450 ;
        RECT 934.950 370.950 937.050 373.050 ;
        RECT 937.950 371.100 940.050 373.200 ;
        RECT 944.400 372.600 945.450 374.400 ;
        RECT 950.400 373.050 951.450 397.950 ;
        RECT 958.950 391.950 961.050 394.050 ;
        RECT 955.950 382.950 958.050 385.050 ;
        RECT 938.400 370.350 939.600 371.100 ;
        RECT 944.400 370.350 945.600 372.600 ;
        RECT 949.950 370.950 952.050 373.050 ;
        RECT 952.950 370.950 955.050 373.050 ;
        RECT 937.950 367.950 940.050 370.050 ;
        RECT 940.950 367.950 943.050 370.050 ;
        RECT 943.950 367.950 946.050 370.050 ;
        RECT 946.950 367.950 949.050 370.050 ;
        RECT 941.400 366.900 942.600 367.650 ;
        RECT 940.950 364.800 943.050 366.900 ;
        RECT 947.400 365.400 948.600 367.650 ;
        RECT 943.950 361.950 946.050 364.050 ;
        RECT 940.950 349.950 943.050 352.050 ;
        RECT 937.950 340.950 940.050 343.050 ;
        RECT 932.400 338.400 936.450 339.450 ;
        RECT 914.400 325.050 915.450 337.950 ;
        RECT 920.400 337.350 921.600 338.100 ;
        RECT 926.400 337.350 927.600 338.100 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 928.950 334.950 931.050 337.050 ;
        RECT 923.400 332.400 924.600 334.650 ;
        RECT 929.400 333.000 930.600 334.650 ;
        RECT 913.950 322.950 916.050 325.050 ;
        RECT 910.950 319.950 913.050 322.050 ;
        RECT 916.950 319.950 919.050 322.050 ;
        RECT 917.400 304.050 918.450 319.950 ;
        RECT 919.950 313.950 922.050 316.050 ;
        RECT 920.400 310.050 921.450 313.950 ;
        RECT 923.400 313.050 924.450 332.400 ;
        RECT 928.950 328.950 931.050 333.000 ;
        RECT 931.950 331.950 934.050 334.050 ;
        RECT 922.950 310.950 925.050 313.050 ;
        RECT 919.950 307.950 922.050 310.050 ;
        RECT 928.950 304.950 931.050 307.050 ;
        RECT 916.950 301.950 919.050 304.050 ;
        RECT 901.950 298.950 904.050 301.050 ;
        RECT 907.950 298.950 910.050 301.050 ;
        RECT 890.400 292.350 891.600 294.000 ;
        RECT 896.400 292.350 897.600 294.000 ;
        RECT 898.950 292.950 901.050 295.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 892.950 289.950 895.050 292.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 887.400 288.000 888.600 289.650 ;
        RECT 886.950 283.950 889.050 288.000 ;
        RECT 893.400 287.400 894.600 289.650 ;
        RECT 878.400 281.400 882.450 282.450 ;
        RECT 875.400 256.350 876.600 258.600 ;
        RECT 874.800 253.950 876.900 256.050 ;
        RECT 878.400 253.050 879.450 281.400 ;
        RECT 893.400 280.050 894.450 287.400 ;
        RECT 892.950 277.950 895.050 280.050 ;
        RECT 892.950 265.950 895.050 268.050 ;
        RECT 886.950 259.950 889.050 262.050 ;
        RECT 883.950 257.100 886.050 259.200 ;
        RECT 884.400 256.350 885.600 257.100 ;
        RECT 883.800 253.950 885.900 256.050 ;
        RECT 869.400 251.400 873.450 252.450 ;
        RECT 865.200 247.500 867.300 249.600 ;
        RECT 865.200 242.700 866.700 247.500 ;
        RECT 865.200 240.600 867.300 242.700 ;
        RECT 844.950 229.950 847.050 232.050 ;
        RECT 826.950 220.950 829.050 223.050 ;
        RECT 838.950 220.950 841.050 223.050 ;
        RECT 823.950 218.100 826.050 220.200 ;
        RECT 824.400 213.450 825.450 218.100 ;
        RECT 827.100 214.950 829.200 217.050 ;
        RECT 833.100 214.950 835.200 217.050 ;
        RECT 827.400 213.450 828.600 214.650 ;
        RECT 824.400 212.400 828.600 213.450 ;
        RECT 820.500 207.300 822.600 209.400 ;
        RECT 820.500 203.700 821.700 207.300 ;
        RECT 814.200 201.600 816.300 203.700 ;
        RECT 817.200 201.600 819.300 203.700 ;
        RECT 820.200 201.600 822.300 203.700 ;
        RECT 839.400 196.050 840.450 220.950 ;
        RECT 845.400 208.050 846.450 229.950 ;
        RECT 856.950 223.950 859.050 226.050 ;
        RECT 857.400 216.600 858.450 223.950 ;
        RECT 862.950 218.100 865.050 220.200 ;
        RECT 863.400 217.350 864.600 218.100 ;
        RECT 857.400 214.350 858.600 216.600 ;
        RECT 862.800 214.950 864.900 217.050 ;
        RECT 868.800 214.950 870.900 217.050 ;
        RECT 853.950 211.950 856.050 214.050 ;
        RECT 856.950 211.950 859.050 214.050 ;
        RECT 854.400 210.000 855.600 211.650 ;
        RECT 844.950 205.950 847.050 208.050 ;
        RECT 853.950 205.950 856.050 210.000 ;
        RECT 872.400 196.050 873.450 251.400 ;
        RECT 877.950 250.950 880.050 253.050 ;
        RECT 875.400 228.300 878.400 230.400 ;
        RECT 879.300 228.300 881.400 230.400 ;
        RECT 875.400 209.400 876.900 228.300 ;
        RECT 879.300 222.300 880.500 228.300 ;
        RECT 878.400 220.200 880.500 222.300 ;
        RECT 875.400 207.300 877.500 209.400 ;
        RECT 876.300 203.700 877.500 207.300 ;
        RECT 879.300 203.700 880.500 220.200 ;
        RECT 881.700 225.300 883.800 227.400 ;
        RECT 881.700 203.700 882.900 225.300 ;
        RECT 887.400 217.200 888.450 259.950 ;
        RECT 893.400 238.050 894.450 265.950 ;
        RECT 902.400 262.050 903.450 298.950 ;
        RECT 904.950 295.950 907.050 298.050 ;
        RECT 909.000 297.900 912.000 298.050 ;
        RECT 907.950 297.450 912.000 297.900 ;
        RECT 907.950 297.000 912.450 297.450 ;
        RECT 907.950 295.950 913.050 297.000 ;
        RECT 901.950 259.950 904.050 262.050 ;
        RECT 905.400 261.600 906.450 295.950 ;
        RECT 907.950 295.800 910.050 295.950 ;
        RECT 908.400 268.050 909.450 295.800 ;
        RECT 910.950 292.950 913.050 295.950 ;
        RECT 917.400 294.600 918.450 301.950 ;
        RECT 922.950 298.950 925.050 301.050 ;
        RECT 923.400 294.600 924.450 298.950 ;
        RECT 917.400 292.350 918.600 294.600 ;
        RECT 923.400 292.350 924.600 294.600 ;
        RECT 913.950 289.950 916.050 292.050 ;
        RECT 916.950 289.950 919.050 292.050 ;
        RECT 919.950 289.950 922.050 292.050 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 914.400 288.900 915.600 289.650 ;
        RECT 913.950 286.800 916.050 288.900 ;
        RECT 920.400 287.400 921.600 289.650 ;
        RECT 907.950 265.950 910.050 268.050 ;
        RECT 914.400 264.450 915.450 286.800 ;
        RECT 920.400 265.050 921.450 287.400 ;
        RECT 925.950 283.950 928.050 286.050 ;
        RECT 926.400 274.050 927.450 283.950 ;
        RECT 925.950 271.950 928.050 274.050 ;
        RECT 914.400 263.400 918.450 264.450 ;
        RECT 905.400 259.350 906.600 261.600 ;
        RECT 910.950 260.100 913.050 262.200 ;
        RECT 917.400 261.450 918.450 263.400 ;
        RECT 919.950 262.950 922.050 265.050 ;
        RECT 917.400 260.400 921.450 261.450 ;
        RECT 911.400 259.350 912.600 260.100 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 904.950 256.950 907.050 259.050 ;
        RECT 907.950 256.950 910.050 259.050 ;
        RECT 910.950 256.950 913.050 259.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 899.400 250.050 900.450 256.950 ;
        RECT 908.400 255.900 909.600 256.650 ;
        RECT 907.950 253.800 910.050 255.900 ;
        RECT 914.400 255.000 915.600 256.650 ;
        RECT 913.950 252.450 916.050 255.000 ;
        RECT 913.950 251.400 918.450 252.450 ;
        RECT 913.950 250.950 916.050 251.400 ;
        RECT 898.950 247.950 901.050 250.050 ;
        RECT 892.950 235.950 895.050 238.050 ;
        RECT 893.400 232.050 894.450 235.950 ;
        RECT 892.950 229.950 895.050 232.050 ;
        RECT 898.200 228.300 900.300 230.400 ;
        RECT 890.400 223.800 892.500 225.900 ;
        RECT 895.800 225.300 897.900 227.400 ;
        RECT 890.400 217.200 891.300 223.800 ;
        RECT 896.100 218.100 897.300 225.300 ;
        RECT 898.800 223.500 900.300 228.300 ;
        RECT 901.200 225.300 903.300 230.400 ;
        RECT 898.800 221.400 900.900 223.500 ;
        RECT 886.950 215.100 889.050 217.200 ;
        RECT 890.400 215.100 892.500 217.200 ;
        RECT 895.800 216.000 897.900 218.100 ;
        RECT 886.950 211.950 889.050 214.050 ;
        RECT 887.400 211.350 888.600 211.950 ;
        RECT 886.800 208.950 888.900 211.050 ;
        RECT 890.400 204.600 891.300 215.100 ;
        RECT 893.100 208.500 895.200 210.600 ;
        RECT 875.700 201.600 877.800 203.700 ;
        RECT 878.700 201.600 880.800 203.700 ;
        RECT 881.700 201.600 883.800 203.700 ;
        RECT 889.800 202.500 891.900 204.600 ;
        RECT 896.100 203.700 897.300 216.000 ;
        RECT 898.800 203.700 900.300 221.400 ;
        RECT 902.100 203.700 903.300 225.300 ;
        RECT 895.200 201.600 897.300 203.700 ;
        RECT 898.200 201.600 900.300 203.700 ;
        RECT 901.200 201.600 903.300 203.700 ;
        RECT 904.200 228.300 906.300 230.400 ;
        RECT 904.200 223.500 905.700 228.300 ;
        RECT 904.200 221.400 906.300 223.500 ;
        RECT 904.200 203.700 905.700 221.400 ;
        RECT 913.800 214.950 915.900 217.050 ;
        RECT 910.950 211.950 913.050 214.050 ;
        RECT 914.400 213.000 915.600 214.650 ;
        RECT 904.200 201.600 906.300 203.700 ;
        RECT 817.950 193.950 820.050 196.050 ;
        RECT 838.950 193.950 841.050 196.050 ;
        RECT 871.950 193.950 874.050 196.050 ;
        RECT 892.950 193.950 895.050 196.050 ;
        RECT 907.950 193.950 910.050 196.050 ;
        RECT 793.950 182.100 796.050 184.200 ;
        RECT 794.400 181.350 795.600 182.100 ;
        RECT 799.950 181.950 802.050 184.050 ;
        RECT 805.950 182.100 808.050 184.200 ;
        RECT 811.950 182.100 814.050 184.200 ;
        RECT 818.400 183.600 819.450 193.950 ;
        RECT 838.950 187.950 841.050 190.050 ;
        RECT 842.700 189.300 844.800 191.400 ;
        RECT 800.400 181.050 801.450 181.950 ;
        RECT 802.950 181.050 805.050 181.200 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 800.400 179.100 805.050 181.050 ;
        RECT 800.400 178.950 804.000 179.100 ;
        RECT 791.400 177.900 792.600 178.650 ;
        RECT 790.950 175.800 793.050 177.900 ;
        RECT 796.950 145.950 799.050 148.050 ;
        RECT 797.400 138.600 798.450 145.950 ;
        RECT 800.400 141.450 801.450 178.950 ;
        RECT 806.400 169.050 807.450 182.100 ;
        RECT 812.400 181.350 813.600 182.100 ;
        RECT 818.400 181.350 819.600 183.600 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 823.950 179.100 826.050 181.200 ;
        RECT 833.400 180.450 834.600 180.600 ;
        RECT 830.400 179.400 834.600 180.450 ;
        RECT 815.400 176.400 816.600 178.650 ;
        RECT 824.400 178.350 825.600 179.100 ;
        RECT 815.400 172.050 816.450 176.400 ;
        RECT 824.100 175.950 826.200 178.050 ;
        RECT 814.950 169.950 817.050 172.050 ;
        RECT 805.950 166.950 808.050 169.050 ;
        RECT 830.400 160.050 831.450 179.400 ;
        RECT 833.400 178.350 834.600 179.400 ;
        RECT 839.400 178.050 840.450 187.950 ;
        RECT 833.100 175.950 835.200 178.050 ;
        RECT 838.950 175.950 841.050 178.050 ;
        RECT 843.300 171.600 844.800 189.300 ;
        RECT 842.700 169.500 844.800 171.600 ;
        RECT 843.300 164.700 844.800 169.500 ;
        RECT 842.700 162.600 844.800 164.700 ;
        RECT 845.700 189.300 847.800 191.400 ;
        RECT 848.700 189.300 850.800 191.400 ;
        RECT 851.700 189.300 853.800 191.400 ;
        RECT 845.700 167.700 846.900 189.300 ;
        RECT 848.700 171.600 850.200 189.300 ;
        RECT 851.700 177.000 852.900 189.300 ;
        RECT 857.100 188.400 859.200 190.500 ;
        RECT 865.200 189.300 867.300 191.400 ;
        RECT 868.200 189.300 870.300 191.400 ;
        RECT 871.200 189.300 873.300 191.400 ;
        RECT 853.800 182.400 855.900 184.500 ;
        RECT 857.700 177.900 858.600 188.400 ;
        RECT 860.100 181.950 862.200 184.050 ;
        RECT 860.400 180.000 861.600 181.650 ;
        RECT 851.100 174.900 853.200 177.000 ;
        RECT 856.500 175.800 858.600 177.900 ;
        RECT 859.950 175.950 862.050 180.000 ;
        RECT 848.100 169.500 850.200 171.600 ;
        RECT 845.700 162.600 847.800 167.700 ;
        RECT 848.700 164.700 850.200 169.500 ;
        RECT 851.700 167.700 852.900 174.900 ;
        RECT 857.700 169.200 858.600 175.800 ;
        RECT 851.100 165.600 853.200 167.700 ;
        RECT 856.500 167.100 858.600 169.200 ;
        RECT 866.100 167.700 867.300 189.300 ;
        RECT 865.200 165.600 867.300 167.700 ;
        RECT 868.500 172.800 869.700 189.300 ;
        RECT 871.500 185.700 872.700 189.300 ;
        RECT 871.500 183.600 873.600 185.700 ;
        RECT 868.500 170.700 870.600 172.800 ;
        RECT 868.500 164.700 869.700 170.700 ;
        RECT 872.100 164.700 873.600 183.600 ;
        RECT 893.400 178.050 894.450 193.950 ;
        RECT 908.400 183.600 909.450 193.950 ;
        RECT 911.400 184.050 912.450 211.950 ;
        RECT 913.950 208.950 916.050 213.000 ;
        RECT 913.950 190.950 916.050 193.050 ;
        RECT 914.400 186.450 915.450 190.950 ;
        RECT 917.400 190.050 918.450 251.400 ;
        RECT 920.400 223.050 921.450 260.400 ;
        RECT 922.950 260.100 925.050 262.200 ;
        RECT 929.400 261.450 930.450 304.950 ;
        RECT 932.400 265.050 933.450 331.950 ;
        RECT 935.400 316.050 936.450 338.400 ;
        RECT 938.400 319.050 939.450 340.950 ;
        RECT 941.400 331.050 942.450 349.950 ;
        RECT 944.400 340.050 945.450 361.950 ;
        RECT 947.400 346.050 948.450 365.400 ;
        RECT 949.950 358.950 952.050 361.050 ;
        RECT 946.950 343.950 949.050 346.050 ;
        RECT 950.400 343.050 951.450 358.950 ;
        RECT 953.400 352.050 954.450 370.950 ;
        RECT 952.950 349.950 955.050 352.050 ;
        RECT 956.400 349.050 957.450 382.950 ;
        RECT 959.400 364.050 960.450 391.950 ;
        RECT 962.400 373.050 963.450 400.950 ;
        RECT 968.400 379.050 969.450 410.400 ;
        RECT 973.950 406.950 976.050 409.050 ;
        RECT 970.950 382.950 973.050 385.050 ;
        RECT 967.950 376.950 970.050 379.050 ;
        RECT 971.400 375.450 972.450 382.950 ;
        RECT 968.400 374.400 972.450 375.450 ;
        RECT 961.950 370.950 964.050 373.050 ;
        RECT 968.400 372.600 969.450 374.400 ;
        RECT 974.400 372.600 975.450 406.950 ;
        RECT 977.400 397.050 978.450 433.950 ;
        RECT 979.950 415.950 982.050 418.050 ;
        RECT 991.950 416.100 994.050 418.200 ;
        RECT 976.950 394.950 979.050 397.050 ;
        RECT 980.400 382.050 981.450 415.950 ;
        RECT 992.400 415.350 993.600 416.100 ;
        RECT 988.950 412.950 991.050 415.050 ;
        RECT 991.950 412.950 994.050 415.050 ;
        RECT 994.950 412.950 997.050 415.050 ;
        RECT 989.400 411.000 990.600 412.650 ;
        RECT 988.950 406.950 991.050 411.000 ;
        RECT 995.400 410.400 996.600 412.650 ;
        RECT 995.400 406.050 996.450 410.400 ;
        RECT 994.950 403.950 997.050 406.050 ;
        RECT 991.950 394.950 994.050 397.050 ;
        RECT 988.950 385.950 991.050 388.050 ;
        RECT 979.950 379.950 982.050 382.050 ;
        RECT 976.950 376.950 979.050 379.050 ;
        RECT 977.400 373.050 978.450 376.950 ;
        RECT 989.400 376.050 990.450 385.950 ;
        RECT 979.950 373.950 982.050 376.050 ;
        RECT 968.400 370.350 969.600 372.600 ;
        RECT 974.400 370.350 975.600 372.600 ;
        RECT 976.950 370.950 979.050 373.050 ;
        RECT 964.950 367.950 967.050 370.050 ;
        RECT 967.950 367.950 970.050 370.050 ;
        RECT 970.950 367.950 973.050 370.050 ;
        RECT 973.950 367.950 976.050 370.050 ;
        RECT 965.400 366.900 966.600 367.650 ;
        RECT 971.400 366.900 972.600 367.650 ;
        RECT 980.400 367.050 981.450 373.950 ;
        RECT 982.950 370.950 985.050 373.050 ;
        RECT 985.950 371.100 988.050 373.200 ;
        RECT 964.950 364.800 967.050 366.900 ;
        RECT 970.950 364.800 973.050 366.900 ;
        RECT 979.950 364.950 982.050 367.050 ;
        RECT 965.400 364.050 966.450 364.800 ;
        RECT 983.400 364.050 984.450 370.950 ;
        RECT 958.950 361.950 961.050 364.050 ;
        RECT 965.400 362.400 970.050 364.050 ;
        RECT 966.000 361.950 970.050 362.400 ;
        RECT 982.950 361.950 985.050 364.050 ;
        RECT 967.950 355.950 970.050 358.050 ;
        RECT 955.950 346.950 958.050 349.050 ;
        RECT 961.950 346.950 964.050 349.050 ;
        RECT 949.950 340.950 952.050 343.050 ;
        RECT 957.000 342.450 961.050 343.050 ;
        RECT 956.400 340.950 961.050 342.450 ;
        RECT 943.950 337.950 946.050 340.050 ;
        RECT 950.400 339.600 951.450 340.950 ;
        RECT 956.400 339.600 957.450 340.950 ;
        RECT 950.400 337.350 951.600 339.600 ;
        RECT 956.400 337.350 957.600 339.600 ;
        RECT 946.950 334.950 949.050 337.050 ;
        RECT 949.950 334.950 952.050 337.050 ;
        RECT 952.950 334.950 955.050 337.050 ;
        RECT 955.950 334.950 958.050 337.050 ;
        RECT 943.950 331.950 946.050 334.050 ;
        RECT 947.400 332.400 948.600 334.650 ;
        RECT 953.400 333.000 954.600 334.650 ;
        RECT 940.950 328.950 943.050 331.050 ;
        RECT 937.950 316.950 940.050 319.050 ;
        RECT 934.950 313.950 937.050 316.050 ;
        RECT 935.400 288.900 936.450 313.950 ;
        RECT 944.400 310.050 945.450 331.950 ;
        RECT 937.950 307.950 940.050 310.050 ;
        RECT 943.950 307.950 946.050 310.050 ;
        RECT 934.950 286.800 937.050 288.900 ;
        RECT 938.400 283.050 939.450 307.950 ;
        RECT 947.400 307.050 948.450 332.400 ;
        RECT 952.950 328.950 955.050 333.000 ;
        RECT 946.950 304.950 949.050 307.050 ;
        RECT 958.950 301.950 961.050 304.050 ;
        RECT 943.500 297.300 945.600 299.400 ;
        RECT 953.100 298.500 955.200 300.600 ;
        RECT 940.950 293.100 943.050 295.200 ;
        RECT 941.400 292.350 942.600 293.100 ;
        RECT 941.100 289.950 943.200 292.050 ;
        RECT 944.400 288.300 945.300 297.300 ;
        RECT 946.800 293.700 948.900 295.800 ;
        RECT 950.400 295.350 951.600 297.600 ;
        RECT 948.000 291.300 948.900 293.700 ;
        RECT 949.800 292.950 951.900 295.050 ;
        RECT 953.700 291.300 954.900 298.500 ;
        RECT 948.000 290.100 954.900 291.300 ;
        RECT 951.000 288.300 953.100 289.200 ;
        RECT 944.400 287.100 953.100 288.300 ;
        RECT 945.900 285.300 948.000 287.100 ;
        RECT 949.800 284.100 951.900 286.200 ;
        RECT 954.000 284.700 954.900 290.100 ;
        RECT 955.800 289.950 957.900 292.050 ;
        RECT 956.400 288.900 957.600 289.650 ;
        RECT 955.950 286.800 958.050 288.900 ;
        RECT 937.950 280.950 940.050 283.050 ;
        RECT 943.950 280.950 946.050 283.050 ;
        RECT 950.400 282.000 951.600 283.800 ;
        RECT 953.100 282.600 955.200 284.700 ;
        RECT 934.950 268.950 937.050 271.050 ;
        RECT 931.950 262.950 934.050 265.050 ;
        RECT 926.400 260.400 930.450 261.450 ;
        RECT 935.400 261.600 936.450 268.950 ;
        RECT 923.400 235.050 924.450 260.100 ;
        RECT 922.950 232.950 925.050 235.050 ;
        RECT 919.950 220.950 922.050 223.050 ;
        RECT 922.800 214.950 924.900 217.050 ;
        RECT 923.400 213.900 924.600 214.650 ;
        RECT 922.950 211.800 925.050 213.900 ;
        RECT 919.950 208.950 922.050 211.050 ;
        RECT 916.950 187.950 919.050 190.050 ;
        RECT 914.400 185.400 918.450 186.450 ;
        RECT 908.400 181.350 909.600 183.600 ;
        RECT 910.950 181.950 913.050 184.050 ;
        RECT 917.400 183.600 918.450 185.400 ;
        RECT 917.400 181.350 918.600 183.600 ;
        RECT 905.100 178.950 907.200 181.050 ;
        RECT 908.100 178.950 910.200 181.050 ;
        RECT 913.800 178.950 915.900 181.050 ;
        RECT 916.800 178.950 918.900 181.050 ;
        RECT 905.400 178.050 906.600 178.650 ;
        RECT 878.100 175.950 880.200 178.050 ;
        RECT 884.100 175.950 886.200 178.050 ;
        RECT 892.950 175.950 895.050 178.050 ;
        RECT 901.950 176.400 906.600 178.050 ;
        RECT 914.400 177.900 915.600 178.650 ;
        RECT 901.950 175.950 906.000 176.400 ;
        RECT 848.700 162.600 850.800 164.700 ;
        RECT 867.600 162.600 869.700 164.700 ;
        RECT 870.600 162.600 873.600 164.700 ;
        RECT 884.400 173.400 885.600 175.650 ;
        RECT 829.950 157.950 832.050 160.050 ;
        RECT 868.950 157.950 871.050 160.050 ;
        RECT 820.950 148.950 823.050 151.050 ;
        RECT 811.950 142.950 814.050 145.050 ;
        RECT 800.400 140.400 804.450 141.450 ;
        RECT 803.400 138.600 804.450 140.400 ;
        RECT 797.400 136.350 798.600 138.600 ;
        RECT 803.400 136.350 804.600 138.600 ;
        RECT 808.950 137.100 811.050 139.200 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 800.400 131.400 801.600 133.650 ;
        RECT 796.950 127.950 799.050 130.050 ;
        RECT 784.950 121.950 787.050 124.050 ;
        RECT 778.950 118.950 781.050 121.050 ;
        RECT 733.950 115.950 736.050 118.050 ;
        RECT 763.950 115.950 766.050 118.050 ;
        RECT 731.700 111.300 733.800 113.400 ;
        RECT 732.300 93.600 733.800 111.300 ;
        RECT 731.700 91.500 733.800 93.600 ;
        RECT 732.300 86.700 733.800 91.500 ;
        RECT 731.700 84.600 733.800 86.700 ;
        RECT 734.700 111.300 736.800 113.400 ;
        RECT 737.700 111.300 739.800 113.400 ;
        RECT 740.700 111.300 742.800 113.400 ;
        RECT 734.700 89.700 735.900 111.300 ;
        RECT 737.700 93.600 739.200 111.300 ;
        RECT 740.700 99.000 741.900 111.300 ;
        RECT 746.100 110.400 748.200 112.500 ;
        RECT 754.200 111.300 756.300 113.400 ;
        RECT 757.200 111.300 759.300 113.400 ;
        RECT 760.200 111.300 762.300 113.400 ;
        RECT 742.800 104.400 744.900 106.500 ;
        RECT 746.700 99.900 747.600 110.400 ;
        RECT 749.100 103.950 751.200 106.050 ;
        RECT 749.400 102.900 750.600 103.650 ;
        RECT 748.950 100.800 751.050 102.900 ;
        RECT 740.100 96.900 742.200 99.000 ;
        RECT 745.500 97.800 747.600 99.900 ;
        RECT 737.100 91.500 739.200 93.600 ;
        RECT 734.700 84.600 736.800 89.700 ;
        RECT 737.700 86.700 739.200 91.500 ;
        RECT 740.700 89.700 741.900 96.900 ;
        RECT 746.700 91.200 747.600 97.800 ;
        RECT 740.100 87.600 742.200 89.700 ;
        RECT 745.500 89.100 747.600 91.200 ;
        RECT 755.100 89.700 756.300 111.300 ;
        RECT 754.200 87.600 756.300 89.700 ;
        RECT 757.500 94.800 758.700 111.300 ;
        RECT 760.500 107.700 761.700 111.300 ;
        RECT 760.500 105.600 762.600 107.700 ;
        RECT 764.400 106.050 765.450 115.950 ;
        RECT 757.500 92.700 759.600 94.800 ;
        RECT 757.500 86.700 758.700 92.700 ;
        RECT 761.100 86.700 762.600 105.600 ;
        RECT 763.950 103.950 766.050 106.050 ;
        RECT 767.100 97.950 769.200 100.050 ;
        RECT 773.100 97.950 775.200 100.050 ;
        RECT 773.400 96.000 774.600 97.650 ;
        RECT 772.950 91.950 775.050 96.000 ;
        RECT 737.700 84.600 739.800 86.700 ;
        RECT 756.600 84.600 758.700 86.700 ;
        RECT 759.600 84.600 762.600 86.700 ;
        RECT 751.950 73.950 754.050 76.050 ;
        RECT 730.950 67.950 733.050 70.050 ;
        RECT 713.400 58.350 714.600 59.100 ;
        RECT 719.400 58.350 720.600 60.600 ;
        RECT 727.950 59.100 730.050 61.200 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 718.950 55.950 721.050 58.050 ;
        RECT 710.400 54.900 711.600 55.650 ;
        RECT 703.950 52.800 706.050 54.900 ;
        RECT 709.950 52.800 712.050 54.900 ;
        RECT 716.400 53.400 717.600 55.650 ;
        RECT 700.950 28.950 703.050 31.050 ;
        RECT 701.400 27.450 702.600 27.600 ;
        RECT 698.400 26.400 702.600 27.450 ;
        RECT 706.950 27.000 709.050 31.050 ;
        RECT 701.400 25.350 702.600 26.400 ;
        RECT 707.400 25.350 708.600 27.000 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 704.400 21.900 705.600 22.650 ;
        RECT 710.400 21.900 711.600 22.650 ;
        RECT 659.400 16.050 660.450 20.400 ;
        RECT 664.950 19.800 667.050 21.900 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 676.950 19.800 679.050 21.900 ;
        RECT 682.950 19.800 685.050 21.900 ;
        RECT 694.950 19.800 697.050 21.900 ;
        RECT 703.950 19.800 706.050 21.900 ;
        RECT 709.950 19.800 712.050 21.900 ;
        RECT 716.400 16.050 717.450 53.400 ;
        RECT 721.950 43.950 724.050 46.050 ;
        RECT 718.950 25.950 721.050 28.050 ;
        RECT 719.400 21.900 720.450 25.950 ;
        RECT 718.950 19.800 721.050 21.900 ;
        RECT 722.400 21.450 723.450 43.950 ;
        RECT 731.400 43.050 732.450 67.950 ;
        RECT 736.950 60.000 739.050 64.050 ;
        RECT 737.400 58.350 738.600 60.000 ;
        RECT 742.950 59.100 745.050 61.200 ;
        RECT 743.400 58.350 744.600 59.100 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 739.950 55.950 742.050 58.050 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 745.950 55.950 748.050 58.050 ;
        RECT 740.400 53.400 741.600 55.650 ;
        RECT 746.400 54.900 747.600 55.650 ;
        RECT 740.400 46.050 741.450 53.400 ;
        RECT 745.950 52.800 748.050 54.900 ;
        RECT 739.950 43.950 742.050 46.050 ;
        RECT 730.950 40.950 733.050 43.050 ;
        RECT 739.950 31.950 742.050 34.050 ;
        RECT 730.950 26.100 733.050 28.200 ;
        RECT 731.400 25.350 732.600 26.100 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 728.400 21.900 729.600 22.650 ;
        RECT 727.950 21.450 730.050 21.900 ;
        RECT 722.400 20.400 730.050 21.450 ;
        RECT 727.950 19.800 730.050 20.400 ;
        RECT 734.400 20.400 735.600 22.650 ;
        RECT 730.950 16.050 733.050 19.050 ;
        RECT 658.950 13.950 661.050 16.050 ;
        RECT 703.950 13.950 706.050 16.050 ;
        RECT 715.950 13.950 718.050 16.050 ;
        RECT 727.950 15.000 733.050 16.050 ;
        RECT 727.950 14.400 732.450 15.000 ;
        RECT 727.950 13.950 732.000 14.400 ;
        RECT 643.950 10.950 646.050 13.050 ;
        RECT 734.400 7.050 735.450 20.400 ;
        RECT 740.400 19.050 741.450 31.950 ;
        RECT 752.400 28.200 753.450 73.950 ;
        RECT 757.950 64.950 760.050 67.050 ;
        RECT 754.950 58.950 757.050 61.050 ;
        RECT 755.400 54.900 756.450 58.950 ;
        RECT 754.950 52.800 757.050 54.900 ;
        RECT 758.400 46.050 759.450 64.950 ;
        RECT 763.950 59.100 766.050 61.200 ;
        RECT 764.400 58.350 765.600 59.100 ;
        RECT 773.100 58.950 775.200 61.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 773.400 57.000 774.600 58.650 ;
        RECT 779.400 57.450 780.450 118.950 ;
        RECT 784.950 115.950 787.050 118.050 ;
        RECT 785.400 109.050 786.450 115.950 ;
        RECT 784.950 106.950 787.050 109.050 ;
        RECT 785.400 99.900 786.450 106.950 ;
        RECT 787.950 104.100 790.050 106.200 ;
        RECT 797.400 105.600 798.450 127.950 ;
        RECT 800.400 121.050 801.450 131.400 ;
        RECT 809.400 130.050 810.450 137.100 ;
        RECT 812.400 133.050 813.450 142.950 ;
        RECT 821.400 139.200 822.450 148.950 ;
        RECT 850.800 142.500 852.900 144.600 ;
        RECT 820.950 137.100 823.050 139.200 ;
        RECT 826.950 138.000 829.050 142.050 ;
        RECT 821.400 136.350 822.600 137.100 ;
        RECT 827.400 136.350 828.600 138.000 ;
        RECT 838.950 136.950 841.050 142.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 826.950 133.950 829.050 136.050 ;
        RECT 829.950 133.950 832.050 136.050 ;
        RECT 811.950 130.950 814.050 133.050 ;
        RECT 824.400 132.900 825.600 133.650 ;
        RECT 823.950 130.800 826.050 132.900 ;
        RECT 830.400 131.400 831.600 133.650 ;
        RECT 808.950 127.950 811.050 130.050 ;
        RECT 811.950 124.950 814.050 127.050 ;
        RECT 799.950 118.950 802.050 121.050 ;
        RECT 812.400 112.050 813.450 124.950 ;
        RECT 830.400 121.050 831.450 131.400 ;
        RECT 829.950 118.950 832.050 121.050 ;
        RECT 839.400 120.450 840.450 136.950 ;
        RECT 848.100 133.950 850.200 136.050 ;
        RECT 851.100 135.300 852.300 142.500 ;
        RECT 854.400 139.350 855.600 141.600 ;
        RECT 860.400 141.300 862.500 143.400 ;
        RECT 854.100 136.950 856.200 139.050 ;
        RECT 857.100 137.700 859.200 139.800 ;
        RECT 857.100 135.300 858.000 137.700 ;
        RECT 851.100 134.100 858.000 135.300 ;
        RECT 848.400 132.450 849.600 133.650 ;
        RECT 845.400 131.400 849.600 132.450 ;
        RECT 845.400 121.050 846.450 131.400 ;
        RECT 851.100 128.700 852.000 134.100 ;
        RECT 852.900 132.300 855.000 133.200 ;
        RECT 860.700 132.300 861.600 141.300 ;
        RECT 863.400 138.450 864.600 138.600 ;
        RECT 863.400 137.400 867.450 138.450 ;
        RECT 863.400 136.350 864.600 137.400 ;
        RECT 862.800 133.950 864.900 136.050 ;
        RECT 866.400 133.050 867.450 137.400 ;
        RECT 852.900 131.100 861.600 132.300 ;
        RECT 850.800 126.600 852.900 128.700 ;
        RECT 854.100 128.100 856.200 130.200 ;
        RECT 858.000 129.300 860.100 131.100 ;
        RECT 865.950 130.950 868.050 133.050 ;
        RECT 854.400 127.050 855.600 127.800 ;
        RECT 853.950 124.950 856.050 127.050 ;
        RECT 865.950 123.450 868.050 124.050 ;
        RECT 869.400 123.450 870.450 157.950 ;
        RECT 880.950 148.950 883.050 151.050 ;
        RECT 874.950 142.950 877.050 145.050 ;
        RECT 871.950 136.950 874.050 139.050 ;
        RECT 872.400 127.050 873.450 136.950 ;
        RECT 871.950 124.950 874.050 127.050 ;
        RECT 865.950 122.400 870.450 123.450 ;
        RECT 865.950 121.950 868.050 122.400 ;
        RECT 836.400 119.400 840.450 120.450 ;
        RECT 823.950 115.950 826.050 118.050 ;
        RECT 811.950 109.950 814.050 112.050 ;
        RECT 784.950 97.800 787.050 99.900 ;
        RECT 788.400 82.050 789.450 104.100 ;
        RECT 797.400 103.350 798.600 105.600 ;
        RECT 817.950 104.100 820.050 106.200 ;
        RECT 824.400 105.600 825.450 115.950 ;
        RECT 818.400 103.350 819.600 104.100 ;
        RECT 824.400 103.350 825.600 105.600 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 794.400 98.400 795.600 100.650 ;
        RECT 800.400 99.900 801.600 100.650 ;
        RECT 821.400 99.900 822.600 100.650 ;
        RECT 836.400 100.050 837.450 119.400 ;
        RECT 844.950 118.950 847.050 121.050 ;
        RECT 850.950 109.950 853.050 112.050 ;
        RECT 844.950 104.100 847.050 106.200 ;
        RECT 845.400 103.350 846.600 104.100 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 794.400 82.050 795.450 98.400 ;
        RECT 799.950 97.800 802.050 99.900 ;
        RECT 820.950 97.800 823.050 99.900 ;
        RECT 835.950 97.950 838.050 100.050 ;
        RECT 842.400 98.400 843.600 100.650 ;
        RECT 787.950 79.950 790.050 82.050 ;
        RECT 793.950 79.950 796.050 82.050 ;
        RECT 782.100 58.950 784.200 61.050 ;
        RECT 782.400 57.450 783.600 58.650 ;
        RECT 767.400 54.900 768.600 55.650 ;
        RECT 766.950 52.800 769.050 54.900 ;
        RECT 772.950 52.950 775.050 57.000 ;
        RECT 779.400 56.400 783.600 57.450 ;
        RECT 757.950 43.950 760.050 46.050 ;
        RECT 782.400 37.050 783.450 56.400 ;
        RECT 788.400 55.050 789.450 79.950 ;
        RECT 842.400 79.050 843.450 98.400 ;
        RECT 851.400 96.900 852.450 109.950 ;
        RECT 866.400 106.200 867.450 121.950 ;
        RECT 875.400 112.050 876.450 142.950 ;
        RECT 881.400 138.600 882.450 148.950 ;
        RECT 884.400 145.050 885.450 173.400 ;
        RECT 893.400 172.050 894.450 175.950 ;
        RECT 913.950 175.800 916.050 177.900 ;
        RECT 892.950 169.950 895.050 172.050 ;
        RECT 886.950 145.950 889.050 148.050 ;
        RECT 907.950 145.950 910.050 148.050 ;
        RECT 916.950 145.950 919.050 148.050 ;
        RECT 883.950 142.950 886.050 145.050 ;
        RECT 887.400 138.600 888.450 145.950 ;
        RECT 908.400 138.600 909.450 145.950 ;
        RECT 881.400 136.350 882.600 138.600 ;
        RECT 887.400 136.350 888.600 138.600 ;
        RECT 908.400 136.350 909.600 138.600 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 884.400 132.900 885.600 133.650 ;
        RECT 883.950 130.800 886.050 132.900 ;
        RECT 905.400 131.400 906.600 133.650 ;
        RECT 917.400 132.900 918.450 145.950 ;
        RECT 905.400 127.050 906.450 131.400 ;
        RECT 916.950 130.800 919.050 132.900 ;
        RECT 904.950 124.950 907.050 127.050 ;
        RECT 920.400 121.050 921.450 208.950 ;
        RECT 922.950 187.950 925.050 190.050 ;
        RECT 923.400 139.200 924.450 187.950 ;
        RECT 926.400 157.050 927.450 260.400 ;
        RECT 935.400 259.350 936.600 261.600 ;
        RECT 931.950 256.950 934.050 259.050 ;
        RECT 934.950 256.950 937.050 259.050 ;
        RECT 937.950 256.950 940.050 259.050 ;
        RECT 928.950 253.950 931.050 256.050 ;
        RECT 932.400 254.400 933.600 256.650 ;
        RECT 938.400 254.400 939.600 256.650 ;
        RECT 929.400 172.050 930.450 253.950 ;
        RECT 932.400 250.050 933.450 254.400 ;
        RECT 931.950 247.950 934.050 250.050 ;
        RECT 938.400 226.050 939.450 254.400 ;
        RECT 944.400 226.050 945.450 280.950 ;
        RECT 949.950 277.950 952.050 282.000 ;
        RECT 959.400 277.050 960.450 301.950 ;
        RECT 962.400 291.450 963.450 346.950 ;
        RECT 964.950 340.950 967.050 343.050 ;
        RECT 965.400 310.050 966.450 340.950 ;
        RECT 964.950 307.950 967.050 310.050 ;
        RECT 968.400 304.050 969.450 355.950 ;
        RECT 979.950 343.950 982.050 346.050 ;
        RECT 973.950 338.100 976.050 343.050 ;
        RECT 980.400 339.600 981.450 343.950 ;
        RECT 974.400 337.350 975.600 338.100 ;
        RECT 980.400 337.350 981.600 339.600 ;
        RECT 973.950 334.950 976.050 337.050 ;
        RECT 976.950 334.950 979.050 337.050 ;
        RECT 979.950 334.950 982.050 337.050 ;
        RECT 977.400 333.900 978.600 334.650 ;
        RECT 976.950 331.800 979.050 333.900 ;
        RECT 976.950 319.950 979.050 322.050 ;
        RECT 970.950 313.950 973.050 316.050 ;
        RECT 967.950 301.950 970.050 304.050 ;
        RECT 967.950 298.800 970.050 300.900 ;
        RECT 962.400 290.400 966.450 291.450 ;
        RECT 961.950 286.950 964.050 289.050 ;
        RECT 962.400 283.050 963.450 286.950 ;
        RECT 961.950 280.950 964.050 283.050 ;
        RECT 961.950 277.800 964.050 279.900 ;
        RECT 949.950 274.800 952.050 276.900 ;
        RECT 958.950 274.950 961.050 277.050 ;
        RECT 946.950 262.950 949.050 265.050 ;
        RECT 947.400 255.900 948.450 262.950 ;
        RECT 946.950 253.800 949.050 255.900 ;
        RECT 937.950 223.950 940.050 226.050 ;
        RECT 943.950 223.950 946.050 226.050 ;
        RECT 931.950 220.950 934.050 223.050 ;
        RECT 928.950 169.950 931.050 172.050 ;
        RECT 925.950 154.950 928.050 157.050 ;
        RECT 929.400 148.050 930.450 169.950 ;
        RECT 932.400 163.050 933.450 220.950 ;
        RECT 944.400 216.600 945.450 223.950 ;
        RECT 950.400 220.200 951.450 274.800 ;
        RECT 955.950 261.000 958.050 265.050 ;
        RECT 962.400 262.200 963.450 277.800 ;
        RECT 965.400 274.050 966.450 290.400 ;
        RECT 968.400 286.050 969.450 298.800 ;
        RECT 971.400 295.200 972.450 313.950 ;
        RECT 970.950 293.100 973.050 295.200 ;
        RECT 977.400 294.600 978.450 319.950 ;
        RECT 979.950 307.950 982.050 310.050 ;
        RECT 980.400 301.050 981.450 307.950 ;
        RECT 986.400 304.050 987.450 371.100 ;
        RECT 988.950 370.950 991.050 376.050 ;
        RECT 992.400 373.200 993.450 394.950 ;
        RECT 1001.400 376.050 1002.450 457.950 ;
        RECT 991.950 371.100 994.050 373.200 ;
        RECT 997.950 372.000 1000.050 376.050 ;
        RECT 1000.950 373.950 1003.050 376.050 ;
        RECT 1004.400 373.050 1005.450 469.950 ;
        RECT 1025.400 469.050 1026.450 488.400 ;
        RECT 1024.950 466.950 1027.050 469.050 ;
        RECT 1018.950 460.950 1021.050 463.050 ;
        RECT 1024.950 460.950 1027.050 463.050 ;
        RECT 1019.400 454.050 1020.450 460.950 ;
        RECT 1006.950 449.100 1009.050 451.200 ;
        RECT 1012.950 449.100 1015.050 451.200 ;
        RECT 1018.950 450.000 1021.050 454.050 ;
        RECT 1025.400 451.050 1026.450 460.950 ;
        RECT 1027.950 454.950 1030.050 457.050 ;
        RECT 1007.400 442.050 1008.450 449.100 ;
        RECT 1013.400 448.350 1014.600 449.100 ;
        RECT 1019.400 448.350 1020.600 450.000 ;
        RECT 1024.950 448.950 1027.050 451.050 ;
        RECT 1012.950 445.950 1015.050 448.050 ;
        RECT 1015.950 445.950 1018.050 448.050 ;
        RECT 1018.950 445.950 1021.050 448.050 ;
        RECT 1021.950 445.950 1024.050 448.050 ;
        RECT 1016.400 443.400 1017.600 445.650 ;
        RECT 1022.400 444.900 1023.600 445.650 ;
        RECT 1006.950 439.950 1009.050 442.050 ;
        RECT 1012.950 439.950 1015.050 442.050 ;
        RECT 1006.950 427.950 1009.050 430.050 ;
        RECT 992.400 370.350 993.600 371.100 ;
        RECT 998.400 370.350 999.600 372.000 ;
        RECT 1003.950 370.950 1006.050 373.050 ;
        RECT 991.950 367.950 994.050 370.050 ;
        RECT 994.950 367.950 997.050 370.050 ;
        RECT 997.950 367.950 1000.050 370.050 ;
        RECT 1000.950 367.950 1003.050 370.050 ;
        RECT 995.400 366.900 996.600 367.650 ;
        RECT 994.950 364.800 997.050 366.900 ;
        RECT 1001.400 365.400 1002.600 367.650 ;
        RECT 1001.400 361.050 1002.450 365.400 ;
        RECT 1003.950 364.950 1006.050 367.050 ;
        RECT 1000.950 358.950 1003.050 361.050 ;
        RECT 1004.400 358.050 1005.450 364.950 ;
        RECT 1003.950 355.950 1006.050 358.050 ;
        RECT 988.950 352.950 991.050 355.050 ;
        RECT 989.400 334.050 990.450 352.950 ;
        RECT 1007.400 352.050 1008.450 427.950 ;
        RECT 1013.400 417.600 1014.450 439.950 ;
        RECT 1016.400 436.050 1017.450 443.400 ;
        RECT 1021.950 442.800 1024.050 444.900 ;
        RECT 1024.950 442.950 1027.050 445.050 ;
        RECT 1028.400 444.900 1029.450 454.950 ;
        RECT 1015.950 433.950 1018.050 436.050 ;
        RECT 1013.400 415.350 1014.600 417.600 ;
        RECT 1018.950 416.100 1021.050 418.200 ;
        RECT 1025.400 418.050 1026.450 442.950 ;
        RECT 1027.950 442.800 1030.050 444.900 ;
        RECT 1019.400 415.350 1020.600 416.100 ;
        RECT 1024.950 415.950 1027.050 418.050 ;
        RECT 1012.950 412.950 1015.050 415.050 ;
        RECT 1015.950 412.950 1018.050 415.050 ;
        RECT 1018.950 412.950 1021.050 415.050 ;
        RECT 1021.950 412.950 1024.050 415.050 ;
        RECT 1016.400 411.900 1017.600 412.650 ;
        RECT 1015.950 409.800 1018.050 411.900 ;
        RECT 1022.400 410.400 1023.600 412.650 ;
        RECT 1009.950 403.950 1012.050 406.050 ;
        RECT 1010.400 367.050 1011.450 403.950 ;
        RECT 1016.400 397.050 1017.450 409.800 ;
        RECT 1022.400 406.050 1023.450 410.400 ;
        RECT 1024.950 409.950 1027.050 412.050 ;
        RECT 1021.950 403.950 1024.050 406.050 ;
        RECT 1015.950 394.950 1018.050 397.050 ;
        RECT 1025.400 394.050 1026.450 409.950 ;
        RECT 1024.950 391.950 1027.050 394.050 ;
        RECT 1012.950 376.950 1015.050 379.050 ;
        RECT 1024.950 376.950 1027.050 379.050 ;
        RECT 1009.950 364.950 1012.050 367.050 ;
        RECT 1013.400 355.050 1014.450 376.950 ;
        RECT 1018.950 372.000 1021.050 376.050 ;
        RECT 1025.400 372.600 1026.450 376.950 ;
        RECT 1028.400 376.050 1029.450 442.800 ;
        RECT 1031.400 403.050 1032.450 505.950 ;
        RECT 1036.950 493.950 1039.050 496.050 ;
        RECT 1033.950 463.950 1036.050 466.050 ;
        RECT 1030.950 400.950 1033.050 403.050 ;
        RECT 1027.950 373.950 1030.050 376.050 ;
        RECT 1019.400 370.350 1020.600 372.000 ;
        RECT 1025.400 370.350 1026.600 372.600 ;
        RECT 1034.400 370.050 1035.450 463.950 ;
        RECT 1037.400 463.050 1038.450 493.950 ;
        RECT 1036.950 460.950 1039.050 463.050 ;
        RECT 1036.950 451.950 1039.050 454.050 ;
        RECT 1037.400 385.050 1038.450 451.950 ;
        RECT 1043.400 400.050 1044.450 514.950 ;
        RECT 1042.950 397.950 1045.050 400.050 ;
        RECT 1036.950 382.950 1039.050 385.050 ;
        RECT 1018.950 367.950 1021.050 370.050 ;
        RECT 1021.950 367.950 1024.050 370.050 ;
        RECT 1024.950 367.950 1027.050 370.050 ;
        RECT 1027.950 367.950 1030.050 370.050 ;
        RECT 1033.950 367.950 1036.050 370.050 ;
        RECT 1022.400 366.900 1023.600 367.650 ;
        RECT 1028.400 366.900 1029.600 367.650 ;
        RECT 1021.950 364.800 1024.050 366.900 ;
        RECT 1027.950 364.800 1030.050 366.900 ;
        RECT 1033.950 364.800 1036.050 366.900 ;
        RECT 1015.950 358.950 1018.050 361.050 ;
        RECT 1012.950 352.950 1015.050 355.050 ;
        RECT 991.950 349.950 994.050 352.050 ;
        RECT 1006.950 349.950 1009.050 352.050 ;
        RECT 988.950 331.950 991.050 334.050 ;
        RECT 988.950 316.950 991.050 319.050 ;
        RECT 985.950 301.950 988.050 304.050 ;
        RECT 979.950 298.950 982.050 301.050 ;
        RECT 984.000 294.600 988.050 295.050 ;
        RECT 977.400 292.350 978.600 294.600 ;
        RECT 983.400 292.950 988.050 294.600 ;
        RECT 983.400 292.350 984.600 292.950 ;
        RECT 973.950 289.950 976.050 292.050 ;
        RECT 976.950 289.950 979.050 292.050 ;
        RECT 979.950 289.950 982.050 292.050 ;
        RECT 982.950 289.950 985.050 292.050 ;
        RECT 974.400 288.000 975.600 289.650 ;
        RECT 967.950 283.950 970.050 286.050 ;
        RECT 973.950 283.950 976.050 288.000 ;
        RECT 980.400 287.400 981.600 289.650 ;
        RECT 980.400 283.050 981.450 287.400 ;
        RECT 982.950 283.950 985.050 286.050 ;
        RECT 970.950 280.950 973.050 283.050 ;
        RECT 979.950 280.950 982.050 283.050 ;
        RECT 971.400 277.050 972.450 280.950 ;
        RECT 970.950 274.950 973.050 277.050 ;
        RECT 983.400 274.050 984.450 283.950 ;
        RECT 964.950 271.950 967.050 274.050 ;
        RECT 973.950 271.950 976.050 274.050 ;
        RECT 982.950 271.950 985.050 274.050 ;
        RECT 965.400 265.050 966.450 271.950 ;
        RECT 970.950 268.950 973.050 271.050 ;
        RECT 964.950 262.950 967.050 265.050 ;
        RECT 956.400 259.350 957.600 261.000 ;
        RECT 961.950 260.100 964.050 262.200 ;
        RECT 962.400 259.350 963.600 260.100 ;
        RECT 955.950 256.950 958.050 259.050 ;
        RECT 958.950 256.950 961.050 259.050 ;
        RECT 961.950 256.950 964.050 259.050 ;
        RECT 964.950 256.950 967.050 259.050 ;
        RECT 952.950 253.950 955.050 256.050 ;
        RECT 959.400 255.000 960.600 256.650 ;
        RECT 965.400 255.900 966.600 256.650 ;
        RECT 971.400 255.900 972.450 268.950 ;
        RECT 949.950 218.100 952.050 220.200 ;
        RECT 953.400 220.050 954.450 253.950 ;
        RECT 958.950 250.950 961.050 255.000 ;
        RECT 964.950 253.800 967.050 255.900 ;
        RECT 970.950 253.800 973.050 255.900 ;
        RECT 974.400 253.050 975.450 271.950 ;
        RECT 989.400 271.050 990.450 316.950 ;
        RECT 992.400 307.050 993.450 349.950 ;
        RECT 1012.950 343.950 1015.050 346.050 ;
        RECT 997.950 338.100 1000.050 340.200 ;
        RECT 1003.950 338.100 1006.050 340.200 ;
        RECT 1013.400 340.050 1014.450 343.950 ;
        RECT 998.400 337.350 999.600 338.100 ;
        RECT 1004.400 337.350 1005.600 338.100 ;
        RECT 1012.950 337.950 1015.050 340.050 ;
        RECT 997.950 334.950 1000.050 337.050 ;
        RECT 1000.950 334.950 1003.050 337.050 ;
        RECT 1003.950 334.950 1006.050 337.050 ;
        RECT 1006.950 334.950 1009.050 337.050 ;
        RECT 1001.400 333.900 1002.600 334.650 ;
        RECT 1000.950 331.800 1003.050 333.900 ;
        RECT 1013.400 316.050 1014.450 337.950 ;
        RECT 1012.950 313.950 1015.050 316.050 ;
        RECT 1009.950 310.950 1012.050 313.050 ;
        RECT 1010.400 307.050 1011.450 310.950 ;
        RECT 1016.400 307.050 1017.450 358.950 ;
        RECT 1018.950 352.950 1021.050 355.050 ;
        RECT 991.950 304.950 994.050 307.050 ;
        RECT 1009.950 304.950 1012.050 307.050 ;
        RECT 1015.950 304.950 1018.050 307.050 ;
        RECT 991.950 301.800 994.050 303.900 ;
        RECT 976.950 268.950 979.050 271.050 ;
        RECT 988.950 268.950 991.050 271.050 ;
        RECT 973.950 250.950 976.050 253.050 ;
        RECT 973.950 220.950 976.050 223.050 ;
        RECT 952.950 217.950 955.050 220.050 ;
        RECT 958.950 217.950 961.050 220.050 ;
        RECT 964.950 217.950 967.050 220.050 ;
        RECT 944.400 214.350 945.600 216.600 ;
        RECT 949.950 214.950 952.050 217.050 ;
        RECT 950.400 214.350 951.600 214.950 ;
        RECT 943.950 211.950 946.050 214.050 ;
        RECT 946.950 211.950 949.050 214.050 ;
        RECT 949.950 211.950 952.050 214.050 ;
        RECT 952.950 211.950 955.050 214.050 ;
        RECT 947.400 209.400 948.600 211.650 ;
        RECT 953.400 209.400 954.600 211.650 ;
        RECT 940.950 189.000 943.050 193.050 ;
        RECT 947.400 190.050 948.450 209.400 ;
        RECT 953.400 205.050 954.450 209.400 ;
        RECT 959.400 205.050 960.450 217.950 ;
        RECT 961.950 214.950 964.050 217.050 ;
        RECT 952.950 202.950 955.050 205.050 ;
        RECT 958.950 204.450 961.050 205.050 ;
        RECT 956.400 203.400 961.050 204.450 ;
        RECT 937.800 186.300 939.900 188.400 ;
        RECT 941.400 187.200 942.600 189.000 ;
        RECT 946.950 187.950 949.050 190.050 ;
        RECT 934.950 182.100 937.050 184.200 ;
        RECT 935.400 181.350 936.600 182.100 ;
        RECT 935.100 178.950 937.200 181.050 ;
        RECT 938.100 180.900 939.000 186.300 ;
        RECT 941.100 184.800 943.200 186.900 ;
        RECT 945.000 183.900 947.100 185.700 ;
        RECT 939.900 182.700 948.600 183.900 ;
        RECT 939.900 181.800 942.000 182.700 ;
        RECT 938.100 179.700 945.000 180.900 ;
        RECT 938.100 172.500 939.300 179.700 ;
        RECT 941.100 175.950 943.200 178.050 ;
        RECT 944.100 177.300 945.000 179.700 ;
        RECT 941.400 173.400 942.600 175.650 ;
        RECT 944.100 175.200 946.200 177.300 ;
        RECT 947.700 173.700 948.600 182.700 ;
        RECT 949.800 178.950 951.900 181.050 ;
        RECT 950.400 177.900 951.600 178.650 ;
        RECT 949.950 175.800 952.050 177.900 ;
        RECT 937.800 170.400 939.900 172.500 ;
        RECT 947.400 171.600 949.500 173.700 ;
        RECT 931.950 160.950 934.050 163.050 ;
        RECT 943.950 154.950 946.050 157.050 ;
        RECT 928.950 145.950 931.050 148.050 ;
        RECT 944.400 145.050 945.450 154.950 ;
        RECT 949.950 148.950 952.050 151.050 ;
        RECT 928.800 142.500 930.900 144.600 ;
        RECT 922.950 137.100 925.050 139.200 ;
        RECT 926.100 133.950 928.200 136.050 ;
        RECT 929.100 135.300 930.300 142.500 ;
        RECT 932.400 139.350 933.600 141.600 ;
        RECT 938.400 141.300 940.500 143.400 ;
        RECT 943.950 142.950 946.050 145.050 ;
        RECT 932.100 136.950 934.200 139.050 ;
        RECT 935.100 137.700 937.200 139.800 ;
        RECT 935.100 135.300 936.000 137.700 ;
        RECT 929.100 134.100 936.000 135.300 ;
        RECT 926.400 132.900 927.600 133.650 ;
        RECT 925.950 130.800 928.050 132.900 ;
        RECT 929.100 128.700 930.000 134.100 ;
        RECT 930.900 132.300 933.000 133.200 ;
        RECT 938.700 132.300 939.600 141.300 ;
        RECT 940.950 137.100 943.050 139.200 ;
        RECT 941.400 136.350 942.600 137.100 ;
        RECT 943.950 136.950 946.050 139.050 ;
        RECT 940.800 133.950 942.900 136.050 ;
        RECT 930.900 131.100 939.600 132.300 ;
        RECT 928.800 126.600 930.900 128.700 ;
        RECT 932.100 128.100 934.200 130.200 ;
        RECT 936.000 129.300 938.100 131.100 ;
        RECT 940.950 127.950 943.050 130.050 ;
        RECT 932.400 125.550 933.600 127.800 ;
        RECT 919.950 118.950 922.050 121.050 ;
        RECT 925.950 118.950 928.050 121.050 ;
        RECT 874.950 109.950 877.050 112.050 ;
        RECT 880.950 109.950 883.050 112.050 ;
        RECT 893.700 111.300 895.800 113.400 ;
        RECT 896.700 111.300 898.800 113.400 ;
        RECT 899.700 111.300 901.800 113.400 ;
        RECT 881.400 106.200 882.450 109.950 ;
        RECT 894.300 107.700 895.500 111.300 ;
        RECT 865.950 104.100 868.050 106.200 ;
        RECT 874.950 104.100 877.050 106.200 ;
        RECT 880.950 104.100 883.050 106.200 ;
        RECT 893.400 105.600 895.500 107.700 ;
        RECT 866.400 103.350 867.600 104.100 ;
        RECT 875.400 103.350 876.600 104.100 ;
        RECT 863.100 100.950 865.200 103.050 ;
        RECT 866.100 100.950 868.200 103.050 ;
        RECT 871.800 100.950 873.900 103.050 ;
        RECT 874.800 100.950 876.900 103.050 ;
        RECT 863.400 98.400 864.600 100.650 ;
        RECT 872.400 98.400 873.600 100.650 ;
        RECT 850.950 94.800 853.050 96.900 ;
        RECT 841.950 76.950 844.050 79.050 ;
        RECT 791.700 72.300 793.800 74.400 ;
        RECT 792.300 67.500 793.800 72.300 ;
        RECT 791.700 65.400 793.800 67.500 ;
        RECT 787.950 52.950 790.050 55.050 ;
        RECT 787.950 46.950 790.050 49.050 ;
        RECT 792.300 47.700 793.800 65.400 ;
        RECT 781.950 34.950 784.050 37.050 ;
        RECT 757.950 31.950 760.050 34.050 ;
        RECT 788.400 33.450 789.450 46.950 ;
        RECT 791.700 45.600 793.800 47.700 ;
        RECT 794.700 69.300 796.800 74.400 ;
        RECT 797.700 72.300 799.800 74.400 ;
        RECT 816.600 72.300 818.700 74.400 ;
        RECT 819.600 72.300 822.600 74.400 ;
        RECT 794.700 47.700 795.900 69.300 ;
        RECT 797.700 67.500 799.200 72.300 ;
        RECT 800.100 69.300 802.200 71.400 ;
        RECT 797.100 65.400 799.200 67.500 ;
        RECT 797.700 47.700 799.200 65.400 ;
        RECT 800.700 62.100 801.900 69.300 ;
        RECT 805.500 67.800 807.600 69.900 ;
        RECT 814.200 69.300 816.300 71.400 ;
        RECT 800.100 60.000 802.200 62.100 ;
        RECT 806.700 61.200 807.600 67.800 ;
        RECT 808.950 64.950 811.050 67.050 ;
        RECT 800.700 47.700 801.900 60.000 ;
        RECT 805.500 59.100 807.600 61.200 ;
        RECT 802.800 52.500 804.900 54.600 ;
        RECT 806.700 48.600 807.600 59.100 ;
        RECT 809.400 57.600 810.450 64.950 ;
        RECT 809.400 55.350 810.600 57.600 ;
        RECT 809.100 52.950 811.200 55.050 ;
        RECT 794.700 45.600 796.800 47.700 ;
        RECT 797.700 45.600 799.800 47.700 ;
        RECT 800.700 45.600 802.800 47.700 ;
        RECT 806.100 46.500 808.200 48.600 ;
        RECT 815.100 47.700 816.300 69.300 ;
        RECT 817.500 66.300 818.700 72.300 ;
        RECT 817.500 64.200 819.600 66.300 ;
        RECT 817.500 47.700 818.700 64.200 ;
        RECT 821.100 53.400 822.600 72.300 ;
        RECT 851.400 64.200 852.450 94.800 ;
        RECT 863.400 91.050 864.450 98.400 ;
        RECT 862.950 88.950 865.050 91.050 ;
        RECT 872.400 76.050 873.450 98.400 ;
        RECT 880.800 97.950 882.900 100.050 ;
        RECT 886.800 97.950 888.900 100.050 ;
        RECT 881.400 96.900 882.600 97.650 ;
        RECT 880.950 94.800 883.050 96.900 ;
        RECT 893.400 86.700 894.900 105.600 ;
        RECT 897.300 94.800 898.500 111.300 ;
        RECT 896.400 92.700 898.500 94.800 ;
        RECT 897.300 86.700 898.500 92.700 ;
        RECT 899.700 89.700 900.900 111.300 ;
        RECT 907.800 110.400 909.900 112.500 ;
        RECT 913.200 111.300 915.300 113.400 ;
        RECT 916.200 111.300 918.300 113.400 ;
        RECT 919.200 111.300 921.300 113.400 ;
        RECT 904.800 103.950 906.900 106.050 ;
        RECT 905.400 102.000 906.600 103.650 ;
        RECT 904.950 97.950 907.050 102.000 ;
        RECT 908.400 99.900 909.300 110.400 ;
        RECT 911.100 104.400 913.200 106.500 ;
        RECT 908.400 97.800 910.500 99.900 ;
        RECT 914.100 99.000 915.300 111.300 ;
        RECT 908.400 91.200 909.300 97.800 ;
        RECT 913.800 96.900 915.900 99.000 ;
        RECT 899.700 87.600 901.800 89.700 ;
        RECT 908.400 89.100 910.500 91.200 ;
        RECT 914.100 89.700 915.300 96.900 ;
        RECT 916.800 93.600 918.300 111.300 ;
        RECT 916.800 91.500 918.900 93.600 ;
        RECT 913.800 87.600 915.900 89.700 ;
        RECT 916.800 86.700 918.300 91.500 ;
        RECT 920.100 89.700 921.300 111.300 ;
        RECT 893.400 84.600 896.400 86.700 ;
        RECT 897.300 84.600 899.400 86.700 ;
        RECT 916.200 84.600 918.300 86.700 ;
        RECT 919.200 84.600 921.300 89.700 ;
        RECT 922.200 111.300 924.300 113.400 ;
        RECT 922.200 93.600 923.700 111.300 ;
        RECT 926.400 106.050 927.450 118.950 ;
        RECT 932.400 108.450 933.450 125.550 ;
        RECT 929.400 107.400 933.450 108.450 ;
        RECT 925.950 103.950 928.050 106.050 ;
        RECT 926.400 94.050 927.450 103.950 ;
        RECT 929.400 103.050 930.450 107.400 ;
        RECT 934.950 106.950 937.050 109.050 ;
        RECT 928.950 100.950 931.050 103.050 ;
        RECT 931.950 102.000 934.050 106.050 ;
        RECT 932.400 100.350 933.600 102.000 ;
        RECT 931.800 97.950 933.900 100.050 ;
        RECT 922.200 91.500 924.300 93.600 ;
        RECT 925.950 91.950 928.050 94.050 ;
        RECT 922.200 86.700 923.700 91.500 ;
        RECT 922.200 84.600 924.300 86.700 ;
        RECT 916.950 79.950 919.050 82.050 ;
        RECT 904.950 76.950 907.050 79.050 ;
        RECT 854.400 72.300 857.400 74.400 ;
        RECT 858.300 72.300 860.400 74.400 ;
        RECT 865.950 73.950 868.050 76.050 ;
        RECT 871.950 73.950 874.050 76.050 ;
        RECT 841.950 62.100 844.050 64.200 ;
        RECT 850.950 62.100 853.050 64.200 ;
        RECT 842.400 61.350 843.600 62.100 ;
        RECT 827.100 58.950 829.200 61.050 ;
        RECT 833.100 58.950 835.200 61.050 ;
        RECT 841.800 58.950 843.900 61.050 ;
        RECT 847.800 58.950 849.900 61.050 ;
        RECT 827.400 57.900 828.600 58.650 ;
        RECT 851.400 57.900 852.450 62.100 ;
        RECT 826.950 55.800 829.050 57.900 ;
        RECT 850.950 55.800 853.050 57.900 ;
        RECT 820.500 51.300 822.600 53.400 ;
        RECT 820.500 47.700 821.700 51.300 ;
        RECT 814.200 45.600 816.300 47.700 ;
        RECT 817.200 45.600 819.300 47.700 ;
        RECT 820.200 45.600 822.300 47.700 ;
        RECT 808.950 34.950 811.050 37.050 ;
        RECT 751.950 26.100 754.050 28.200 ;
        RECT 758.400 27.600 759.450 31.950 ;
        RECT 781.500 29.400 783.600 31.500 ;
        RECT 788.400 31.200 789.600 33.450 ;
        RECT 752.400 25.350 753.600 26.100 ;
        RECT 758.400 25.350 759.600 27.600 ;
        RECT 775.950 25.950 778.050 28.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 755.400 20.400 756.600 22.650 ;
        RECT 761.400 21.900 762.600 22.650 ;
        RECT 739.950 16.950 742.050 19.050 ;
        RECT 755.400 7.050 756.450 20.400 ;
        RECT 760.950 19.800 763.050 21.900 ;
        RECT 776.400 21.450 777.450 25.950 ;
        RECT 779.100 22.950 781.200 25.050 ;
        RECT 779.400 21.450 780.600 22.650 ;
        RECT 776.400 20.400 780.600 21.450 ;
        RECT 782.100 16.800 783.000 29.400 ;
        RECT 788.100 28.800 790.200 30.900 ;
        RECT 791.400 29.100 793.500 31.200 ;
        RECT 783.900 27.000 786.000 27.900 ;
        RECT 783.900 25.800 791.100 27.000 ;
        RECT 789.000 24.900 791.100 25.800 ;
        RECT 783.900 24.000 786.000 24.900 ;
        RECT 792.000 24.000 792.900 29.100 ;
        RECT 794.400 27.450 795.600 27.600 ;
        RECT 794.400 26.400 798.450 27.450 ;
        RECT 794.400 25.350 795.600 26.400 ;
        RECT 783.900 23.100 792.900 24.000 ;
        RECT 783.900 22.800 786.000 23.100 ;
        RECT 788.100 19.950 790.200 22.050 ;
        RECT 788.400 17.400 789.600 19.650 ;
        RECT 781.800 14.700 783.900 16.800 ;
        RECT 792.000 16.500 792.900 23.100 ;
        RECT 793.800 22.950 795.900 25.050 ;
        RECT 797.400 24.450 798.450 26.400 ;
        RECT 809.400 24.600 810.450 34.950 ;
        RECT 818.700 33.300 820.800 35.400 ;
        RECT 800.400 24.450 801.600 24.600 ;
        RECT 797.400 24.000 801.600 24.450 ;
        RECT 796.950 23.400 801.600 24.000 ;
        RECT 796.950 19.950 799.050 23.400 ;
        RECT 800.400 22.350 801.600 23.400 ;
        RECT 809.400 22.350 810.600 24.600 ;
        RECT 800.100 19.950 802.200 22.050 ;
        RECT 809.100 19.950 811.200 22.050 ;
        RECT 790.800 14.400 792.900 16.500 ;
        RECT 819.300 15.600 820.800 33.300 ;
        RECT 818.700 13.500 820.800 15.600 ;
        RECT 819.300 8.700 820.800 13.500 ;
        RECT 370.950 4.950 373.050 7.050 ;
        RECT 541.950 4.950 544.050 7.050 ;
        RECT 733.950 4.950 736.050 7.050 ;
        RECT 754.950 4.950 757.050 7.050 ;
        RECT 818.700 6.600 820.800 8.700 ;
        RECT 821.700 33.300 823.800 35.400 ;
        RECT 824.700 33.300 826.800 35.400 ;
        RECT 827.700 33.300 829.800 35.400 ;
        RECT 821.700 11.700 822.900 33.300 ;
        RECT 824.700 15.600 826.200 33.300 ;
        RECT 827.700 21.000 828.900 33.300 ;
        RECT 833.100 32.400 835.200 34.500 ;
        RECT 841.200 33.300 843.300 35.400 ;
        RECT 844.200 33.300 846.300 35.400 ;
        RECT 847.200 33.300 849.300 35.400 ;
        RECT 829.800 26.400 831.900 28.500 ;
        RECT 833.700 21.900 834.600 32.400 ;
        RECT 836.100 25.950 838.200 28.050 ;
        RECT 827.100 18.900 829.200 21.000 ;
        RECT 832.500 19.800 834.600 21.900 ;
        RECT 824.100 13.500 826.200 15.600 ;
        RECT 821.700 6.600 823.800 11.700 ;
        RECT 824.700 8.700 826.200 13.500 ;
        RECT 827.700 11.700 828.900 18.900 ;
        RECT 833.700 13.200 834.600 19.800 ;
        RECT 836.400 23.400 837.600 25.650 ;
        RECT 836.400 16.050 837.450 23.400 ;
        RECT 835.950 13.950 838.050 16.050 ;
        RECT 827.100 9.600 829.200 11.700 ;
        RECT 832.500 11.100 834.600 13.200 ;
        RECT 842.100 11.700 843.300 33.300 ;
        RECT 841.200 9.600 843.300 11.700 ;
        RECT 844.500 16.800 845.700 33.300 ;
        RECT 847.500 29.700 848.700 33.300 ;
        RECT 847.500 27.600 849.600 29.700 ;
        RECT 844.500 14.700 846.600 16.800 ;
        RECT 844.500 8.700 845.700 14.700 ;
        RECT 848.100 8.700 849.600 27.600 ;
        RECT 851.400 19.050 852.450 55.800 ;
        RECT 854.400 53.400 855.900 72.300 ;
        RECT 858.300 66.300 859.500 72.300 ;
        RECT 857.400 64.200 859.500 66.300 ;
        RECT 854.400 51.300 856.500 53.400 ;
        RECT 855.300 47.700 856.500 51.300 ;
        RECT 858.300 47.700 859.500 64.200 ;
        RECT 860.700 69.300 862.800 71.400 ;
        RECT 860.700 47.700 861.900 69.300 ;
        RECT 866.400 57.600 867.450 73.950 ;
        RECT 877.200 72.300 879.300 74.400 ;
        RECT 869.400 67.800 871.500 69.900 ;
        RECT 874.800 69.300 876.900 71.400 ;
        RECT 869.400 61.200 870.300 67.800 ;
        RECT 875.100 62.100 876.300 69.300 ;
        RECT 877.800 67.500 879.300 72.300 ;
        RECT 880.200 69.300 882.300 74.400 ;
        RECT 877.800 65.400 879.900 67.500 ;
        RECT 869.400 59.100 871.500 61.200 ;
        RECT 874.800 60.000 876.900 62.100 ;
        RECT 866.400 55.350 867.600 57.600 ;
        RECT 865.800 52.950 867.900 55.050 ;
        RECT 869.400 48.600 870.300 59.100 ;
        RECT 872.100 52.500 874.200 54.600 ;
        RECT 854.700 45.600 856.800 47.700 ;
        RECT 857.700 45.600 859.800 47.700 ;
        RECT 860.700 45.600 862.800 47.700 ;
        RECT 868.800 46.500 870.900 48.600 ;
        RECT 875.100 47.700 876.300 60.000 ;
        RECT 877.800 47.700 879.300 65.400 ;
        RECT 881.100 47.700 882.300 69.300 ;
        RECT 874.200 45.600 876.300 47.700 ;
        RECT 877.200 45.600 879.300 47.700 ;
        RECT 880.200 45.600 882.300 47.700 ;
        RECT 883.200 72.300 885.300 74.400 ;
        RECT 883.200 67.500 884.700 72.300 ;
        RECT 883.200 65.400 885.300 67.500 ;
        RECT 883.200 47.700 884.700 65.400 ;
        RECT 892.800 58.950 894.900 61.050 ;
        RECT 901.800 58.950 903.900 61.050 ;
        RECT 893.400 56.400 894.600 58.650 ;
        RECT 902.400 57.450 903.600 58.650 ;
        RECT 905.400 57.450 906.450 76.950 ;
        RECT 902.400 56.400 906.450 57.450 ;
        RECT 883.200 45.600 885.300 47.700 ;
        RECT 880.950 37.950 883.050 40.050 ;
        RECT 881.400 27.600 882.450 37.950 ;
        RECT 893.400 37.050 894.450 56.400 ;
        RECT 917.400 55.050 918.450 79.950 ;
        RECT 935.400 73.050 936.450 106.950 ;
        RECT 941.400 102.600 942.450 127.950 ;
        RECT 941.400 100.350 942.600 102.600 ;
        RECT 940.800 97.950 942.900 100.050 ;
        RECT 940.950 91.950 943.050 94.050 ;
        RECT 934.950 70.950 937.050 73.050 ;
        RECT 931.950 64.950 934.050 67.050 ;
        RECT 925.950 60.000 928.050 64.050 ;
        RECT 932.400 60.600 933.450 64.950 ;
        RECT 935.400 64.050 936.450 70.950 ;
        RECT 934.950 61.950 937.050 64.050 ;
        RECT 926.400 58.350 927.600 60.000 ;
        RECT 932.400 58.350 933.600 60.600 ;
        RECT 937.950 58.950 940.050 61.050 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 928.950 55.950 931.050 58.050 ;
        RECT 931.950 55.950 934.050 58.050 ;
        RECT 916.950 52.950 919.050 55.050 ;
        RECT 923.400 54.000 924.600 55.650 ;
        RECT 929.400 54.900 930.600 55.650 ;
        RECT 922.950 49.950 925.050 54.000 ;
        RECT 928.950 52.800 931.050 54.900 ;
        RECT 892.950 34.950 895.050 37.050 ;
        RECT 905.700 33.300 907.800 35.400 ;
        RECT 908.700 33.300 910.800 35.400 ;
        RECT 911.700 33.300 913.800 35.400 ;
        RECT 906.300 29.700 907.500 33.300 ;
        RECT 905.400 27.600 907.500 29.700 ;
        RECT 881.400 25.350 882.600 27.600 ;
        RECT 881.400 22.950 883.500 25.050 ;
        RECT 886.800 22.950 888.900 25.050 ;
        RECT 854.100 19.950 856.200 22.050 ;
        RECT 860.100 19.950 862.200 22.050 ;
        RECT 887.400 21.000 888.600 22.650 ;
        RECT 850.950 16.950 853.050 19.050 ;
        RECT 860.400 18.900 861.600 19.650 ;
        RECT 859.950 16.800 862.050 18.900 ;
        RECT 886.950 16.800 889.050 21.000 ;
        RECT 892.800 19.950 894.900 22.050 ;
        RECT 898.800 19.950 900.900 22.050 ;
        RECT 893.400 18.900 894.600 19.650 ;
        RECT 892.950 16.800 895.050 18.900 ;
        RECT 824.700 6.600 826.800 8.700 ;
        RECT 843.600 6.600 845.700 8.700 ;
        RECT 846.600 6.600 849.600 8.700 ;
        RECT 905.400 8.700 906.900 27.600 ;
        RECT 909.300 16.800 910.500 33.300 ;
        RECT 908.400 14.700 910.500 16.800 ;
        RECT 909.300 8.700 910.500 14.700 ;
        RECT 911.700 11.700 912.900 33.300 ;
        RECT 919.800 32.400 921.900 34.500 ;
        RECT 925.200 33.300 927.300 35.400 ;
        RECT 928.200 33.300 930.300 35.400 ;
        RECT 931.200 33.300 933.300 35.400 ;
        RECT 916.800 25.950 918.900 28.050 ;
        RECT 917.400 24.900 918.600 25.650 ;
        RECT 916.950 22.800 919.050 24.900 ;
        RECT 920.400 21.900 921.300 32.400 ;
        RECT 923.100 26.400 925.200 28.500 ;
        RECT 920.400 19.800 922.500 21.900 ;
        RECT 926.100 21.000 927.300 33.300 ;
        RECT 920.400 13.200 921.300 19.800 ;
        RECT 925.800 18.900 927.900 21.000 ;
        RECT 911.700 9.600 913.800 11.700 ;
        RECT 920.400 11.100 922.500 13.200 ;
        RECT 926.100 11.700 927.300 18.900 ;
        RECT 928.800 15.600 930.300 33.300 ;
        RECT 928.800 13.500 930.900 15.600 ;
        RECT 925.800 9.600 927.900 11.700 ;
        RECT 928.800 8.700 930.300 13.500 ;
        RECT 932.100 11.700 933.300 33.300 ;
        RECT 905.400 6.600 908.400 8.700 ;
        RECT 909.300 6.600 911.400 8.700 ;
        RECT 928.200 6.600 930.300 8.700 ;
        RECT 931.200 6.600 933.300 11.700 ;
        RECT 934.200 33.300 936.300 35.400 ;
        RECT 934.200 15.600 935.700 33.300 ;
        RECT 938.400 19.050 939.450 58.950 ;
        RECT 941.400 36.450 942.450 91.950 ;
        RECT 944.400 79.050 945.450 136.950 ;
        RECT 946.950 133.950 949.050 136.050 ;
        RECT 947.400 91.050 948.450 133.950 ;
        RECT 946.950 88.950 949.050 91.050 ;
        RECT 943.950 76.950 946.050 79.050 ;
        RECT 943.950 61.950 946.050 64.050 ;
        RECT 944.400 52.050 945.450 61.950 ;
        RECT 947.400 61.200 948.450 88.950 ;
        RECT 950.400 76.050 951.450 148.950 ;
        RECT 952.950 142.950 955.050 145.050 ;
        RECT 953.400 132.900 954.450 142.950 ;
        RECT 956.400 139.050 957.450 203.400 ;
        RECT 958.950 202.950 961.050 203.400 ;
        RECT 958.950 187.950 961.050 190.050 ;
        RECT 959.400 148.050 960.450 187.950 ;
        RECT 962.400 151.050 963.450 214.950 ;
        RECT 965.400 210.900 966.450 217.950 ;
        RECT 974.400 216.600 975.450 220.950 ;
        RECT 977.400 217.050 978.450 268.950 ;
        RECT 979.950 261.450 982.050 265.050 ;
        RECT 983.400 261.450 984.600 261.600 ;
        RECT 979.950 261.000 984.600 261.450 ;
        RECT 980.400 260.400 984.600 261.000 ;
        RECT 983.400 259.350 984.600 260.400 ;
        RECT 982.950 256.950 985.050 259.050 ;
        RECT 985.950 256.950 988.050 259.050 ;
        RECT 986.400 255.000 987.600 256.650 ;
        RECT 985.950 250.950 988.050 255.000 ;
        RECT 992.400 247.050 993.450 301.800 ;
        RECT 997.950 294.600 1002.000 295.050 ;
        RECT 1010.400 294.600 1011.450 304.950 ;
        RECT 1015.950 298.950 1018.050 301.050 ;
        RECT 997.950 292.950 1002.600 294.600 ;
        RECT 998.400 286.050 999.450 292.950 ;
        RECT 1001.400 292.350 1002.600 292.950 ;
        RECT 1010.400 294.450 1011.600 294.600 ;
        RECT 1010.400 293.400 1014.450 294.450 ;
        RECT 1010.400 292.350 1011.600 293.400 ;
        RECT 1001.100 289.950 1003.200 292.050 ;
        RECT 1006.500 289.950 1008.600 292.050 ;
        RECT 1009.800 289.950 1011.900 292.050 ;
        RECT 1007.400 288.900 1008.600 289.650 ;
        RECT 1006.950 286.800 1009.050 288.900 ;
        RECT 997.950 283.950 1000.050 286.050 ;
        RECT 994.950 274.950 997.050 277.050 ;
        RECT 995.400 253.050 996.450 274.950 ;
        RECT 997.950 265.950 1000.050 268.050 ;
        RECT 998.400 255.900 999.450 265.950 ;
        RECT 1013.400 265.200 1014.450 293.400 ;
        RECT 1012.950 263.100 1015.050 265.200 ;
        RECT 1016.400 265.050 1017.450 298.950 ;
        RECT 1015.950 262.950 1018.050 265.050 ;
        RECT 1000.950 259.950 1003.050 262.050 ;
        RECT 1006.950 260.100 1009.050 262.200 ;
        RECT 1007.400 259.350 1008.600 260.100 ;
        RECT 1012.950 259.950 1015.050 262.050 ;
        RECT 1013.400 259.350 1014.600 259.950 ;
        RECT 1003.950 256.950 1006.050 259.050 ;
        RECT 1006.950 256.950 1009.050 259.050 ;
        RECT 1009.950 256.950 1012.050 259.050 ;
        RECT 1012.950 256.950 1015.050 259.050 ;
        RECT 997.950 253.800 1000.050 255.900 ;
        RECT 1000.950 253.950 1003.050 256.050 ;
        RECT 1004.400 255.900 1005.600 256.650 ;
        RECT 1010.400 255.900 1011.600 256.650 ;
        RECT 1019.400 255.900 1020.450 352.950 ;
        RECT 1024.950 334.950 1027.050 337.050 ;
        RECT 1027.950 334.950 1030.050 337.050 ;
        RECT 1028.400 333.900 1029.600 334.650 ;
        RECT 1034.400 334.050 1035.450 364.800 ;
        RECT 1037.400 346.050 1038.450 382.950 ;
        RECT 1039.950 367.950 1042.050 370.050 ;
        RECT 1036.950 343.950 1039.050 346.050 ;
        RECT 1040.400 336.450 1041.450 367.950 ;
        RECT 1037.400 335.400 1041.450 336.450 ;
        RECT 1027.950 331.800 1030.050 333.900 ;
        RECT 1033.950 331.950 1036.050 334.050 ;
        RECT 1037.400 319.050 1038.450 335.400 ;
        RECT 1039.950 331.950 1042.050 334.050 ;
        RECT 1036.950 316.950 1039.050 319.050 ;
        RECT 1027.950 304.950 1030.050 307.050 ;
        RECT 1021.950 293.100 1024.050 295.200 ;
        RECT 1028.400 294.600 1029.450 304.950 ;
        RECT 1022.400 288.450 1023.450 293.100 ;
        RECT 1028.400 292.350 1029.600 294.600 ;
        RECT 1033.950 293.100 1036.050 295.200 ;
        RECT 1034.400 292.350 1035.600 293.100 ;
        RECT 1027.950 289.950 1030.050 292.050 ;
        RECT 1030.950 289.950 1033.050 292.050 ;
        RECT 1033.950 289.950 1036.050 292.050 ;
        RECT 1024.950 288.450 1027.050 288.900 ;
        RECT 1022.400 287.400 1027.050 288.450 ;
        RECT 1024.950 286.800 1027.050 287.400 ;
        RECT 1031.400 287.400 1032.600 289.650 ;
        RECT 1021.950 262.950 1024.050 265.050 ;
        RECT 994.950 250.950 997.050 253.050 ;
        RECT 979.950 244.950 982.050 247.050 ;
        RECT 991.950 244.950 994.050 247.050 ;
        RECT 974.400 214.350 975.600 216.600 ;
        RECT 976.950 214.950 979.050 217.050 ;
        RECT 970.950 211.950 973.050 214.050 ;
        RECT 973.950 211.950 976.050 214.050 ;
        RECT 971.400 210.900 972.600 211.650 ;
        RECT 964.950 208.800 967.050 210.900 ;
        RECT 970.950 208.800 973.050 210.900 ;
        RECT 967.950 187.950 970.050 190.050 ;
        RECT 968.400 183.600 969.450 187.950 ;
        RECT 968.400 181.350 969.600 183.600 ;
        RECT 973.950 182.100 976.050 184.200 ;
        RECT 974.400 181.350 975.600 182.100 ;
        RECT 967.950 178.950 970.050 181.050 ;
        RECT 970.950 178.950 973.050 181.050 ;
        RECT 973.950 178.950 976.050 181.050 ;
        RECT 971.400 177.900 972.600 178.650 ;
        RECT 970.950 175.800 973.050 177.900 ;
        RECT 980.400 169.050 981.450 244.950 ;
        RECT 998.400 238.050 999.450 253.800 ;
        RECT 985.950 235.950 988.050 238.050 ;
        RECT 997.950 235.950 1000.050 238.050 ;
        RECT 982.950 214.950 985.050 217.050 ;
        RECT 983.400 190.050 984.450 214.950 ;
        RECT 986.400 210.900 987.450 235.950 ;
        RECT 1001.400 217.200 1002.450 253.950 ;
        RECT 1003.950 253.800 1006.050 255.900 ;
        RECT 1009.950 253.800 1012.050 255.900 ;
        RECT 1018.950 253.800 1021.050 255.900 ;
        RECT 1022.400 241.050 1023.450 262.950 ;
        RECT 1025.400 262.050 1026.450 286.800 ;
        RECT 1031.400 283.050 1032.450 287.400 ;
        RECT 1030.950 280.950 1033.050 283.050 ;
        RECT 1024.950 259.950 1027.050 262.050 ;
        RECT 1033.950 261.000 1036.050 265.050 ;
        RECT 1040.400 262.200 1041.450 331.950 ;
        RECT 1025.400 253.050 1026.450 259.950 ;
        RECT 1034.400 259.350 1035.600 261.000 ;
        RECT 1039.800 260.100 1041.900 262.200 ;
        RECT 1043.400 262.050 1044.450 397.950 ;
        RECT 1040.400 259.350 1041.600 260.100 ;
        RECT 1042.950 259.950 1045.050 262.050 ;
        RECT 1030.950 256.950 1033.050 259.050 ;
        RECT 1033.950 256.950 1036.050 259.050 ;
        RECT 1036.950 256.950 1039.050 259.050 ;
        RECT 1039.950 256.950 1042.050 259.050 ;
        RECT 1031.400 256.050 1032.600 256.650 ;
        RECT 1027.950 254.400 1032.600 256.050 ;
        RECT 1037.400 255.900 1038.600 256.650 ;
        RECT 1027.950 253.950 1032.000 254.400 ;
        RECT 1024.950 250.950 1027.050 253.050 ;
        RECT 1003.950 238.950 1006.050 241.050 ;
        RECT 1021.950 238.950 1024.050 241.050 ;
        RECT 994.950 215.100 997.050 217.200 ;
        RECT 1000.950 215.100 1003.050 217.200 ;
        RECT 995.400 214.350 996.600 215.100 ;
        RECT 991.950 211.950 994.050 214.050 ;
        RECT 994.950 211.950 997.050 214.050 ;
        RECT 997.950 211.950 1000.050 214.050 ;
        RECT 985.950 208.800 988.050 210.900 ;
        RECT 992.400 209.400 993.600 211.650 ;
        RECT 998.400 210.900 999.600 211.650 ;
        RECT 982.950 187.950 985.050 190.050 ;
        RECT 982.950 182.100 985.050 184.200 ;
        RECT 983.400 178.050 984.450 182.100 ;
        RECT 982.950 175.950 985.050 178.050 ;
        RECT 979.950 166.950 982.050 169.050 ;
        RECT 976.950 157.950 979.050 160.050 ;
        RECT 961.950 148.950 964.050 151.050 ;
        RECT 958.950 145.950 961.050 148.050 ;
        RECT 955.950 136.950 958.050 139.050 ;
        RECT 962.400 138.600 963.450 148.950 ;
        RECT 967.950 142.950 970.050 145.050 ;
        RECT 962.400 136.350 963.600 138.600 ;
        RECT 958.950 133.950 961.050 136.050 ;
        RECT 961.950 133.950 964.050 136.050 ;
        RECT 959.400 132.900 960.600 133.650 ;
        RECT 952.950 130.800 955.050 132.900 ;
        RECT 958.950 130.800 961.050 132.900 ;
        RECT 949.950 73.950 952.050 76.050 ;
        RECT 949.950 64.950 952.050 67.050 ;
        RECT 946.950 59.100 949.050 61.200 ;
        RECT 950.400 60.600 951.450 64.950 ;
        RECT 953.400 64.050 954.450 130.800 ;
        RECT 964.500 107.400 966.600 109.500 ;
        RECT 968.400 109.050 969.450 142.950 ;
        RECT 977.400 132.450 978.450 157.950 ;
        RECT 986.400 145.050 987.450 208.800 ;
        RECT 992.400 199.050 993.450 209.400 ;
        RECT 997.950 208.800 1000.050 210.900 ;
        RECT 997.950 199.950 1000.050 202.050 ;
        RECT 991.950 196.950 994.050 199.050 ;
        RECT 998.400 187.050 999.450 199.950 ;
        RECT 1000.950 187.950 1003.050 190.050 ;
        RECT 994.950 183.000 997.050 187.050 ;
        RECT 997.950 184.950 1000.050 187.050 ;
        RECT 995.400 181.350 996.600 183.000 ;
        RECT 1001.400 181.050 1002.450 187.950 ;
        RECT 1004.400 187.050 1005.450 238.950 ;
        RECT 1006.950 232.950 1009.050 235.050 ;
        RECT 1007.400 211.050 1008.450 232.950 ;
        RECT 1015.950 220.950 1018.050 223.050 ;
        RECT 1016.400 216.600 1017.450 220.950 ;
        RECT 1016.400 214.350 1017.600 216.600 ;
        RECT 1021.950 215.100 1024.050 217.200 ;
        RECT 1022.400 214.350 1023.600 215.100 ;
        RECT 1015.950 211.950 1018.050 214.050 ;
        RECT 1018.950 211.950 1021.050 214.050 ;
        RECT 1021.950 211.950 1024.050 214.050 ;
        RECT 1006.950 208.950 1009.050 211.050 ;
        RECT 1019.400 210.900 1020.600 211.650 ;
        RECT 1018.950 208.800 1021.050 210.900 ;
        RECT 1028.400 199.050 1029.450 253.950 ;
        RECT 1036.950 253.800 1039.050 255.900 ;
        RECT 1042.950 253.950 1045.050 256.050 ;
        RECT 1030.950 250.950 1033.050 253.050 ;
        RECT 1027.950 196.950 1030.050 199.050 ;
        RECT 1031.400 195.450 1032.450 250.950 ;
        RECT 1033.950 235.950 1036.050 238.050 ;
        RECT 1028.400 194.400 1032.450 195.450 ;
        RECT 1003.950 184.950 1006.050 187.050 ;
        RECT 991.950 178.950 994.050 181.050 ;
        RECT 994.950 178.950 997.050 181.050 ;
        RECT 1000.950 178.950 1003.050 181.050 ;
        RECT 992.400 177.900 993.600 178.650 ;
        RECT 1004.400 177.900 1005.450 184.950 ;
        RECT 1006.950 182.100 1009.050 184.200 ;
        RECT 1015.950 182.100 1018.050 184.200 ;
        RECT 1021.950 182.100 1024.050 184.200 ;
        RECT 991.950 175.800 994.050 177.900 ;
        RECT 1003.950 175.800 1006.050 177.900 ;
        RECT 1007.400 172.050 1008.450 182.100 ;
        RECT 1016.400 181.350 1017.600 182.100 ;
        RECT 1022.400 181.350 1023.600 182.100 ;
        RECT 1012.950 178.950 1015.050 181.050 ;
        RECT 1015.950 178.950 1018.050 181.050 ;
        RECT 1018.950 178.950 1021.050 181.050 ;
        RECT 1021.950 178.950 1024.050 181.050 ;
        RECT 1013.400 177.900 1014.600 178.650 ;
        RECT 1019.400 177.900 1020.600 178.650 ;
        RECT 1012.950 175.800 1015.050 177.900 ;
        RECT 1018.950 175.800 1021.050 177.900 ;
        RECT 1028.400 177.450 1029.450 194.400 ;
        RECT 1030.950 181.950 1033.050 184.050 ;
        RECT 1025.400 176.400 1029.450 177.450 ;
        RECT 1006.950 169.950 1009.050 172.050 ;
        RECT 1000.950 166.950 1003.050 169.050 ;
        RECT 982.800 142.500 984.900 144.600 ;
        RECT 985.950 142.950 988.050 145.050 ;
        RECT 980.100 133.950 982.200 136.050 ;
        RECT 983.100 135.300 984.300 142.500 ;
        RECT 986.400 139.350 987.600 141.600 ;
        RECT 992.400 141.300 994.500 143.400 ;
        RECT 986.100 136.950 988.200 139.050 ;
        RECT 989.100 137.700 991.200 139.800 ;
        RECT 989.100 135.300 990.000 137.700 ;
        RECT 983.100 134.100 990.000 135.300 ;
        RECT 980.400 132.450 981.600 133.650 ;
        RECT 977.400 131.400 981.600 132.450 ;
        RECT 983.100 128.700 984.000 134.100 ;
        RECT 984.900 132.300 987.000 133.200 ;
        RECT 992.700 132.300 993.600 141.300 ;
        RECT 997.950 139.950 1000.050 142.050 ;
        RECT 994.950 137.100 997.050 139.200 ;
        RECT 995.400 136.350 996.600 137.100 ;
        RECT 994.800 133.950 996.900 136.050 ;
        RECT 984.900 131.100 993.600 132.300 ;
        RECT 982.800 126.600 984.900 128.700 ;
        RECT 986.100 128.100 988.200 130.200 ;
        RECT 990.000 129.300 992.100 131.100 ;
        RECT 986.400 125.550 987.600 127.800 ;
        RECT 970.950 109.950 973.050 112.050 ;
        RECT 971.400 109.200 972.600 109.950 ;
        RECT 962.100 100.950 964.200 103.050 ;
        RECT 962.400 99.450 963.600 100.650 ;
        RECT 959.400 98.400 963.600 99.450 ;
        RECT 959.400 82.050 960.450 98.400 ;
        RECT 965.100 94.800 966.000 107.400 ;
        RECT 967.950 106.950 970.050 109.050 ;
        RECT 971.100 106.800 973.200 108.900 ;
        RECT 974.400 107.100 976.500 109.200 ;
        RECT 966.900 105.000 969.000 105.900 ;
        RECT 966.900 103.800 974.100 105.000 ;
        RECT 972.000 102.900 974.100 103.800 ;
        RECT 966.900 102.000 969.000 102.900 ;
        RECT 975.000 102.000 975.900 107.100 ;
        RECT 986.400 106.200 987.450 125.550 ;
        RECT 976.950 104.100 979.050 106.200 ;
        RECT 985.950 104.100 988.050 106.200 ;
        RECT 998.400 105.600 999.450 139.950 ;
        RECT 1001.400 133.050 1002.450 166.950 ;
        RECT 1025.400 166.050 1026.450 176.400 ;
        RECT 1006.950 163.950 1009.050 166.050 ;
        RECT 1024.950 163.950 1027.050 166.050 ;
        RECT 1000.950 130.950 1003.050 133.050 ;
        RECT 977.400 103.350 978.600 104.100 ;
        RECT 966.900 101.100 975.900 102.000 ;
        RECT 966.900 100.800 969.000 101.100 ;
        RECT 971.100 97.950 973.200 100.050 ;
        RECT 971.400 95.400 972.600 97.650 ;
        RECT 964.800 92.700 966.900 94.800 ;
        RECT 975.000 94.500 975.900 101.100 ;
        RECT 976.800 100.950 978.900 103.050 ;
        RECT 986.400 97.050 987.450 104.100 ;
        RECT 998.400 103.350 999.600 105.600 ;
        RECT 994.950 100.950 997.050 103.050 ;
        RECT 997.950 100.950 1000.050 103.050 ;
        RECT 1000.950 100.950 1003.050 103.050 ;
        RECT 995.400 98.400 996.600 100.650 ;
        RECT 1001.400 99.000 1002.600 100.650 ;
        RECT 985.950 94.950 988.050 97.050 ;
        RECT 973.800 92.400 975.900 94.500 ;
        RECT 958.950 79.950 961.050 82.050 ;
        RECT 985.950 79.950 988.050 82.050 ;
        RECT 970.950 73.950 973.050 76.050 ;
        RECT 952.950 61.950 955.050 64.050 ;
        RECT 950.400 58.350 951.600 60.600 ;
        RECT 955.950 59.100 958.050 61.200 ;
        RECT 956.400 58.350 957.600 59.100 ;
        RECT 964.950 58.950 967.050 61.050 ;
        RECT 949.950 55.950 952.050 58.050 ;
        RECT 952.950 55.950 955.050 58.050 ;
        RECT 955.950 55.950 958.050 58.050 ;
        RECT 958.950 55.950 961.050 58.050 ;
        RECT 953.400 53.400 954.600 55.650 ;
        RECT 959.400 53.400 960.600 55.650 ;
        RECT 943.950 49.950 946.050 52.050 ;
        RECT 953.400 46.050 954.450 53.400 ;
        RECT 955.950 49.950 958.050 52.050 ;
        RECT 952.950 43.950 955.050 46.050 ;
        RECT 956.400 40.050 957.450 49.950 ;
        RECT 955.950 37.950 958.050 40.050 ;
        RECT 943.950 36.450 946.050 37.050 ;
        RECT 941.400 35.400 946.050 36.450 ;
        RECT 943.950 34.950 946.050 35.400 ;
        RECT 944.400 24.600 945.450 34.950 ;
        RECT 952.950 31.950 955.050 34.050 ;
        RECT 953.400 24.600 954.450 31.950 ;
        RECT 959.400 25.050 960.450 53.400 ;
        RECT 965.400 46.050 966.450 58.950 ;
        RECT 964.950 43.950 967.050 46.050 ;
        RECT 971.400 34.050 972.450 73.950 ;
        RECT 973.950 64.950 976.050 67.050 ;
        RECT 974.400 55.050 975.450 64.950 ;
        RECT 976.950 59.100 979.050 61.200 ;
        RECT 986.400 60.600 987.450 79.950 ;
        RECT 995.400 61.200 996.450 98.400 ;
        RECT 1000.950 94.950 1003.050 99.000 ;
        RECT 1007.400 94.050 1008.450 163.950 ;
        RECT 1027.950 160.950 1030.050 163.050 ;
        RECT 1012.950 145.950 1015.050 148.050 ;
        RECT 1013.400 138.600 1014.450 145.950 ;
        RECT 1013.400 136.350 1014.600 138.600 ;
        RECT 1018.950 138.000 1021.050 142.050 ;
        RECT 1019.400 136.350 1020.600 138.000 ;
        RECT 1012.950 133.950 1015.050 136.050 ;
        RECT 1015.950 133.950 1018.050 136.050 ;
        RECT 1018.950 133.950 1021.050 136.050 ;
        RECT 1021.950 133.950 1024.050 136.050 ;
        RECT 1016.400 132.900 1017.600 133.650 ;
        RECT 1015.950 130.800 1018.050 132.900 ;
        RECT 1022.400 131.400 1023.600 133.650 ;
        RECT 1022.400 127.050 1023.450 131.400 ;
        RECT 1021.950 124.950 1024.050 127.050 ;
        RECT 1022.400 105.600 1023.450 124.950 ;
        RECT 1022.400 103.350 1023.600 105.600 ;
        RECT 1018.950 100.950 1021.050 103.050 ;
        RECT 1021.950 100.950 1024.050 103.050 ;
        RECT 1019.400 98.400 1020.600 100.650 ;
        RECT 1006.950 91.950 1009.050 94.050 ;
        RECT 1019.400 82.050 1020.450 98.400 ;
        RECT 1021.950 91.950 1024.050 94.050 ;
        RECT 1003.950 79.950 1006.050 82.050 ;
        RECT 1018.950 79.950 1021.050 82.050 ;
        RECT 977.400 58.350 978.600 59.100 ;
        RECT 986.400 58.350 987.600 60.600 ;
        RECT 994.950 59.100 997.050 61.200 ;
        RECT 1004.400 60.600 1005.450 79.950 ;
        RECT 1018.950 70.950 1021.050 73.050 ;
        RECT 1015.950 64.950 1018.050 67.050 ;
        RECT 977.100 55.950 979.200 58.050 ;
        RECT 982.500 55.950 984.600 58.050 ;
        RECT 985.800 55.950 987.900 58.050 ;
        RECT 973.950 52.950 976.050 55.050 ;
        RECT 983.400 53.400 984.600 55.650 ;
        RECT 983.400 49.050 984.450 53.400 ;
        RECT 995.400 49.050 996.450 59.100 ;
        RECT 1004.400 58.350 1005.600 60.600 ;
        RECT 1009.950 59.100 1012.050 61.200 ;
        RECT 1010.400 58.350 1011.600 59.100 ;
        RECT 1003.950 55.950 1006.050 58.050 ;
        RECT 1006.950 55.950 1009.050 58.050 ;
        RECT 1009.950 55.950 1012.050 58.050 ;
        RECT 1007.400 54.900 1008.600 55.650 ;
        RECT 1006.950 52.800 1009.050 54.900 ;
        RECT 982.950 46.950 985.050 49.050 ;
        RECT 994.950 46.950 997.050 49.050 ;
        RECT 1006.950 46.950 1009.050 49.050 ;
        RECT 982.950 37.950 985.050 40.050 ;
        RECT 970.950 31.950 973.050 34.050 ;
        RECT 983.400 28.200 984.450 37.950 ;
        RECT 1007.400 33.450 1008.450 46.950 ;
        RECT 1003.800 30.300 1005.900 32.400 ;
        RECT 1007.400 31.200 1008.600 33.450 ;
        RECT 1016.400 31.050 1017.450 64.950 ;
        RECT 961.950 25.950 964.050 28.050 ;
        RECT 976.950 26.100 979.050 28.200 ;
        RECT 982.950 26.100 985.050 28.200 ;
        RECT 1000.950 26.100 1003.050 28.200 ;
        RECT 944.400 22.350 945.600 24.600 ;
        RECT 953.400 22.350 954.600 24.600 ;
        RECT 958.950 22.950 961.050 25.050 ;
        RECT 962.400 22.050 963.450 25.950 ;
        RECT 977.400 25.350 978.600 26.100 ;
        RECT 983.400 25.350 984.600 26.100 ;
        RECT 1001.400 25.350 1002.600 26.100 ;
        RECT 973.950 22.950 976.050 25.050 ;
        RECT 976.950 22.950 979.050 25.050 ;
        RECT 979.950 22.950 982.050 25.050 ;
        RECT 982.950 22.950 985.050 25.050 ;
        RECT 1001.100 22.950 1003.200 25.050 ;
        RECT 1004.100 24.900 1005.000 30.300 ;
        RECT 1007.100 28.800 1009.200 30.900 ;
        RECT 1011.000 27.900 1013.100 29.700 ;
        RECT 1015.950 28.950 1018.050 31.050 ;
        RECT 1005.900 26.700 1014.600 27.900 ;
        RECT 1005.900 25.800 1008.000 26.700 ;
        RECT 1004.100 23.700 1011.000 24.900 ;
        RECT 943.800 19.950 945.900 22.050 ;
        RECT 952.800 19.950 954.900 22.050 ;
        RECT 961.950 19.950 964.050 22.050 ;
        RECT 974.400 21.900 975.600 22.650 ;
        RECT 973.950 19.800 976.050 21.900 ;
        RECT 980.400 21.000 981.600 22.650 ;
        RECT 937.950 16.950 940.050 19.050 ;
        RECT 979.950 16.950 982.050 21.000 ;
        RECT 1004.100 16.500 1005.300 23.700 ;
        RECT 1007.100 19.950 1009.200 22.050 ;
        RECT 1010.100 21.300 1011.000 23.700 ;
        RECT 1007.400 17.400 1008.600 19.650 ;
        RECT 1010.100 19.200 1012.200 21.300 ;
        RECT 1013.700 17.700 1014.600 26.700 ;
        RECT 1015.800 22.950 1017.900 25.050 ;
        RECT 1016.400 21.450 1017.600 22.650 ;
        RECT 1019.400 21.450 1020.450 70.950 ;
        RECT 1022.400 43.050 1023.450 91.950 ;
        RECT 1028.400 60.600 1029.450 160.950 ;
        RECT 1031.400 127.050 1032.450 181.950 ;
        RECT 1030.950 124.950 1033.050 127.050 ;
        RECT 1034.400 67.050 1035.450 235.950 ;
        RECT 1033.950 64.950 1036.050 67.050 ;
        RECT 1037.400 63.450 1038.450 253.800 ;
        RECT 1039.950 250.950 1042.050 253.050 ;
        RECT 1040.400 202.050 1041.450 250.950 ;
        RECT 1039.950 199.950 1042.050 202.050 ;
        RECT 1034.400 62.400 1038.450 63.450 ;
        RECT 1034.400 60.600 1035.450 62.400 ;
        RECT 1028.400 58.350 1029.600 60.600 ;
        RECT 1034.400 58.350 1035.600 60.600 ;
        RECT 1027.950 55.950 1030.050 58.050 ;
        RECT 1030.950 55.950 1033.050 58.050 ;
        RECT 1033.950 55.950 1036.050 58.050 ;
        RECT 1036.950 55.950 1039.050 58.050 ;
        RECT 1031.400 53.400 1032.600 55.650 ;
        RECT 1037.400 53.400 1038.600 55.650 ;
        RECT 1021.950 40.950 1024.050 43.050 ;
        RECT 1024.950 28.950 1027.050 31.050 ;
        RECT 1016.400 20.400 1020.450 21.450 ;
        RECT 1025.400 19.050 1026.450 28.950 ;
        RECT 1031.400 27.450 1032.450 53.400 ;
        RECT 1037.400 49.050 1038.450 53.400 ;
        RECT 1043.400 49.050 1044.450 253.950 ;
        RECT 1036.950 46.950 1039.050 49.050 ;
        RECT 1042.950 46.950 1045.050 49.050 ;
        RECT 1036.950 40.950 1039.050 43.050 ;
        RECT 1028.400 26.400 1032.450 27.450 ;
        RECT 1037.400 27.600 1038.450 40.950 ;
        RECT 1028.400 21.900 1029.450 26.400 ;
        RECT 1037.400 25.350 1038.600 27.600 ;
        RECT 1033.950 22.950 1036.050 25.050 ;
        RECT 1036.950 22.950 1039.050 25.050 ;
        RECT 1039.950 22.950 1042.050 25.050 ;
        RECT 1027.950 19.800 1030.050 21.900 ;
        RECT 1034.400 21.000 1035.600 22.650 ;
        RECT 1040.400 21.900 1041.600 22.650 ;
        RECT 934.200 13.500 936.300 15.600 ;
        RECT 1003.800 14.400 1005.900 16.500 ;
        RECT 1013.400 15.600 1015.500 17.700 ;
        RECT 1024.950 16.950 1027.050 19.050 ;
        RECT 1033.950 16.950 1036.050 21.000 ;
        RECT 1039.950 19.800 1042.050 21.900 ;
        RECT 934.200 8.700 935.700 13.500 ;
        RECT 934.200 6.600 936.300 8.700 ;
      LAYER metal3 ;
        RECT 406.950 969.600 409.050 970.050 ;
        RECT 445.950 969.600 448.050 970.050 ;
        RECT 406.950 968.400 448.050 969.600 ;
        RECT 406.950 967.950 409.050 968.400 ;
        RECT 445.950 967.950 448.050 968.400 ;
        RECT 451.950 969.600 454.050 970.050 ;
        RECT 472.950 969.600 475.050 970.050 ;
        RECT 451.950 968.400 475.050 969.600 ;
        RECT 451.950 967.950 454.050 968.400 ;
        RECT 472.950 967.950 475.050 968.400 ;
        RECT 490.950 969.600 493.050 970.050 ;
        RECT 619.950 969.600 622.050 970.050 ;
        RECT 631.950 969.600 634.050 970.050 ;
        RECT 490.950 968.400 634.050 969.600 ;
        RECT 490.950 967.950 493.050 968.400 ;
        RECT 619.950 967.950 622.050 968.400 ;
        RECT 631.950 967.950 634.050 968.400 ;
        RECT 664.950 969.600 667.050 970.050 ;
        RECT 736.950 969.600 739.050 970.050 ;
        RECT 664.950 968.400 739.050 969.600 ;
        RECT 664.950 967.950 667.050 968.400 ;
        RECT 736.950 967.950 739.050 968.400 ;
        RECT 742.950 969.600 745.050 970.050 ;
        RECT 766.950 969.600 769.050 970.050 ;
        RECT 742.950 968.400 769.050 969.600 ;
        RECT 742.950 967.950 745.050 968.400 ;
        RECT 766.950 967.950 769.050 968.400 ;
        RECT 949.950 969.600 952.050 970.050 ;
        RECT 967.950 969.600 970.050 970.050 ;
        RECT 949.950 968.400 970.050 969.600 ;
        RECT 949.950 967.950 952.050 968.400 ;
        RECT 967.950 967.950 970.050 968.400 ;
        RECT 358.950 966.600 361.050 967.050 ;
        RECT 373.950 966.600 376.050 967.050 ;
        RECT 358.950 965.400 376.050 966.600 ;
        RECT 358.950 964.950 361.050 965.400 ;
        RECT 373.950 964.950 376.050 965.400 ;
        RECT 448.950 966.600 451.050 967.050 ;
        RECT 520.950 966.600 523.050 967.050 ;
        RECT 448.950 965.400 523.050 966.600 ;
        RECT 448.950 964.950 451.050 965.400 ;
        RECT 520.950 964.950 523.050 965.400 ;
        RECT 592.950 966.600 595.050 967.050 ;
        RECT 598.950 966.600 601.050 967.050 ;
        RECT 592.950 965.400 601.050 966.600 ;
        RECT 592.950 964.950 595.050 965.400 ;
        RECT 598.950 964.950 601.050 965.400 ;
        RECT 835.950 966.600 838.050 967.050 ;
        RECT 898.950 966.600 901.050 967.050 ;
        RECT 970.950 966.600 973.050 967.050 ;
        RECT 835.950 965.400 973.050 966.600 ;
        RECT 835.950 964.950 838.050 965.400 ;
        RECT 898.950 964.950 901.050 965.400 ;
        RECT 970.950 964.950 973.050 965.400 ;
        RECT 979.950 966.600 982.050 967.050 ;
        RECT 1030.950 966.600 1033.050 967.050 ;
        RECT 979.950 965.400 1033.050 966.600 ;
        RECT 979.950 964.950 982.050 965.400 ;
        RECT 1030.950 964.950 1033.050 965.400 ;
        RECT 22.950 963.600 25.050 964.200 ;
        RECT 40.950 963.750 43.050 964.200 ;
        RECT 61.950 963.750 64.050 964.200 ;
        RECT 40.950 963.600 64.050 963.750 ;
        RECT 22.950 962.550 64.050 963.600 ;
        RECT 22.950 962.400 43.050 962.550 ;
        RECT 22.950 962.100 25.050 962.400 ;
        RECT 40.950 962.100 43.050 962.400 ;
        RECT 61.950 962.100 64.050 962.550 ;
        RECT 121.950 963.600 124.050 964.050 ;
        RECT 136.950 963.600 139.050 964.050 ;
        RECT 121.950 962.400 139.050 963.600 ;
        RECT 121.950 961.950 124.050 962.400 ;
        RECT 136.950 961.950 139.050 962.400 ;
        RECT 205.950 963.600 208.050 964.050 ;
        RECT 259.950 963.600 262.050 964.050 ;
        RECT 367.950 963.600 370.050 964.200 ;
        RECT 205.950 962.400 262.050 963.600 ;
        RECT 305.400 963.000 370.050 963.600 ;
        RECT 205.950 961.950 208.050 962.400 ;
        RECT 259.950 961.950 262.050 962.400 ;
        RECT 304.950 962.400 370.050 963.000 ;
        RECT 199.950 960.750 202.050 961.200 ;
        RECT 265.950 960.750 268.050 961.200 ;
        RECT 199.950 959.550 268.050 960.750 ;
        RECT 199.950 959.100 202.050 959.550 ;
        RECT 265.950 959.100 268.050 959.550 ;
        RECT 304.950 958.950 307.050 962.400 ;
        RECT 367.950 962.100 370.050 962.400 ;
        RECT 379.950 963.600 382.050 964.050 ;
        RECT 391.950 963.600 394.050 964.200 ;
        RECT 379.950 962.400 394.050 963.600 ;
        RECT 379.950 961.950 382.050 962.400 ;
        RECT 391.950 962.100 394.050 962.400 ;
        RECT 397.950 963.600 400.050 964.200 ;
        RECT 421.950 963.600 424.050 964.200 ;
        RECT 397.950 962.400 424.050 963.600 ;
        RECT 397.950 962.100 400.050 962.400 ;
        RECT 421.950 962.100 424.050 962.400 ;
        RECT 430.950 963.600 433.050 964.050 ;
        RECT 442.950 963.600 445.050 964.200 ;
        RECT 430.950 962.400 445.050 963.600 ;
        RECT 430.950 961.950 433.050 962.400 ;
        RECT 442.950 962.100 445.050 962.400 ;
        RECT 448.950 962.100 451.050 964.200 ;
        RECT 478.950 963.750 481.050 964.200 ;
        RECT 484.950 963.750 487.050 964.200 ;
        RECT 478.950 962.550 487.050 963.750 ;
        RECT 478.950 962.100 481.050 962.550 ;
        RECT 484.950 962.100 487.050 962.550 ;
        RECT 499.950 963.750 502.050 964.200 ;
        RECT 505.950 963.750 508.050 964.200 ;
        RECT 499.950 962.550 508.050 963.750 ;
        RECT 499.950 962.100 502.050 962.550 ;
        RECT 505.950 962.100 508.050 962.550 ;
        RECT 541.950 963.600 544.050 964.200 ;
        RECT 562.950 963.600 565.050 964.200 ;
        RECT 541.950 962.400 565.050 963.600 ;
        RECT 541.950 962.100 544.050 962.400 ;
        RECT 562.950 962.100 565.050 962.400 ;
        RECT 568.950 963.600 571.050 964.200 ;
        RECT 580.950 963.600 583.050 964.050 ;
        RECT 586.950 963.600 589.050 964.200 ;
        RECT 568.950 962.400 583.050 963.600 ;
        RECT 568.950 962.100 571.050 962.400 ;
        RECT 394.950 957.450 397.050 957.900 ;
        RECT 406.950 957.450 409.050 957.900 ;
        RECT 394.950 956.250 409.050 957.450 ;
        RECT 394.950 955.800 397.050 956.250 ;
        RECT 406.950 955.800 409.050 956.250 ;
        RECT 424.950 957.600 427.050 957.900 ;
        RECT 449.400 957.600 450.600 962.100 ;
        RECT 580.950 961.950 583.050 962.400 ;
        RECT 584.400 962.400 589.050 963.600 ;
        RECT 526.950 960.600 529.050 961.050 ;
        RECT 584.400 960.600 585.600 962.400 ;
        RECT 586.950 962.100 589.050 962.400 ;
        RECT 604.950 963.600 607.050 964.050 ;
        RECT 613.950 963.600 616.050 964.200 ;
        RECT 604.950 962.400 616.050 963.600 ;
        RECT 604.950 961.950 607.050 962.400 ;
        RECT 613.950 962.100 616.050 962.400 ;
        RECT 640.950 963.600 643.050 964.200 ;
        RECT 655.950 963.600 658.050 964.050 ;
        RECT 640.950 962.400 658.050 963.600 ;
        RECT 640.950 962.100 643.050 962.400 ;
        RECT 655.950 961.950 658.050 962.400 ;
        RECT 670.950 963.600 673.050 964.200 ;
        RECT 676.950 963.600 679.050 964.050 ;
        RECT 691.950 963.600 694.050 964.200 ;
        RECT 670.950 962.400 675.600 963.600 ;
        RECT 670.950 962.100 673.050 962.400 ;
        RECT 526.950 959.400 585.600 960.600 ;
        RECT 674.400 960.600 675.600 962.400 ;
        RECT 676.950 962.400 694.050 963.600 ;
        RECT 676.950 961.950 679.050 962.400 ;
        RECT 691.950 962.100 694.050 962.400 ;
        RECT 703.950 963.600 706.050 964.050 ;
        RECT 712.950 963.600 715.050 964.200 ;
        RECT 703.950 962.400 715.050 963.600 ;
        RECT 703.950 961.950 706.050 962.400 ;
        RECT 712.950 962.100 715.050 962.400 ;
        RECT 748.950 963.750 751.050 964.200 ;
        RECT 760.950 963.750 763.050 964.200 ;
        RECT 748.950 962.550 763.050 963.750 ;
        RECT 748.950 962.100 751.050 962.550 ;
        RECT 760.950 962.100 763.050 962.550 ;
        RECT 766.950 963.750 769.050 964.200 ;
        RECT 772.950 963.750 775.050 964.200 ;
        RECT 766.950 962.550 775.050 963.750 ;
        RECT 766.950 962.100 769.050 962.550 ;
        RECT 772.950 962.100 775.050 962.550 ;
        RECT 778.950 963.750 781.050 964.200 ;
        RECT 787.950 963.750 790.050 964.200 ;
        RECT 778.950 962.550 790.050 963.750 ;
        RECT 778.950 962.100 781.050 962.550 ;
        RECT 787.950 962.100 790.050 962.550 ;
        RECT 793.950 962.100 796.050 964.200 ;
        RECT 817.950 962.100 820.050 964.200 ;
        RECT 826.950 963.600 829.050 964.050 ;
        RECT 844.950 963.600 847.050 964.200 ;
        RECT 859.950 963.600 862.050 964.050 ;
        RECT 826.950 962.400 862.050 963.600 ;
        RECT 775.950 960.600 778.050 961.050 ;
        RECT 794.400 960.600 795.600 962.100 ;
        RECT 674.400 959.400 690.600 960.600 ;
        RECT 526.950 958.950 529.050 959.400 ;
        RECT 424.950 956.400 450.600 957.600 ;
        RECT 484.950 957.600 487.050 958.050 ;
        RECT 539.400 957.900 540.600 959.400 ;
        RECT 689.400 957.900 690.600 959.400 ;
        RECT 775.950 959.400 795.600 960.600 ;
        RECT 818.400 960.600 819.600 962.100 ;
        RECT 826.950 961.950 829.050 962.400 ;
        RECT 844.950 962.100 847.050 962.400 ;
        RECT 859.950 961.950 862.050 962.400 ;
        RECT 868.950 963.600 871.050 964.200 ;
        RECT 883.950 963.600 886.050 964.050 ;
        RECT 868.950 962.400 886.050 963.600 ;
        RECT 868.950 962.100 871.050 962.400 ;
        RECT 883.950 961.950 886.050 962.400 ;
        RECT 892.950 963.600 895.050 964.200 ;
        RECT 907.950 963.600 910.050 964.050 ;
        RECT 892.950 962.400 910.050 963.600 ;
        RECT 892.950 962.100 895.050 962.400 ;
        RECT 907.950 961.950 910.050 962.400 ;
        RECT 919.950 963.600 922.050 964.200 ;
        RECT 931.800 963.600 933.900 964.050 ;
        RECT 919.950 962.400 933.900 963.600 ;
        RECT 919.950 962.100 922.050 962.400 ;
        RECT 931.800 961.950 933.900 962.400 ;
        RECT 934.950 963.750 937.050 964.200 ;
        RECT 943.950 963.750 946.050 964.200 ;
        RECT 934.950 962.550 946.050 963.750 ;
        RECT 934.950 962.100 937.050 962.550 ;
        RECT 943.950 962.100 946.050 962.550 ;
        RECT 988.950 963.750 991.050 964.200 ;
        RECT 997.950 963.750 1000.050 964.200 ;
        RECT 988.950 962.550 1000.050 963.750 ;
        RECT 988.950 962.100 991.050 962.550 ;
        RECT 997.950 962.100 1000.050 962.550 ;
        RECT 1006.950 963.750 1009.050 964.200 ;
        RECT 1012.950 963.750 1015.050 964.200 ;
        RECT 1006.950 962.550 1015.050 963.750 ;
        RECT 1006.950 962.100 1009.050 962.550 ;
        RECT 1012.950 962.100 1015.050 962.550 ;
        RECT 818.400 959.400 846.600 960.600 ;
        RECT 775.950 958.950 778.050 959.400 ;
        RECT 496.950 957.600 499.050 957.900 ;
        RECT 484.950 956.400 499.050 957.600 ;
        RECT 424.950 955.800 427.050 956.400 ;
        RECT 484.950 955.950 487.050 956.400 ;
        RECT 496.950 955.800 499.050 956.400 ;
        RECT 538.950 955.800 541.050 957.900 ;
        RECT 565.950 957.600 568.050 957.900 ;
        RECT 589.950 957.600 592.050 957.900 ;
        RECT 565.950 956.400 592.050 957.600 ;
        RECT 565.950 955.800 568.050 956.400 ;
        RECT 589.950 955.800 592.050 956.400 ;
        RECT 655.950 957.450 658.050 957.900 ;
        RECT 661.950 957.450 664.050 957.900 ;
        RECT 655.950 956.250 664.050 957.450 ;
        RECT 655.950 955.800 658.050 956.250 ;
        RECT 661.950 955.800 664.050 956.250 ;
        RECT 688.950 955.800 691.050 957.900 ;
        RECT 763.950 957.600 766.050 957.900 ;
        RECT 778.950 957.600 781.050 958.050 ;
        RECT 763.950 956.400 781.050 957.600 ;
        RECT 763.950 955.800 766.050 956.400 ;
        RECT 778.950 955.950 781.050 956.400 ;
        RECT 796.950 957.600 799.050 957.900 ;
        RECT 814.950 957.600 817.050 957.900 ;
        RECT 796.950 956.400 817.050 957.600 ;
        RECT 796.950 955.800 799.050 956.400 ;
        RECT 814.950 955.800 817.050 956.400 ;
        RECT 823.950 957.600 826.050 957.900 ;
        RECT 841.950 957.600 844.050 957.900 ;
        RECT 823.950 956.400 844.050 957.600 ;
        RECT 845.400 957.600 846.600 959.400 ;
        RECT 847.950 957.600 850.050 957.900 ;
        RECT 845.400 956.400 850.050 957.600 ;
        RECT 823.950 955.800 826.050 956.400 ;
        RECT 841.950 955.800 844.050 956.400 ;
        RECT 847.950 955.800 850.050 956.400 ;
        RECT 883.950 957.450 886.050 957.900 ;
        RECT 889.950 957.450 892.050 957.900 ;
        RECT 883.950 956.250 892.050 957.450 ;
        RECT 883.950 955.800 886.050 956.250 ;
        RECT 889.950 955.800 892.050 956.250 ;
        RECT 931.950 957.450 934.050 957.900 ;
        RECT 940.950 957.450 943.050 957.900 ;
        RECT 931.950 956.250 943.050 957.450 ;
        RECT 931.950 955.800 934.050 956.250 ;
        RECT 940.950 955.800 943.050 956.250 ;
        RECT 1000.950 957.450 1003.050 957.900 ;
        RECT 1009.950 957.450 1012.050 957.900 ;
        RECT 1000.950 956.250 1012.050 957.450 ;
        RECT 1000.950 955.800 1003.050 956.250 ;
        RECT 1009.950 955.800 1012.050 956.250 ;
        RECT 370.950 954.600 373.050 955.050 ;
        RECT 379.950 954.600 382.050 955.050 ;
        RECT 370.950 953.400 382.050 954.600 ;
        RECT 370.950 952.950 373.050 953.400 ;
        RECT 379.950 952.950 382.050 953.400 ;
        RECT 544.950 954.600 547.050 955.050 ;
        RECT 598.950 954.600 601.050 955.050 ;
        RECT 544.950 953.400 601.050 954.600 ;
        RECT 544.950 952.950 547.050 953.400 ;
        RECT 598.950 952.950 601.050 953.400 ;
        RECT 631.950 954.600 634.050 955.050 ;
        RECT 637.950 954.600 640.050 955.050 ;
        RECT 631.950 953.400 640.050 954.600 ;
        RECT 631.950 952.950 634.050 953.400 ;
        RECT 637.950 952.950 640.050 953.400 ;
        RECT 904.950 954.600 907.050 955.050 ;
        RECT 922.950 954.600 925.050 955.050 ;
        RECT 955.950 954.600 958.050 955.050 ;
        RECT 904.950 953.400 958.050 954.600 ;
        RECT 904.950 952.950 907.050 953.400 ;
        RECT 922.950 952.950 925.050 953.400 ;
        RECT 955.950 952.950 958.050 953.400 ;
        RECT 130.950 951.600 133.050 952.050 ;
        RECT 136.950 951.600 139.050 952.050 ;
        RECT 199.950 951.600 202.050 952.050 ;
        RECT 205.950 951.600 208.050 952.050 ;
        RECT 130.950 950.400 208.050 951.600 ;
        RECT 130.950 949.950 133.050 950.400 ;
        RECT 136.950 949.950 139.050 950.400 ;
        RECT 199.950 949.950 202.050 950.400 ;
        RECT 205.950 949.950 208.050 950.400 ;
        RECT 415.950 951.600 418.050 952.050 ;
        RECT 445.950 951.600 448.050 952.050 ;
        RECT 415.950 950.400 448.050 951.600 ;
        RECT 415.950 949.950 418.050 950.400 ;
        RECT 445.950 949.950 448.050 950.400 ;
        RECT 472.950 951.600 475.050 952.050 ;
        RECT 559.950 951.600 562.050 952.050 ;
        RECT 472.950 950.400 562.050 951.600 ;
        RECT 472.950 949.950 475.050 950.400 ;
        RECT 559.950 949.950 562.050 950.400 ;
        RECT 580.950 951.600 583.050 952.050 ;
        RECT 595.950 951.600 598.050 952.050 ;
        RECT 580.950 950.400 598.050 951.600 ;
        RECT 580.950 949.950 583.050 950.400 ;
        RECT 595.950 949.950 598.050 950.400 ;
        RECT 814.950 951.600 817.050 952.050 ;
        RECT 895.950 951.600 898.050 952.050 ;
        RECT 814.950 950.400 898.050 951.600 ;
        RECT 814.950 949.950 817.050 950.400 ;
        RECT 895.950 949.950 898.050 950.400 ;
        RECT 52.950 948.600 55.050 949.050 ;
        RECT 85.950 948.600 88.050 949.050 ;
        RECT 52.950 947.400 88.050 948.600 ;
        RECT 52.950 946.950 55.050 947.400 ;
        RECT 85.950 946.950 88.050 947.400 ;
        RECT 346.950 948.600 349.050 949.050 ;
        RECT 424.950 948.600 427.050 949.050 ;
        RECT 346.950 947.400 427.050 948.600 ;
        RECT 346.950 946.950 349.050 947.400 ;
        RECT 424.950 946.950 427.050 947.400 ;
        RECT 448.950 948.600 451.050 949.050 ;
        RECT 469.950 948.600 472.050 949.050 ;
        RECT 517.950 948.600 520.050 949.050 ;
        RECT 448.950 947.400 520.050 948.600 ;
        RECT 448.950 946.950 451.050 947.400 ;
        RECT 469.950 946.950 472.050 947.400 ;
        RECT 517.950 946.950 520.050 947.400 ;
        RECT 604.950 948.600 607.050 949.050 ;
        RECT 667.950 948.600 670.050 949.050 ;
        RECT 604.950 947.400 670.050 948.600 ;
        RECT 604.950 946.950 607.050 947.400 ;
        RECT 667.950 946.950 670.050 947.400 ;
        RECT 739.950 948.600 742.050 949.050 ;
        RECT 784.950 948.600 787.050 949.050 ;
        RECT 739.950 947.400 787.050 948.600 ;
        RECT 739.950 946.950 742.050 947.400 ;
        RECT 784.950 946.950 787.050 947.400 ;
        RECT 880.950 948.600 883.050 949.050 ;
        RECT 1012.950 948.600 1015.050 949.050 ;
        RECT 880.950 947.400 1015.050 948.600 ;
        RECT 880.950 946.950 883.050 947.400 ;
        RECT 1012.950 946.950 1015.050 947.400 ;
        RECT 619.950 945.600 622.050 946.050 ;
        RECT 643.950 945.600 646.050 946.050 ;
        RECT 619.950 944.400 646.050 945.600 ;
        RECT 619.950 943.950 622.050 944.400 ;
        RECT 643.950 943.950 646.050 944.400 ;
        RECT 694.950 945.600 697.050 946.050 ;
        RECT 790.950 945.600 793.050 946.050 ;
        RECT 694.950 944.400 793.050 945.600 ;
        RECT 694.950 943.950 697.050 944.400 ;
        RECT 790.950 943.950 793.050 944.400 ;
        RECT 868.950 945.600 871.050 946.050 ;
        RECT 934.950 945.600 937.050 946.050 ;
        RECT 868.950 944.400 937.050 945.600 ;
        RECT 868.950 943.950 871.050 944.400 ;
        RECT 934.950 943.950 937.050 944.400 ;
        RECT 85.950 942.600 88.050 943.050 ;
        RECT 145.950 942.600 148.050 943.050 ;
        RECT 214.950 942.600 217.050 943.050 ;
        RECT 85.950 941.400 217.050 942.600 ;
        RECT 85.950 940.950 88.050 941.400 ;
        RECT 145.950 940.950 148.050 941.400 ;
        RECT 214.950 940.950 217.050 941.400 ;
        RECT 277.950 942.600 280.050 943.050 ;
        RECT 313.950 942.600 316.050 943.050 ;
        RECT 277.950 941.400 316.050 942.600 ;
        RECT 277.950 940.950 280.050 941.400 ;
        RECT 313.950 940.950 316.050 941.400 ;
        RECT 328.950 942.600 331.050 943.050 ;
        RECT 715.950 942.600 718.050 943.050 ;
        RECT 775.950 942.600 778.050 943.050 ;
        RECT 328.950 941.400 423.600 942.600 ;
        RECT 328.950 940.950 331.050 941.400 ;
        RECT 422.400 940.050 423.600 941.400 ;
        RECT 715.950 941.400 778.050 942.600 ;
        RECT 715.950 940.950 718.050 941.400 ;
        RECT 775.950 940.950 778.050 941.400 ;
        RECT 796.950 942.600 799.050 943.050 ;
        RECT 823.950 942.600 826.050 943.050 ;
        RECT 796.950 941.400 826.050 942.600 ;
        RECT 796.950 940.950 799.050 941.400 ;
        RECT 823.950 940.950 826.050 941.400 ;
        RECT 853.950 942.600 856.050 943.050 ;
        RECT 853.950 941.400 933.600 942.600 ;
        RECT 853.950 940.950 856.050 941.400 ;
        RECT 268.950 939.600 271.050 940.050 ;
        RECT 364.950 939.600 367.050 940.050 ;
        RECT 268.950 938.400 367.050 939.600 ;
        RECT 268.950 937.950 271.050 938.400 ;
        RECT 364.950 937.950 367.050 938.400 ;
        RECT 421.950 939.600 424.050 940.050 ;
        RECT 475.950 939.600 478.050 940.050 ;
        RECT 505.950 939.600 508.050 940.050 ;
        RECT 601.950 939.600 604.050 940.050 ;
        RECT 421.950 938.400 604.050 939.600 ;
        RECT 932.400 939.600 933.600 941.400 ;
        RECT 946.950 939.600 949.050 940.050 ;
        RECT 932.400 938.400 949.050 939.600 ;
        RECT 421.950 937.950 424.050 938.400 ;
        RECT 475.950 937.950 478.050 938.400 ;
        RECT 505.950 937.950 508.050 938.400 ;
        RECT 601.950 937.950 604.050 938.400 ;
        RECT 946.950 937.950 949.050 938.400 ;
        RECT 100.950 936.600 103.050 937.050 ;
        RECT 106.950 936.600 109.050 937.050 ;
        RECT 100.950 935.400 109.050 936.600 ;
        RECT 100.950 934.950 103.050 935.400 ;
        RECT 106.950 934.950 109.050 935.400 ;
        RECT 700.950 936.600 703.050 937.050 ;
        RECT 826.950 936.600 829.050 937.050 ;
        RECT 700.950 935.400 829.050 936.600 ;
        RECT 700.950 934.950 703.050 935.400 ;
        RECT 826.950 934.950 829.050 935.400 ;
        RECT 859.950 936.600 862.050 937.050 ;
        RECT 883.950 936.600 886.050 937.050 ;
        RECT 916.950 936.600 919.050 937.050 ;
        RECT 859.950 935.400 919.050 936.600 ;
        RECT 859.950 934.950 862.050 935.400 ;
        RECT 883.950 934.950 886.050 935.400 ;
        RECT 916.950 934.950 919.050 935.400 ;
        RECT 121.950 933.600 124.050 934.050 ;
        RECT 139.950 933.600 142.050 934.050 ;
        RECT 121.950 932.400 142.050 933.600 ;
        RECT 121.950 931.950 124.050 932.400 ;
        RECT 139.950 931.950 142.050 932.400 ;
        RECT 214.950 933.600 217.050 934.050 ;
        RECT 283.950 933.600 286.050 934.050 ;
        RECT 214.950 932.400 286.050 933.600 ;
        RECT 214.950 931.950 217.050 932.400 ;
        RECT 283.950 931.950 286.050 932.400 ;
        RECT 331.950 933.600 334.050 934.050 ;
        RECT 478.950 933.600 481.050 934.050 ;
        RECT 721.950 933.600 724.050 934.050 ;
        RECT 331.950 932.400 481.050 933.600 ;
        RECT 331.950 931.950 334.050 932.400 ;
        RECT 478.950 931.950 481.050 932.400 ;
        RECT 704.400 932.400 724.050 933.600 ;
        RECT 145.950 930.600 148.050 931.050 ;
        RECT 160.950 930.600 163.050 931.050 ;
        RECT 145.950 929.400 163.050 930.600 ;
        RECT 145.950 928.950 148.050 929.400 ;
        RECT 160.950 928.950 163.050 929.400 ;
        RECT 259.950 930.600 262.050 931.050 ;
        RECT 328.950 930.600 331.050 931.050 ;
        RECT 259.950 929.400 279.600 930.600 ;
        RECT 259.950 928.950 262.050 929.400 ;
        RECT 184.950 927.600 187.050 928.050 ;
        RECT 226.950 927.600 229.050 928.050 ;
        RECT 184.950 926.400 229.050 927.600 ;
        RECT 278.400 927.600 279.600 929.400 ;
        RECT 287.400 929.400 331.050 930.600 ;
        RECT 287.400 927.600 288.600 929.400 ;
        RECT 328.950 928.950 331.050 929.400 ;
        RECT 364.950 930.600 367.050 931.050 ;
        RECT 466.950 930.600 469.050 931.050 ;
        RECT 364.950 929.400 469.050 930.600 ;
        RECT 364.950 928.950 367.050 929.400 ;
        RECT 466.950 928.950 469.050 929.400 ;
        RECT 595.950 930.600 598.050 931.050 ;
        RECT 704.400 930.600 705.600 932.400 ;
        RECT 721.950 931.950 724.050 932.400 ;
        RECT 727.950 933.600 730.050 934.050 ;
        RECT 778.950 933.600 781.050 934.050 ;
        RECT 784.950 933.600 787.050 934.050 ;
        RECT 727.950 932.400 787.050 933.600 ;
        RECT 727.950 931.950 730.050 932.400 ;
        RECT 778.950 931.950 781.050 932.400 ;
        RECT 784.950 931.950 787.050 932.400 ;
        RECT 817.950 933.600 820.050 934.050 ;
        RECT 853.950 933.600 856.050 934.050 ;
        RECT 817.950 932.400 856.050 933.600 ;
        RECT 817.950 931.950 820.050 932.400 ;
        RECT 853.950 931.950 856.050 932.400 ;
        RECT 595.950 929.400 705.600 930.600 ;
        RECT 865.950 930.600 868.050 931.050 ;
        RECT 877.950 930.600 880.050 931.050 ;
        RECT 865.950 929.400 880.050 930.600 ;
        RECT 595.950 928.950 598.050 929.400 ;
        RECT 865.950 928.950 868.050 929.400 ;
        RECT 877.950 928.950 880.050 929.400 ;
        RECT 278.400 926.400 288.600 927.600 ;
        RECT 343.950 927.600 346.050 928.050 ;
        RECT 361.950 927.600 364.050 928.050 ;
        RECT 343.950 926.400 364.050 927.600 ;
        RECT 184.950 925.950 187.050 926.400 ;
        RECT 226.950 925.950 229.050 926.400 ;
        RECT 343.950 925.950 346.050 926.400 ;
        RECT 361.950 925.950 364.050 926.400 ;
        RECT 499.950 927.600 502.050 928.050 ;
        RECT 649.950 927.600 652.050 928.050 ;
        RECT 499.950 926.400 652.050 927.600 ;
        RECT 499.950 925.950 502.050 926.400 ;
        RECT 649.950 925.950 652.050 926.400 ;
        RECT 706.950 927.600 709.050 928.050 ;
        RECT 715.950 927.600 718.050 928.050 ;
        RECT 706.950 926.400 718.050 927.600 ;
        RECT 706.950 925.950 709.050 926.400 ;
        RECT 715.950 925.950 718.050 926.400 ;
        RECT 766.950 927.600 769.050 928.050 ;
        RECT 799.950 927.600 802.050 928.050 ;
        RECT 766.950 926.400 802.050 927.600 ;
        RECT 766.950 925.950 769.050 926.400 ;
        RECT 799.950 925.950 802.050 926.400 ;
        RECT 808.950 927.600 811.050 928.050 ;
        RECT 856.950 927.600 859.050 928.050 ;
        RECT 808.950 926.400 859.050 927.600 ;
        RECT 808.950 925.950 811.050 926.400 ;
        RECT 856.950 925.950 859.050 926.400 ;
        RECT 973.950 927.600 976.050 928.050 ;
        RECT 991.950 927.600 994.050 928.050 ;
        RECT 973.950 926.400 994.050 927.600 ;
        RECT 973.950 925.950 976.050 926.400 ;
        RECT 991.950 925.950 994.050 926.400 ;
        RECT 151.950 924.600 154.050 925.050 ;
        RECT 223.950 924.600 226.050 925.050 ;
        RECT 274.950 924.600 277.050 925.050 ;
        RECT 298.950 924.600 301.050 925.050 ;
        RECT 151.950 923.400 301.050 924.600 ;
        RECT 151.950 922.950 154.050 923.400 ;
        RECT 223.950 922.950 226.050 923.400 ;
        RECT 274.950 922.950 277.050 923.400 ;
        RECT 298.950 922.950 301.050 923.400 ;
        RECT 340.950 924.600 343.050 925.050 ;
        RECT 379.950 924.600 382.050 925.050 ;
        RECT 400.950 924.600 403.050 925.050 ;
        RECT 340.950 923.400 403.050 924.600 ;
        RECT 340.950 922.950 343.050 923.400 ;
        RECT 379.950 922.950 382.050 923.400 ;
        RECT 400.950 922.950 403.050 923.400 ;
        RECT 406.950 924.600 409.050 925.050 ;
        RECT 418.950 924.600 421.050 925.050 ;
        RECT 496.950 924.600 499.050 925.050 ;
        RECT 406.950 923.400 499.050 924.600 ;
        RECT 406.950 922.950 409.050 923.400 ;
        RECT 418.950 922.950 421.050 923.400 ;
        RECT 496.950 922.950 499.050 923.400 ;
        RECT 583.950 924.600 586.050 925.050 ;
        RECT 634.950 924.600 637.050 925.050 ;
        RECT 583.950 923.400 637.050 924.600 ;
        RECT 583.950 922.950 586.050 923.400 ;
        RECT 634.950 922.950 637.050 923.400 ;
        RECT 643.950 924.600 646.050 925.050 ;
        RECT 715.950 924.600 718.050 924.900 ;
        RECT 643.950 923.400 718.050 924.600 ;
        RECT 643.950 922.950 646.050 923.400 ;
        RECT 715.950 922.800 718.050 923.400 ;
        RECT 721.950 924.600 724.050 925.050 ;
        RECT 775.950 924.600 778.050 925.050 ;
        RECT 721.950 923.400 778.050 924.600 ;
        RECT 721.950 922.950 724.050 923.400 ;
        RECT 775.950 922.950 778.050 923.400 ;
        RECT 889.950 924.600 892.050 925.050 ;
        RECT 904.950 924.600 907.050 925.050 ;
        RECT 889.950 923.400 907.050 924.600 ;
        RECT 889.950 922.950 892.050 923.400 ;
        RECT 904.950 922.950 907.050 923.400 ;
        RECT 1006.950 924.600 1009.050 925.050 ;
        RECT 1027.950 924.600 1030.050 925.050 ;
        RECT 1006.950 923.400 1030.050 924.600 ;
        RECT 1006.950 922.950 1009.050 923.400 ;
        RECT 1027.950 922.950 1030.050 923.400 ;
        RECT 124.950 921.600 127.050 922.050 ;
        RECT 133.950 921.600 136.050 922.050 ;
        RECT 124.950 920.400 136.050 921.600 ;
        RECT 124.950 919.950 127.050 920.400 ;
        RECT 133.950 919.950 136.050 920.400 ;
        RECT 169.950 921.600 172.050 922.050 ;
        RECT 214.950 921.600 217.050 922.050 ;
        RECT 169.950 920.400 217.050 921.600 ;
        RECT 169.950 919.950 172.050 920.400 ;
        RECT 214.950 919.950 217.050 920.400 ;
        RECT 244.950 921.600 247.050 922.050 ;
        RECT 256.950 921.600 259.050 922.050 ;
        RECT 244.950 920.400 259.050 921.600 ;
        RECT 244.950 919.950 247.050 920.400 ;
        RECT 256.950 919.950 259.050 920.400 ;
        RECT 304.950 921.600 307.050 922.050 ;
        RECT 346.950 921.600 349.050 922.050 ;
        RECT 304.950 920.400 349.050 921.600 ;
        RECT 304.950 919.950 307.050 920.400 ;
        RECT 346.950 919.950 349.050 920.400 ;
        RECT 724.950 921.600 727.050 922.050 ;
        RECT 739.950 921.600 742.050 922.050 ;
        RECT 724.950 920.400 742.050 921.600 ;
        RECT 724.950 919.950 727.050 920.400 ;
        RECT 739.950 919.950 742.050 920.400 ;
        RECT 952.950 921.600 955.050 922.050 ;
        RECT 991.950 921.600 994.050 922.050 ;
        RECT 952.950 920.400 994.050 921.600 ;
        RECT 952.950 919.950 955.050 920.400 ;
        RECT 991.950 919.950 994.050 920.400 ;
        RECT 25.950 918.750 28.050 919.200 ;
        RECT 37.950 918.750 40.050 919.200 ;
        RECT 25.950 917.550 40.050 918.750 ;
        RECT 25.950 917.100 28.050 917.550 ;
        RECT 37.950 917.100 40.050 917.550 ;
        RECT 79.950 918.750 82.050 919.200 ;
        RECT 97.950 918.750 100.050 919.200 ;
        RECT 79.950 917.550 100.050 918.750 ;
        RECT 79.950 917.100 82.050 917.550 ;
        RECT 97.950 917.100 100.050 917.550 ;
        RECT 118.950 917.100 121.050 919.200 ;
        RECT 139.950 918.750 142.050 919.200 ;
        RECT 145.950 918.750 148.050 919.200 ;
        RECT 139.950 917.550 148.050 918.750 ;
        RECT 268.950 918.600 271.050 919.200 ;
        RECT 139.950 917.100 142.050 917.550 ;
        RECT 145.950 917.100 148.050 917.550 ;
        RECT 227.400 917.400 271.050 918.600 ;
        RECT 119.400 915.600 120.600 917.100 ;
        RECT 220.950 915.600 223.050 915.900 ;
        RECT 227.400 915.600 228.600 917.400 ;
        RECT 268.950 917.100 271.050 917.400 ;
        RECT 325.950 918.750 328.050 919.200 ;
        RECT 340.950 918.750 343.050 919.200 ;
        RECT 325.950 917.550 343.050 918.750 ;
        RECT 325.950 917.100 328.050 917.550 ;
        RECT 340.950 917.100 343.050 917.550 ;
        RECT 352.950 918.600 355.050 919.200 ;
        RECT 385.950 918.600 388.050 919.050 ;
        RECT 430.950 918.600 433.050 919.050 ;
        RECT 352.950 917.400 381.600 918.600 ;
        RECT 352.950 917.100 355.050 917.400 ;
        RECT 119.400 914.400 129.600 915.600 ;
        RECT 37.950 912.450 40.050 912.900 ;
        RECT 46.950 912.450 49.050 912.900 ;
        RECT 37.950 911.250 49.050 912.450 ;
        RECT 37.950 910.800 40.050 911.250 ;
        RECT 46.950 910.800 49.050 911.250 ;
        RECT 106.950 912.600 109.050 913.050 ;
        RECT 121.950 912.600 124.050 912.900 ;
        RECT 106.950 911.400 124.050 912.600 ;
        RECT 128.400 912.600 129.600 914.400 ;
        RECT 220.950 914.400 228.600 915.600 ;
        RECT 380.400 915.600 381.600 917.400 ;
        RECT 385.950 917.400 433.050 918.600 ;
        RECT 385.950 916.950 388.050 917.400 ;
        RECT 430.950 916.950 433.050 917.400 ;
        RECT 439.950 918.600 442.050 919.200 ;
        RECT 460.950 918.600 463.050 919.200 ;
        RECT 439.950 917.400 463.050 918.600 ;
        RECT 439.950 917.100 442.050 917.400 ;
        RECT 460.950 917.100 463.050 917.400 ;
        RECT 466.950 918.600 469.050 919.200 ;
        RECT 490.950 918.750 493.050 919.200 ;
        RECT 496.950 918.750 499.050 919.200 ;
        RECT 490.950 918.600 499.050 918.750 ;
        RECT 466.950 917.550 499.050 918.600 ;
        RECT 466.950 917.400 493.050 917.550 ;
        RECT 466.950 917.100 469.050 917.400 ;
        RECT 490.950 917.100 493.050 917.400 ;
        RECT 496.950 917.100 499.050 917.550 ;
        RECT 511.950 918.600 514.050 919.200 ;
        RECT 532.950 918.600 535.050 919.200 ;
        RECT 511.950 917.400 535.050 918.600 ;
        RECT 511.950 917.100 514.050 917.400 ;
        RECT 532.950 917.100 535.050 917.400 ;
        RECT 538.950 918.750 541.050 919.200 ;
        RECT 547.950 918.750 550.050 919.200 ;
        RECT 538.950 917.550 550.050 918.750 ;
        RECT 538.950 917.100 541.050 917.550 ;
        RECT 547.950 917.100 550.050 917.550 ;
        RECT 553.950 918.600 556.050 919.050 ;
        RECT 562.950 918.600 565.050 919.200 ;
        RECT 553.950 917.400 565.050 918.600 ;
        RECT 553.950 916.950 556.050 917.400 ;
        RECT 562.950 917.100 565.050 917.400 ;
        RECT 589.950 917.100 592.050 919.200 ;
        RECT 610.950 918.600 613.050 919.200 ;
        RECT 625.950 918.600 628.050 919.050 ;
        RECT 610.950 917.400 628.050 918.600 ;
        RECT 610.950 917.100 613.050 917.400 ;
        RECT 380.400 914.400 402.600 915.600 ;
        RECT 220.950 913.800 223.050 914.400 ;
        RECT 148.950 912.600 151.050 912.900 ;
        RECT 128.400 911.400 151.050 912.600 ;
        RECT 106.950 910.950 109.050 911.400 ;
        RECT 121.950 910.800 124.050 911.400 ;
        RECT 148.950 910.800 151.050 911.400 ;
        RECT 226.950 912.600 229.050 913.050 ;
        RECT 247.950 912.600 250.050 912.900 ;
        RECT 226.950 911.400 250.050 912.600 ;
        RECT 226.950 910.950 229.050 911.400 ;
        RECT 247.950 910.800 250.050 911.400 ;
        RECT 259.950 912.600 262.050 913.050 ;
        RECT 271.950 912.600 274.050 912.900 ;
        RECT 259.950 911.400 274.050 912.600 ;
        RECT 259.950 910.950 262.050 911.400 ;
        RECT 271.950 910.800 274.050 911.400 ;
        RECT 277.950 912.600 280.050 912.900 ;
        RECT 295.950 912.600 298.050 912.900 ;
        RECT 277.950 911.400 298.050 912.600 ;
        RECT 277.950 910.800 280.050 911.400 ;
        RECT 295.950 910.800 298.050 911.400 ;
        RECT 301.950 912.600 304.050 912.900 ;
        RECT 343.950 912.600 346.050 913.050 ;
        RECT 401.400 912.900 402.600 914.400 ;
        RECT 590.400 913.050 591.600 917.100 ;
        RECT 625.950 916.950 628.050 917.400 ;
        RECT 646.950 918.750 649.050 919.200 ;
        RECT 658.950 918.750 661.050 919.200 ;
        RECT 646.950 917.550 661.050 918.750 ;
        RECT 646.950 917.100 649.050 917.550 ;
        RECT 658.950 917.100 661.050 917.550 ;
        RECT 676.950 918.750 679.050 918.900 ;
        RECT 682.950 918.750 685.050 919.200 ;
        RECT 676.950 917.550 685.050 918.750 ;
        RECT 688.950 918.600 691.050 919.200 ;
        RECT 676.950 916.800 679.050 917.550 ;
        RECT 682.950 917.100 685.050 917.550 ;
        RECT 686.400 917.400 691.050 918.600 ;
        RECT 686.400 915.600 687.600 917.400 ;
        RECT 688.950 917.100 691.050 917.400 ;
        RECT 694.950 918.750 697.050 919.200 ;
        RECT 703.950 918.750 706.050 919.200 ;
        RECT 694.950 917.550 706.050 918.750 ;
        RECT 694.950 917.100 697.050 917.550 ;
        RECT 703.950 917.100 706.050 917.550 ;
        RECT 748.950 918.750 751.050 919.200 ;
        RECT 760.950 918.750 763.050 919.200 ;
        RECT 748.950 917.550 763.050 918.750 ;
        RECT 748.950 917.100 751.050 917.550 ;
        RECT 760.950 917.100 763.050 917.550 ;
        RECT 790.950 918.750 793.050 919.200 ;
        RECT 802.950 918.750 805.050 919.200 ;
        RECT 790.950 917.550 805.050 918.750 ;
        RECT 790.950 917.100 793.050 917.550 ;
        RECT 802.950 917.100 805.050 917.550 ;
        RECT 826.950 918.600 829.050 919.050 ;
        RECT 835.950 918.600 838.050 919.200 ;
        RECT 868.950 918.600 871.050 919.200 ;
        RECT 826.950 917.400 838.050 918.600 ;
        RECT 826.950 916.950 829.050 917.400 ;
        RECT 835.950 917.100 838.050 917.400 ;
        RECT 863.400 917.400 871.050 918.600 ;
        RECT 863.400 915.600 864.600 917.400 ;
        RECT 868.950 917.100 871.050 917.400 ;
        RECT 895.950 918.750 898.050 919.200 ;
        RECT 904.950 918.750 907.050 919.200 ;
        RECT 895.950 917.550 907.050 918.750 ;
        RECT 895.950 917.100 898.050 917.550 ;
        RECT 904.950 917.100 907.050 917.550 ;
        RECT 910.950 918.750 913.050 919.200 ;
        RECT 922.950 918.750 925.050 919.200 ;
        RECT 910.950 917.550 925.050 918.750 ;
        RECT 910.950 917.100 913.050 917.550 ;
        RECT 922.950 917.100 925.050 917.550 ;
        RECT 934.950 918.750 937.050 919.200 ;
        RECT 940.950 918.750 943.050 919.200 ;
        RECT 934.950 917.550 943.050 918.750 ;
        RECT 934.950 917.100 937.050 917.550 ;
        RECT 940.950 917.100 943.050 917.550 ;
        RECT 946.950 917.100 949.050 919.200 ;
        RECT 958.950 918.750 961.050 919.200 ;
        RECT 967.950 918.750 970.050 919.200 ;
        RECT 958.950 917.550 970.050 918.750 ;
        RECT 958.950 917.100 961.050 917.550 ;
        RECT 967.950 917.100 970.050 917.550 ;
        RECT 997.950 918.600 1000.050 919.200 ;
        RECT 1021.950 918.600 1024.050 919.200 ;
        RECT 997.950 917.400 1024.050 918.600 ;
        RECT 997.950 917.100 1000.050 917.400 ;
        RECT 1021.950 917.100 1024.050 917.400 ;
        RECT 662.400 914.400 687.600 915.600 ;
        RECT 851.400 914.400 864.600 915.600 ;
        RECT 301.950 911.400 346.050 912.600 ;
        RECT 301.950 910.800 304.050 911.400 ;
        RECT 343.950 910.950 346.050 911.400 ;
        RECT 349.950 912.450 352.050 912.900 ;
        RECT 364.950 912.450 367.050 912.900 ;
        RECT 349.950 911.250 367.050 912.450 ;
        RECT 349.950 910.800 352.050 911.250 ;
        RECT 364.950 910.800 367.050 911.250 ;
        RECT 376.950 912.450 379.050 912.900 ;
        RECT 385.950 912.450 388.050 912.900 ;
        RECT 376.950 911.250 388.050 912.450 ;
        RECT 376.950 910.800 379.050 911.250 ;
        RECT 385.950 910.800 388.050 911.250 ;
        RECT 400.950 910.800 403.050 912.900 ;
        RECT 409.950 912.600 412.050 912.900 ;
        RECT 436.950 912.600 439.050 912.900 ;
        RECT 409.950 911.400 439.050 912.600 ;
        RECT 409.950 910.800 412.050 911.400 ;
        RECT 436.950 910.800 439.050 911.400 ;
        RECT 463.950 912.450 466.050 912.900 ;
        RECT 475.800 912.450 477.900 912.900 ;
        RECT 463.950 911.250 477.900 912.450 ;
        RECT 463.950 910.800 466.050 911.250 ;
        RECT 475.800 910.800 477.900 911.250 ;
        RECT 478.950 912.600 481.050 913.050 ;
        RECT 487.950 912.600 490.050 912.900 ;
        RECT 478.950 911.400 490.050 912.600 ;
        RECT 478.950 910.950 481.050 911.400 ;
        RECT 487.950 910.800 490.050 911.400 ;
        RECT 541.950 912.450 544.050 912.900 ;
        RECT 556.950 912.450 559.050 912.900 ;
        RECT 541.950 911.250 559.050 912.450 ;
        RECT 541.950 910.800 544.050 911.250 ;
        RECT 556.950 910.800 559.050 911.250 ;
        RECT 565.950 912.600 568.050 912.900 ;
        RECT 586.950 912.600 589.050 912.900 ;
        RECT 565.950 911.400 589.050 912.600 ;
        RECT 590.400 911.400 595.050 913.050 ;
        RECT 565.950 910.800 568.050 911.400 ;
        RECT 586.950 910.800 589.050 911.400 ;
        RECT 591.000 910.950 595.050 911.400 ;
        RECT 604.950 912.600 607.050 913.050 ;
        RECT 662.400 912.900 663.600 914.400 ;
        RECT 625.950 912.600 628.050 912.900 ;
        RECT 604.950 912.450 628.050 912.600 ;
        RECT 631.950 912.450 634.050 912.900 ;
        RECT 604.950 911.400 634.050 912.450 ;
        RECT 604.950 910.950 607.050 911.400 ;
        RECT 625.950 911.250 634.050 911.400 ;
        RECT 625.950 910.800 628.050 911.250 ;
        RECT 631.950 910.800 634.050 911.250 ;
        RECT 637.950 912.450 640.050 912.900 ;
        RECT 643.950 912.450 646.050 912.900 ;
        RECT 637.950 911.250 646.050 912.450 ;
        RECT 637.950 910.800 640.050 911.250 ;
        RECT 643.950 910.800 646.050 911.250 ;
        RECT 661.950 910.800 664.050 912.900 ;
        RECT 670.950 912.450 673.050 912.900 ;
        RECT 685.950 912.450 688.050 912.900 ;
        RECT 670.950 911.250 688.050 912.450 ;
        RECT 670.950 910.800 673.050 911.250 ;
        RECT 685.950 910.800 688.050 911.250 ;
        RECT 718.950 912.450 721.050 912.900 ;
        RECT 724.950 912.450 727.050 912.900 ;
        RECT 718.950 911.250 727.050 912.450 ;
        RECT 718.950 910.800 721.050 911.250 ;
        RECT 724.950 910.800 727.050 911.250 ;
        RECT 730.950 912.450 733.050 912.900 ;
        RECT 736.950 912.450 739.050 912.900 ;
        RECT 730.950 911.250 739.050 912.450 ;
        RECT 730.950 910.800 733.050 911.250 ;
        RECT 736.950 910.800 739.050 911.250 ;
        RECT 787.950 912.600 790.050 912.900 ;
        RECT 796.950 912.600 799.050 913.050 ;
        RECT 787.950 911.400 799.050 912.600 ;
        RECT 787.950 910.800 790.050 911.400 ;
        RECT 796.950 910.950 799.050 911.400 ;
        RECT 844.950 912.600 847.050 912.900 ;
        RECT 851.400 912.600 852.600 914.400 ;
        RECT 947.400 913.050 948.600 917.100 ;
        RECT 844.950 911.400 852.600 912.600 ;
        RECT 856.950 912.450 859.050 912.900 ;
        RECT 865.950 912.450 868.050 912.900 ;
        RECT 844.950 910.800 847.050 911.400 ;
        RECT 856.950 911.250 868.050 912.450 ;
        RECT 856.950 910.800 859.050 911.250 ;
        RECT 865.950 910.800 868.050 911.250 ;
        RECT 883.950 912.450 886.050 912.900 ;
        RECT 892.950 912.450 895.050 912.900 ;
        RECT 883.950 911.250 895.050 912.450 ;
        RECT 883.950 910.800 886.050 911.250 ;
        RECT 892.950 910.800 895.050 911.250 ;
        RECT 925.950 912.600 928.050 912.900 ;
        RECT 934.950 912.600 937.050 913.050 ;
        RECT 925.950 911.400 937.050 912.600 ;
        RECT 947.400 911.400 952.050 913.050 ;
        RECT 925.950 910.800 928.050 911.400 ;
        RECT 934.950 910.950 937.050 911.400 ;
        RECT 948.000 910.950 952.050 911.400 ;
        RECT 1012.950 912.450 1015.050 912.900 ;
        RECT 1018.950 912.450 1021.050 912.900 ;
        RECT 1012.950 911.250 1021.050 912.450 ;
        RECT 1012.950 910.800 1015.050 911.250 ;
        RECT 1018.950 910.800 1021.050 911.250 ;
        RECT 61.950 909.600 64.050 910.050 ;
        RECT 73.950 909.600 76.050 910.050 ;
        RECT 61.950 908.400 76.050 909.600 ;
        RECT 61.950 907.950 64.050 908.400 ;
        RECT 73.950 907.950 76.050 908.400 ;
        RECT 157.950 909.600 160.050 910.050 ;
        RECT 646.950 909.600 649.050 910.050 ;
        RECT 655.950 909.600 658.050 910.050 ;
        RECT 157.950 908.400 225.600 909.600 ;
        RECT 157.950 907.950 160.050 908.400 ;
        RECT 139.950 906.600 142.050 907.050 ;
        RECT 148.950 906.600 151.050 907.050 ;
        RECT 139.950 905.400 151.050 906.600 ;
        RECT 139.950 904.950 142.050 905.400 ;
        RECT 148.950 904.950 151.050 905.400 ;
        RECT 154.950 906.600 157.050 907.050 ;
        RECT 163.950 906.600 166.050 907.050 ;
        RECT 154.950 905.400 166.050 906.600 ;
        RECT 154.950 904.950 157.050 905.400 ;
        RECT 163.950 904.950 166.050 905.400 ;
        RECT 205.950 906.600 208.050 907.050 ;
        RECT 211.950 906.600 214.050 907.050 ;
        RECT 220.950 906.600 223.050 907.050 ;
        RECT 205.950 905.400 223.050 906.600 ;
        RECT 224.400 906.600 225.600 908.400 ;
        RECT 646.950 908.400 658.050 909.600 ;
        RECT 646.950 907.950 649.050 908.400 ;
        RECT 655.950 907.950 658.050 908.400 ;
        RECT 691.950 909.600 694.050 910.050 ;
        RECT 700.950 909.600 703.050 910.050 ;
        RECT 691.950 908.400 703.050 909.600 ;
        RECT 691.950 907.950 694.050 908.400 ;
        RECT 700.950 907.950 703.050 908.400 ;
        RECT 757.950 909.600 760.050 910.050 ;
        RECT 772.950 909.600 775.050 910.050 ;
        RECT 757.950 908.400 775.050 909.600 ;
        RECT 757.950 907.950 760.050 908.400 ;
        RECT 772.950 907.950 775.050 908.400 ;
        RECT 799.950 909.600 802.050 910.050 ;
        RECT 823.950 909.600 826.050 910.050 ;
        RECT 799.950 908.400 826.050 909.600 ;
        RECT 799.950 907.950 802.050 908.400 ;
        RECT 823.950 907.950 826.050 908.400 ;
        RECT 994.950 909.600 997.050 910.050 ;
        RECT 1000.950 909.600 1003.050 910.050 ;
        RECT 994.950 908.400 1003.050 909.600 ;
        RECT 994.950 907.950 997.050 908.400 ;
        RECT 1000.950 907.950 1003.050 908.400 ;
        RECT 367.950 906.600 370.050 907.050 ;
        RECT 224.400 905.400 370.050 906.600 ;
        RECT 205.950 904.950 208.050 905.400 ;
        RECT 211.950 904.950 214.050 905.400 ;
        RECT 220.950 904.950 223.050 905.400 ;
        RECT 367.950 904.950 370.050 905.400 ;
        RECT 439.950 906.600 442.050 907.050 ;
        RECT 448.950 906.600 451.050 907.050 ;
        RECT 439.950 905.400 451.050 906.600 ;
        RECT 439.950 904.950 442.050 905.400 ;
        RECT 448.950 904.950 451.050 905.400 ;
        RECT 601.950 906.600 604.050 907.050 ;
        RECT 613.950 906.600 616.050 907.050 ;
        RECT 721.950 906.600 724.050 907.050 ;
        RECT 601.950 905.400 724.050 906.600 ;
        RECT 601.950 904.950 604.050 905.400 ;
        RECT 613.950 904.950 616.050 905.400 ;
        RECT 721.950 904.950 724.050 905.400 ;
        RECT 763.950 906.600 766.050 907.050 ;
        RECT 805.950 906.600 808.050 907.050 ;
        RECT 763.950 905.400 808.050 906.600 ;
        RECT 763.950 904.950 766.050 905.400 ;
        RECT 805.950 904.950 808.050 905.400 ;
        RECT 814.950 906.600 817.050 907.050 ;
        RECT 853.950 906.600 856.050 907.050 ;
        RECT 814.950 905.400 856.050 906.600 ;
        RECT 814.950 904.950 817.050 905.400 ;
        RECT 853.950 904.950 856.050 905.400 ;
        RECT 871.950 906.600 874.050 907.050 ;
        RECT 904.950 906.600 907.050 907.050 ;
        RECT 871.950 905.400 907.050 906.600 ;
        RECT 871.950 904.950 874.050 905.400 ;
        RECT 904.950 904.950 907.050 905.400 ;
        RECT 970.950 906.600 973.050 907.050 ;
        RECT 995.400 906.600 996.600 907.950 ;
        RECT 970.950 905.400 996.600 906.600 ;
        RECT 1009.950 906.600 1012.050 907.050 ;
        RECT 1018.950 906.600 1021.050 907.050 ;
        RECT 1024.950 906.600 1027.050 907.050 ;
        RECT 1009.950 905.400 1027.050 906.600 ;
        RECT 970.950 904.950 973.050 905.400 ;
        RECT 1009.950 904.950 1012.050 905.400 ;
        RECT 1018.950 904.950 1021.050 905.400 ;
        RECT 1024.950 904.950 1027.050 905.400 ;
        RECT 256.950 903.600 259.050 904.050 ;
        RECT 322.950 903.600 325.050 904.050 ;
        RECT 256.950 902.400 325.050 903.600 ;
        RECT 256.950 901.950 259.050 902.400 ;
        RECT 322.950 901.950 325.050 902.400 ;
        RECT 388.950 903.600 391.050 904.050 ;
        RECT 433.950 903.600 436.050 904.050 ;
        RECT 388.950 902.400 436.050 903.600 ;
        RECT 388.950 901.950 391.050 902.400 ;
        RECT 433.950 901.950 436.050 902.400 ;
        RECT 451.950 903.600 454.050 904.050 ;
        RECT 460.950 903.600 463.050 904.050 ;
        RECT 493.950 903.600 496.050 904.050 ;
        RECT 451.950 902.400 496.050 903.600 ;
        RECT 451.950 901.950 454.050 902.400 ;
        RECT 460.950 901.950 463.050 902.400 ;
        RECT 493.950 901.950 496.050 902.400 ;
        RECT 547.950 903.600 550.050 904.050 ;
        RECT 595.950 903.600 598.050 904.050 ;
        RECT 547.950 902.400 598.050 903.600 ;
        RECT 547.950 901.950 550.050 902.400 ;
        RECT 595.950 901.950 598.050 902.400 ;
        RECT 667.950 903.600 670.050 904.050 ;
        RECT 676.950 903.600 679.050 904.050 ;
        RECT 730.950 903.600 733.050 903.900 ;
        RECT 667.950 902.400 733.050 903.600 ;
        RECT 667.950 901.950 670.050 902.400 ;
        RECT 676.950 901.950 679.050 902.400 ;
        RECT 730.950 901.800 733.050 902.400 ;
        RECT 841.950 903.600 844.050 904.050 ;
        RECT 877.950 903.600 880.050 904.050 ;
        RECT 841.950 902.400 880.050 903.600 ;
        RECT 841.950 901.950 844.050 902.400 ;
        RECT 877.950 901.950 880.050 902.400 ;
        RECT 922.950 903.600 925.050 904.050 ;
        RECT 964.950 903.600 967.050 904.050 ;
        RECT 922.950 902.400 967.050 903.600 ;
        RECT 922.950 901.950 925.050 902.400 ;
        RECT 964.950 901.950 967.050 902.400 ;
        RECT 133.950 900.600 136.050 901.050 ;
        RECT 157.800 900.600 159.900 901.050 ;
        RECT 133.950 899.400 159.900 900.600 ;
        RECT 133.950 898.950 136.050 899.400 ;
        RECT 157.800 898.950 159.900 899.400 ;
        RECT 160.950 900.600 163.050 901.050 ;
        RECT 241.950 900.600 244.050 901.050 ;
        RECT 160.950 899.400 244.050 900.600 ;
        RECT 160.950 898.950 163.050 899.400 ;
        RECT 241.950 898.950 244.050 899.400 ;
        RECT 394.950 900.600 397.050 901.050 ;
        RECT 421.950 900.600 424.050 901.050 ;
        RECT 394.950 899.400 424.050 900.600 ;
        RECT 394.950 898.950 397.050 899.400 ;
        RECT 421.950 898.950 424.050 899.400 ;
        RECT 607.950 900.600 610.050 901.050 ;
        RECT 619.950 900.600 622.050 901.050 ;
        RECT 607.950 899.400 622.050 900.600 ;
        RECT 607.950 898.950 610.050 899.400 ;
        RECT 619.950 898.950 622.050 899.400 ;
        RECT 703.950 900.600 706.050 901.050 ;
        RECT 727.800 900.600 729.900 901.050 ;
        RECT 703.950 899.400 729.900 900.600 ;
        RECT 731.400 900.600 732.600 901.800 ;
        RECT 835.950 900.600 838.050 901.050 ;
        RECT 731.400 899.400 838.050 900.600 ;
        RECT 703.950 898.950 706.050 899.400 ;
        RECT 727.800 898.950 729.900 899.400 ;
        RECT 835.950 898.950 838.050 899.400 ;
        RECT 892.950 900.600 895.050 901.050 ;
        RECT 919.950 900.600 922.050 901.050 ;
        RECT 892.950 899.400 922.050 900.600 ;
        RECT 892.950 898.950 895.050 899.400 ;
        RECT 919.950 898.950 922.050 899.400 ;
        RECT 79.950 897.600 82.050 898.050 ;
        RECT 136.950 897.600 139.050 898.050 ;
        RECT 79.950 896.400 139.050 897.600 ;
        RECT 79.950 895.950 82.050 896.400 ;
        RECT 136.950 895.950 139.050 896.400 ;
        RECT 235.950 897.600 238.050 898.050 ;
        RECT 256.950 897.600 259.050 898.050 ;
        RECT 235.950 896.400 259.050 897.600 ;
        RECT 235.950 895.950 238.050 896.400 ;
        RECT 256.950 895.950 259.050 896.400 ;
        RECT 466.950 897.600 469.050 898.050 ;
        RECT 526.950 897.600 529.050 898.050 ;
        RECT 466.950 896.400 529.050 897.600 ;
        RECT 466.950 895.950 469.050 896.400 ;
        RECT 526.950 895.950 529.050 896.400 ;
        RECT 538.950 897.600 541.050 898.050 ;
        RECT 553.950 897.600 556.050 898.050 ;
        RECT 538.950 896.400 556.050 897.600 ;
        RECT 538.950 895.950 541.050 896.400 ;
        RECT 553.950 895.950 556.050 896.400 ;
        RECT 625.950 897.600 628.050 898.050 ;
        RECT 673.950 897.600 676.050 898.050 ;
        RECT 625.950 896.400 676.050 897.600 ;
        RECT 625.950 895.950 628.050 896.400 ;
        RECT 673.950 895.950 676.050 896.400 ;
        RECT 679.950 897.600 682.050 898.050 ;
        RECT 700.950 897.600 703.050 898.050 ;
        RECT 679.950 896.400 703.050 897.600 ;
        RECT 679.950 895.950 682.050 896.400 ;
        RECT 700.950 895.950 703.050 896.400 ;
        RECT 859.950 897.600 862.050 898.050 ;
        RECT 880.950 897.600 883.050 898.050 ;
        RECT 859.950 896.400 883.050 897.600 ;
        RECT 859.950 895.950 862.050 896.400 ;
        RECT 880.950 895.950 883.050 896.400 ;
        RECT 928.950 897.600 931.050 898.050 ;
        RECT 1003.950 897.600 1006.050 898.050 ;
        RECT 928.950 896.400 1006.050 897.600 ;
        RECT 928.950 895.950 931.050 896.400 ;
        RECT 1003.950 895.950 1006.050 896.400 ;
        RECT 127.950 894.600 130.050 895.050 ;
        RECT 160.950 894.600 163.050 895.050 ;
        RECT 127.950 893.400 163.050 894.600 ;
        RECT 127.950 892.950 130.050 893.400 ;
        RECT 160.950 892.950 163.050 893.400 ;
        RECT 220.950 894.600 223.050 895.050 ;
        RECT 298.950 894.600 301.050 895.050 ;
        RECT 337.950 894.600 340.050 895.050 ;
        RECT 220.950 893.400 340.050 894.600 ;
        RECT 220.950 892.950 223.050 893.400 ;
        RECT 298.950 892.950 301.050 893.400 ;
        RECT 337.950 892.950 340.050 893.400 ;
        RECT 751.950 894.600 754.050 895.050 ;
        RECT 793.950 894.600 796.050 895.050 ;
        RECT 751.950 893.400 796.050 894.600 ;
        RECT 751.950 892.950 754.050 893.400 ;
        RECT 793.950 892.950 796.050 893.400 ;
        RECT 838.950 894.600 841.050 895.050 ;
        RECT 847.950 894.600 850.050 895.050 ;
        RECT 838.950 893.400 850.050 894.600 ;
        RECT 838.950 892.950 841.050 893.400 ;
        RECT 847.950 892.950 850.050 893.400 ;
        RECT 907.950 894.600 910.050 895.050 ;
        RECT 964.950 894.600 967.050 895.050 ;
        RECT 907.950 893.400 967.050 894.600 ;
        RECT 907.950 892.950 910.050 893.400 ;
        RECT 964.950 892.950 967.050 893.400 ;
        RECT 250.950 891.600 253.050 892.050 ;
        RECT 385.950 891.600 388.050 892.050 ;
        RECT 412.950 891.600 415.050 892.050 ;
        RECT 250.950 890.400 357.600 891.600 ;
        RECT 250.950 889.950 253.050 890.400 ;
        RECT 356.400 888.600 357.600 890.400 ;
        RECT 385.950 890.400 415.050 891.600 ;
        RECT 385.950 889.950 388.050 890.400 ;
        RECT 412.950 889.950 415.050 890.400 ;
        RECT 508.950 889.950 511.050 892.050 ;
        RECT 598.950 891.600 601.050 892.050 ;
        RECT 637.950 891.600 640.050 892.050 ;
        RECT 598.950 890.400 640.050 891.600 ;
        RECT 598.950 889.950 601.050 890.400 ;
        RECT 637.950 889.950 640.050 890.400 ;
        RECT 643.950 891.600 646.050 892.050 ;
        RECT 694.950 891.600 697.050 892.050 ;
        RECT 706.950 891.600 709.050 892.050 ;
        RECT 643.950 890.400 654.600 891.600 ;
        RECT 643.950 889.950 646.050 890.400 ;
        RECT 361.950 888.600 364.050 889.050 ;
        RECT 356.400 887.400 364.050 888.600 ;
        RECT 361.950 886.950 364.050 887.400 ;
        RECT 22.950 885.750 25.050 886.200 ;
        RECT 37.950 885.750 40.050 886.200 ;
        RECT 22.950 884.550 40.050 885.750 ;
        RECT 22.950 884.100 25.050 884.550 ;
        RECT 37.950 884.100 40.050 884.550 ;
        RECT 115.950 885.600 118.050 886.200 ;
        RECT 139.950 885.600 142.050 886.200 ;
        RECT 115.950 884.400 142.050 885.600 ;
        RECT 115.950 884.100 118.050 884.400 ;
        RECT 139.950 884.100 142.050 884.400 ;
        RECT 241.950 885.750 244.050 886.200 ;
        RECT 250.950 885.750 253.050 886.200 ;
        RECT 241.950 884.550 253.050 885.750 ;
        RECT 241.950 884.100 244.050 884.550 ;
        RECT 250.950 884.100 253.050 884.550 ;
        RECT 265.950 885.600 268.050 886.050 ;
        RECT 283.950 885.600 286.050 886.200 ;
        RECT 265.950 884.400 286.050 885.600 ;
        RECT 265.950 883.950 268.050 884.400 ;
        RECT 283.950 884.100 286.050 884.400 ;
        RECT 304.950 885.750 307.050 886.200 ;
        RECT 313.800 885.750 315.900 886.200 ;
        RECT 304.950 884.550 315.900 885.750 ;
        RECT 304.950 884.100 307.050 884.550 ;
        RECT 313.800 884.100 315.900 884.550 ;
        RECT 316.950 885.750 319.050 886.200 ;
        RECT 325.950 885.750 328.050 886.200 ;
        RECT 316.950 884.550 328.050 885.750 ;
        RECT 355.950 885.600 358.050 886.200 ;
        RECT 316.950 884.100 319.050 884.550 ;
        RECT 325.950 884.100 328.050 884.550 ;
        RECT 329.400 884.400 358.050 885.600 ;
        RECT 88.950 882.600 91.050 883.200 ;
        RECT 319.950 882.600 322.050 883.050 ;
        RECT 329.400 882.600 330.600 884.400 ;
        RECT 355.950 884.100 358.050 884.400 ;
        RECT 367.950 885.600 370.050 886.050 ;
        RECT 379.950 885.600 382.050 886.200 ;
        RECT 367.950 884.400 382.050 885.600 ;
        RECT 367.950 883.950 370.050 884.400 ;
        RECT 379.950 884.100 382.050 884.400 ;
        RECT 400.950 885.750 403.050 886.200 ;
        RECT 406.950 885.750 409.050 886.200 ;
        RECT 400.950 884.550 409.050 885.750 ;
        RECT 442.950 885.600 445.050 886.050 ;
        RECT 400.950 884.100 403.050 884.550 ;
        RECT 406.950 884.100 409.050 884.550 ;
        RECT 410.400 884.400 445.050 885.600 ;
        RECT 410.400 882.600 411.600 884.400 ;
        RECT 442.950 883.950 445.050 884.400 ;
        RECT 481.950 885.600 484.050 886.200 ;
        RECT 502.950 885.600 505.050 886.200 ;
        RECT 509.400 886.050 510.600 889.950 ;
        RECT 514.950 888.600 517.050 889.050 ;
        RECT 529.950 888.600 532.050 889.050 ;
        RECT 514.950 887.400 532.050 888.600 ;
        RECT 514.950 886.950 517.050 887.400 ;
        RECT 529.950 886.950 532.050 887.400 ;
        RECT 481.950 884.400 507.600 885.600 ;
        RECT 509.400 884.400 514.050 886.050 ;
        RECT 481.950 884.100 484.050 884.400 ;
        RECT 502.950 884.100 505.050 884.400 ;
        RECT 88.950 881.400 114.600 882.600 ;
        RECT 88.950 881.100 91.050 881.400 ;
        RECT 100.950 879.600 103.050 880.050 ;
        RECT 109.950 879.600 112.050 879.900 ;
        RECT 100.950 878.400 112.050 879.600 ;
        RECT 113.400 879.600 114.600 881.400 ;
        RECT 319.950 881.400 330.600 882.600 ;
        RECT 392.400 881.400 411.600 882.600 ;
        RECT 506.400 882.600 507.600 884.400 ;
        RECT 510.000 883.950 514.050 884.400 ;
        RECT 517.950 885.750 520.050 886.200 ;
        RECT 523.950 885.750 526.050 886.200 ;
        RECT 517.950 884.550 526.050 885.750 ;
        RECT 517.950 884.100 520.050 884.550 ;
        RECT 523.950 884.100 526.050 884.550 ;
        RECT 550.950 885.600 553.050 886.200 ;
        RECT 577.950 885.600 580.050 886.200 ;
        RECT 550.950 884.400 580.050 885.600 ;
        RECT 550.950 884.100 553.050 884.400 ;
        RECT 577.950 884.100 580.050 884.400 ;
        RECT 613.950 885.600 616.050 886.050 ;
        RECT 625.950 885.600 628.050 886.200 ;
        RECT 613.950 884.400 628.050 885.600 ;
        RECT 613.950 883.950 616.050 884.400 ;
        RECT 625.950 884.100 628.050 884.400 ;
        RECT 649.950 884.100 652.050 886.200 ;
        RECT 506.400 881.400 528.600 882.600 ;
        RECT 319.950 880.950 322.050 881.400 ;
        RECT 121.950 879.600 124.050 880.050 ;
        RECT 160.950 879.600 163.050 879.900 ;
        RECT 113.400 878.400 163.050 879.600 ;
        RECT 100.950 877.950 103.050 878.400 ;
        RECT 109.950 877.800 112.050 878.400 ;
        RECT 121.950 877.950 124.050 878.400 ;
        RECT 160.950 877.800 163.050 878.400 ;
        RECT 241.950 879.600 244.050 880.050 ;
        RECT 247.950 879.600 250.050 880.050 ;
        RECT 241.950 878.400 250.050 879.600 ;
        RECT 241.950 877.950 244.050 878.400 ;
        RECT 247.950 877.950 250.050 878.400 ;
        RECT 259.950 879.450 262.050 879.900 ;
        RECT 265.950 879.450 268.050 879.900 ;
        RECT 259.950 878.250 268.050 879.450 ;
        RECT 259.950 877.800 262.050 878.250 ;
        RECT 265.950 877.800 268.050 878.250 ;
        RECT 295.950 879.600 298.050 880.050 ;
        RECT 301.950 879.600 304.050 880.050 ;
        RECT 295.950 878.400 304.050 879.600 ;
        RECT 295.950 877.950 298.050 878.400 ;
        RECT 301.950 877.950 304.050 878.400 ;
        RECT 307.950 879.600 310.050 879.900 ;
        RECT 316.950 879.600 319.050 880.050 ;
        RECT 307.950 878.400 319.050 879.600 ;
        RECT 307.950 877.800 310.050 878.400 ;
        RECT 316.950 877.950 319.050 878.400 ;
        RECT 358.950 879.450 361.050 879.900 ;
        RECT 367.950 879.450 370.050 879.900 ;
        RECT 358.950 878.250 370.050 879.450 ;
        RECT 358.950 877.800 361.050 878.250 ;
        RECT 367.950 877.800 370.050 878.250 ;
        RECT 388.950 879.600 391.050 879.900 ;
        RECT 392.400 879.600 393.600 881.400 ;
        RECT 388.950 878.400 393.600 879.600 ;
        RECT 415.950 879.450 418.050 879.900 ;
        RECT 421.950 879.450 424.050 879.900 ;
        RECT 388.950 877.800 391.050 878.400 ;
        RECT 415.950 878.250 424.050 879.450 ;
        RECT 415.950 877.800 418.050 878.250 ;
        RECT 421.950 877.800 424.050 878.250 ;
        RECT 436.950 879.450 439.050 879.900 ;
        RECT 445.950 879.450 448.050 879.900 ;
        RECT 436.950 878.250 448.050 879.450 ;
        RECT 436.950 877.800 439.050 878.250 ;
        RECT 445.950 877.800 448.050 878.250 ;
        RECT 457.950 879.600 460.050 879.900 ;
        RECT 478.950 879.600 481.050 879.900 ;
        RECT 457.950 878.400 481.050 879.600 ;
        RECT 457.950 877.800 460.050 878.400 ;
        RECT 478.950 877.800 481.050 878.400 ;
        RECT 505.950 879.600 508.050 879.900 ;
        RECT 511.950 879.600 514.050 880.050 ;
        RECT 505.950 878.400 514.050 879.600 ;
        RECT 527.400 879.600 528.600 881.400 ;
        RECT 650.400 880.050 651.600 884.100 ;
        RECT 547.950 879.600 550.050 879.900 ;
        RECT 527.400 878.400 550.050 879.600 ;
        RECT 505.950 877.800 508.050 878.400 ;
        RECT 511.950 877.950 514.050 878.400 ;
        RECT 547.950 877.800 550.050 878.400 ;
        RECT 592.950 879.600 595.050 880.050 ;
        RECT 607.950 879.600 610.050 879.900 ;
        RECT 628.950 879.600 631.050 879.900 ;
        RECT 592.950 878.400 631.050 879.600 ;
        RECT 592.950 877.950 595.050 878.400 ;
        RECT 607.950 877.800 610.050 878.400 ;
        RECT 628.950 877.800 631.050 878.400 ;
        RECT 646.950 878.400 651.600 880.050 ;
        RECT 653.400 879.900 654.600 890.400 ;
        RECT 694.950 890.400 709.050 891.600 ;
        RECT 694.950 889.950 697.050 890.400 ;
        RECT 706.950 889.950 709.050 890.400 ;
        RECT 778.950 891.600 781.050 892.050 ;
        RECT 787.950 891.600 790.050 892.050 ;
        RECT 778.950 890.400 790.050 891.600 ;
        RECT 778.950 889.950 781.050 890.400 ;
        RECT 787.950 889.950 790.050 890.400 ;
        RECT 940.950 891.600 943.050 892.050 ;
        RECT 949.950 891.600 952.050 892.050 ;
        RECT 985.950 891.600 988.050 892.050 ;
        RECT 940.950 890.400 988.050 891.600 ;
        RECT 940.950 889.950 943.050 890.400 ;
        RECT 949.950 889.950 952.050 890.400 ;
        RECT 985.950 889.950 988.050 890.400 ;
        RECT 685.950 888.600 688.050 889.050 ;
        RECT 691.950 888.600 694.050 889.050 ;
        RECT 685.950 887.400 694.050 888.600 ;
        RECT 685.950 886.950 688.050 887.400 ;
        RECT 691.950 886.950 694.050 887.400 ;
        RECT 751.950 888.600 754.050 889.050 ;
        RECT 796.950 888.600 799.050 889.050 ;
        RECT 751.950 887.400 799.050 888.600 ;
        RECT 751.950 886.950 754.050 887.400 ;
        RECT 796.950 886.950 799.050 887.400 ;
        RECT 835.950 888.600 838.050 889.200 ;
        RECT 907.950 888.600 910.050 889.050 ;
        RECT 835.950 887.400 910.050 888.600 ;
        RECT 835.950 887.100 838.050 887.400 ;
        RECT 907.950 886.950 910.050 887.400 ;
        RECT 661.950 885.750 664.050 886.200 ;
        RECT 670.950 885.750 673.050 886.200 ;
        RECT 661.950 884.550 673.050 885.750 ;
        RECT 661.950 884.100 664.050 884.550 ;
        RECT 670.950 884.100 673.050 884.550 ;
        RECT 703.950 884.100 706.050 886.200 ;
        RECT 724.950 885.600 727.050 886.050 ;
        RECT 742.950 885.600 745.050 886.050 ;
        RECT 724.950 884.400 745.050 885.600 ;
        RECT 704.400 882.600 705.600 884.100 ;
        RECT 724.950 883.950 727.050 884.400 ;
        RECT 742.950 883.950 745.050 884.400 ;
        RECT 757.950 885.750 760.050 886.200 ;
        RECT 766.950 885.750 769.050 886.200 ;
        RECT 757.950 884.550 769.050 885.750 ;
        RECT 781.950 885.600 784.050 886.200 ;
        RECT 757.950 884.100 760.050 884.550 ;
        RECT 766.950 884.100 769.050 884.550 ;
        RECT 770.400 884.400 784.050 885.600 ;
        RECT 770.400 882.600 771.600 884.400 ;
        RECT 781.950 884.100 784.050 884.400 ;
        RECT 802.950 885.600 805.050 886.050 ;
        RECT 808.950 885.600 811.050 886.200 ;
        RECT 835.950 885.600 838.050 886.050 ;
        RECT 802.950 884.400 838.050 885.600 ;
        RECT 802.950 883.950 805.050 884.400 ;
        RECT 808.950 884.100 811.050 884.400 ;
        RECT 809.400 882.600 810.600 884.100 ;
        RECT 835.950 883.950 838.050 884.400 ;
        RECT 877.950 885.750 880.050 886.200 ;
        RECT 886.950 885.750 889.050 886.200 ;
        RECT 877.950 884.550 889.050 885.750 ;
        RECT 877.950 884.100 880.050 884.550 ;
        RECT 886.950 884.100 889.050 884.550 ;
        RECT 910.950 884.100 913.050 886.200 ;
        RECT 916.950 885.600 919.050 886.200 ;
        RECT 925.950 885.600 928.050 886.050 ;
        RECT 916.950 884.400 928.050 885.600 ;
        RECT 916.950 884.100 919.050 884.400 ;
        RECT 898.950 882.600 901.050 883.050 ;
        RECT 701.400 882.000 705.600 882.600 ;
        RECT 700.950 881.400 705.600 882.000 ;
        RECT 758.400 881.400 771.600 882.600 ;
        RECT 788.400 881.400 810.600 882.600 ;
        RECT 890.400 881.400 901.050 882.600 ;
        RECT 646.950 877.950 651.000 878.400 ;
        RECT 652.950 877.800 655.050 879.900 ;
        RECT 658.950 879.450 661.050 879.900 ;
        RECT 667.950 879.450 670.050 879.900 ;
        RECT 658.950 878.250 670.050 879.450 ;
        RECT 658.950 877.800 661.050 878.250 ;
        RECT 667.950 877.800 670.050 878.250 ;
        RECT 673.950 879.600 676.050 880.050 ;
        RECT 682.950 879.600 685.050 879.900 ;
        RECT 673.950 878.400 685.050 879.600 ;
        RECT 673.950 877.950 676.050 878.400 ;
        RECT 682.950 877.800 685.050 878.400 ;
        RECT 700.950 877.950 703.050 881.400 ;
        RECT 706.950 879.600 709.050 879.900 ;
        RECT 712.950 879.600 715.050 880.050 ;
        RECT 706.950 878.400 715.050 879.600 ;
        RECT 706.950 877.800 709.050 878.400 ;
        RECT 712.950 877.950 715.050 878.400 ;
        RECT 754.950 879.600 757.050 879.900 ;
        RECT 758.400 879.600 759.600 881.400 ;
        RECT 754.950 878.400 759.600 879.600 ;
        RECT 784.950 879.600 787.050 879.900 ;
        RECT 788.400 879.600 789.600 881.400 ;
        RECT 784.950 878.400 789.600 879.600 ;
        RECT 799.950 879.600 802.050 880.050 ;
        RECT 890.400 879.600 891.600 881.400 ;
        RECT 898.950 880.950 901.050 881.400 ;
        RECT 799.950 878.400 891.600 879.600 ;
        RECT 911.400 879.600 912.600 884.100 ;
        RECT 925.950 883.950 928.050 884.400 ;
        RECT 931.800 885.000 933.900 886.050 ;
        RECT 934.950 885.600 937.050 886.200 ;
        RECT 949.950 885.600 952.050 886.050 ;
        RECT 931.800 883.950 934.050 885.000 ;
        RECT 934.950 884.400 952.050 885.600 ;
        RECT 934.950 884.100 937.050 884.400 ;
        RECT 949.950 883.950 952.050 884.400 ;
        RECT 970.950 885.600 973.050 886.200 ;
        RECT 976.950 885.600 979.050 886.050 ;
        RECT 970.950 884.400 979.050 885.600 ;
        RECT 970.950 884.100 973.050 884.400 ;
        RECT 976.950 883.950 979.050 884.400 ;
        RECT 994.950 885.750 997.050 886.200 ;
        RECT 1003.950 885.750 1006.050 886.200 ;
        RECT 994.950 884.550 1006.050 885.750 ;
        RECT 994.950 884.100 997.050 884.550 ;
        RECT 1003.950 884.100 1006.050 884.550 ;
        RECT 931.950 882.600 934.050 883.950 ;
        RECT 931.950 882.000 945.600 882.600 ;
        RECT 932.400 881.400 945.600 882.000 ;
        RECT 919.950 879.600 922.050 880.050 ;
        RECT 944.400 879.900 945.600 881.400 ;
        RECT 911.400 878.400 922.050 879.600 ;
        RECT 754.950 877.800 757.050 878.400 ;
        RECT 784.950 877.800 787.050 878.400 ;
        RECT 799.950 877.950 802.050 878.400 ;
        RECT 919.950 877.950 922.050 878.400 ;
        RECT 928.950 879.450 931.050 879.900 ;
        RECT 937.950 879.450 940.050 879.900 ;
        RECT 928.950 878.250 940.050 879.450 ;
        RECT 928.950 877.800 931.050 878.250 ;
        RECT 937.950 877.800 940.050 878.250 ;
        RECT 943.950 877.800 946.050 879.900 ;
        RECT 967.950 879.450 970.050 879.900 ;
        RECT 982.950 879.450 985.050 879.900 ;
        RECT 967.950 878.250 985.050 879.450 ;
        RECT 967.950 877.800 970.050 878.250 ;
        RECT 982.950 877.800 985.050 878.250 ;
        RECT 1003.950 879.600 1006.050 880.050 ;
        RECT 1015.950 879.600 1018.050 879.900 ;
        RECT 1003.950 878.400 1018.050 879.600 ;
        RECT 1003.950 877.950 1006.050 878.400 ;
        RECT 1015.950 877.800 1018.050 878.400 ;
        RECT 16.950 876.450 19.050 876.900 ;
        RECT 28.950 876.450 31.050 876.900 ;
        RECT 697.950 876.600 700.050 877.050 ;
        RECT 16.950 875.250 31.050 876.450 ;
        RECT 16.950 874.800 19.050 875.250 ;
        RECT 28.950 874.800 31.050 875.250 ;
        RECT 635.400 875.400 700.050 876.600 ;
        RECT 148.950 873.600 151.050 874.050 ;
        RECT 163.950 873.600 166.050 874.050 ;
        RECT 148.950 872.400 166.050 873.600 ;
        RECT 148.950 871.950 151.050 872.400 ;
        RECT 163.950 871.950 166.050 872.400 ;
        RECT 214.950 873.600 217.050 874.050 ;
        RECT 319.950 873.600 322.050 874.050 ;
        RECT 214.950 872.400 322.050 873.600 ;
        RECT 214.950 871.950 217.050 872.400 ;
        RECT 319.950 871.950 322.050 872.400 ;
        RECT 325.950 873.600 328.050 874.050 ;
        RECT 352.950 873.600 355.050 874.050 ;
        RECT 325.950 872.400 355.050 873.600 ;
        RECT 325.950 871.950 328.050 872.400 ;
        RECT 352.950 871.950 355.050 872.400 ;
        RECT 376.950 873.600 379.050 874.050 ;
        RECT 394.950 873.600 397.050 874.050 ;
        RECT 376.950 872.400 397.050 873.600 ;
        RECT 376.950 871.950 379.050 872.400 ;
        RECT 394.950 871.950 397.050 872.400 ;
        RECT 424.950 873.600 427.050 874.050 ;
        RECT 469.950 873.600 472.050 874.050 ;
        RECT 604.950 873.600 607.050 874.050 ;
        RECT 635.400 873.600 636.600 875.400 ;
        RECT 697.950 874.950 700.050 875.400 ;
        RECT 703.950 876.600 706.050 877.050 ;
        RECT 745.950 876.600 748.050 877.050 ;
        RECT 703.950 875.400 748.050 876.600 ;
        RECT 703.950 874.950 706.050 875.400 ;
        RECT 745.950 874.950 748.050 875.400 ;
        RECT 826.950 876.600 829.050 877.050 ;
        RECT 895.950 876.600 898.050 877.050 ;
        RECT 826.950 875.400 898.050 876.600 ;
        RECT 826.950 874.950 829.050 875.400 ;
        RECT 895.950 874.950 898.050 875.400 ;
        RECT 901.950 876.600 904.050 877.050 ;
        RECT 913.950 876.600 916.050 877.050 ;
        RECT 952.950 876.600 955.050 877.050 ;
        RECT 901.950 875.400 955.050 876.600 ;
        RECT 983.400 876.600 984.600 877.800 ;
        RECT 1021.950 876.600 1024.050 877.050 ;
        RECT 983.400 875.400 1024.050 876.600 ;
        RECT 901.950 874.950 904.050 875.400 ;
        RECT 913.950 874.950 916.050 875.400 ;
        RECT 952.950 874.950 955.050 875.400 ;
        RECT 1021.950 874.950 1024.050 875.400 ;
        RECT 646.800 873.600 648.900 874.050 ;
        RECT 424.950 872.400 636.600 873.600 ;
        RECT 638.400 872.400 648.900 873.600 ;
        RECT 424.950 871.950 427.050 872.400 ;
        RECT 469.950 871.950 472.050 872.400 ;
        RECT 604.950 871.950 607.050 872.400 ;
        RECT 355.950 870.600 358.050 871.050 ;
        RECT 397.950 870.600 400.050 871.050 ;
        RECT 409.950 870.600 412.050 871.050 ;
        RECT 355.950 869.400 412.050 870.600 ;
        RECT 355.950 868.950 358.050 869.400 ;
        RECT 397.950 868.950 400.050 869.400 ;
        RECT 409.950 868.950 412.050 869.400 ;
        RECT 493.950 870.600 496.050 871.050 ;
        RECT 574.950 870.600 577.050 871.050 ;
        RECT 493.950 869.400 577.050 870.600 ;
        RECT 493.950 868.950 496.050 869.400 ;
        RECT 574.950 868.950 577.050 869.400 ;
        RECT 613.950 870.600 616.050 871.050 ;
        RECT 638.400 870.600 639.600 872.400 ;
        RECT 646.800 871.950 648.900 872.400 ;
        RECT 649.950 873.600 652.050 874.050 ;
        RECT 688.950 873.600 691.050 874.050 ;
        RECT 649.950 872.400 691.050 873.600 ;
        RECT 649.950 871.950 652.050 872.400 ;
        RECT 688.950 871.950 691.050 872.400 ;
        RECT 772.950 873.600 775.050 874.050 ;
        RECT 787.950 873.600 790.050 874.050 ;
        RECT 772.950 872.400 790.050 873.600 ;
        RECT 772.950 871.950 775.050 872.400 ;
        RECT 787.950 871.950 790.050 872.400 ;
        RECT 805.950 873.600 808.050 874.050 ;
        RECT 838.950 873.600 841.050 874.050 ;
        RECT 805.950 872.400 841.050 873.600 ;
        RECT 805.950 871.950 808.050 872.400 ;
        RECT 838.950 871.950 841.050 872.400 ;
        RECT 856.950 873.600 859.050 874.050 ;
        RECT 880.950 873.600 883.050 874.050 ;
        RECT 856.950 872.400 883.050 873.600 ;
        RECT 856.950 871.950 859.050 872.400 ;
        RECT 880.950 871.950 883.050 872.400 ;
        RECT 898.950 873.600 901.050 874.050 ;
        RECT 928.950 873.600 931.050 874.050 ;
        RECT 898.950 872.400 931.050 873.600 ;
        RECT 898.950 871.950 901.050 872.400 ;
        RECT 928.950 871.950 931.050 872.400 ;
        RECT 985.950 873.600 988.050 874.050 ;
        RECT 997.950 873.600 1000.050 874.050 ;
        RECT 985.950 872.400 1000.050 873.600 ;
        RECT 985.950 871.950 988.050 872.400 ;
        RECT 997.950 871.950 1000.050 872.400 ;
        RECT 613.950 869.400 639.600 870.600 ;
        RECT 640.950 870.600 643.050 871.050 ;
        RECT 712.950 870.600 715.050 871.050 ;
        RECT 640.950 869.400 715.050 870.600 ;
        RECT 613.950 868.950 616.050 869.400 ;
        RECT 640.950 868.950 643.050 869.400 ;
        RECT 712.950 868.950 715.050 869.400 ;
        RECT 727.950 870.600 730.050 871.050 ;
        RECT 754.950 870.600 757.050 871.050 ;
        RECT 727.950 869.400 757.050 870.600 ;
        RECT 727.950 868.950 730.050 869.400 ;
        RECT 754.950 868.950 757.050 869.400 ;
        RECT 760.950 870.600 763.050 871.050 ;
        RECT 799.950 870.600 802.050 871.050 ;
        RECT 760.950 869.400 802.050 870.600 ;
        RECT 760.950 868.950 763.050 869.400 ;
        RECT 799.950 868.950 802.050 869.400 ;
        RECT 811.950 870.600 814.050 871.050 ;
        RECT 832.950 870.600 835.050 871.050 ;
        RECT 811.950 869.400 835.050 870.600 ;
        RECT 811.950 868.950 814.050 869.400 ;
        RECT 832.950 868.950 835.050 869.400 ;
        RECT 949.950 870.600 952.050 870.900 ;
        RECT 955.950 870.600 958.050 871.050 ;
        RECT 949.950 869.400 958.050 870.600 ;
        RECT 949.950 868.800 952.050 869.400 ;
        RECT 955.950 868.950 958.050 869.400 ;
        RECT 961.950 870.600 964.050 871.050 ;
        RECT 997.950 870.600 1000.050 870.900 ;
        RECT 961.950 869.400 1000.050 870.600 ;
        RECT 961.950 868.950 964.050 869.400 ;
        RECT 997.950 868.800 1000.050 869.400 ;
        RECT 52.950 867.600 55.050 868.050 ;
        RECT 100.950 867.600 103.050 868.050 ;
        RECT 154.950 867.600 157.050 868.050 ;
        RECT 52.950 866.400 157.050 867.600 ;
        RECT 52.950 865.950 55.050 866.400 ;
        RECT 100.950 865.950 103.050 866.400 ;
        RECT 154.950 865.950 157.050 866.400 ;
        RECT 163.950 867.600 166.050 868.050 ;
        RECT 196.950 867.600 199.050 868.050 ;
        RECT 343.950 867.600 346.050 868.050 ;
        RECT 163.950 866.400 346.050 867.600 ;
        RECT 163.950 865.950 166.050 866.400 ;
        RECT 196.950 865.950 199.050 866.400 ;
        RECT 343.950 865.950 346.050 866.400 ;
        RECT 394.950 867.600 397.050 868.050 ;
        RECT 451.950 867.600 454.050 868.050 ;
        RECT 394.950 866.400 454.050 867.600 ;
        RECT 394.950 865.950 397.050 866.400 ;
        RECT 451.950 865.950 454.050 866.400 ;
        RECT 484.950 867.600 487.050 868.050 ;
        RECT 622.950 867.600 625.050 868.050 ;
        RECT 484.950 866.400 625.050 867.600 ;
        RECT 484.950 865.950 487.050 866.400 ;
        RECT 622.950 865.950 625.050 866.400 ;
        RECT 679.950 867.600 682.050 868.050 ;
        RECT 700.950 867.600 703.050 868.050 ;
        RECT 679.950 866.400 703.050 867.600 ;
        RECT 679.950 865.950 682.050 866.400 ;
        RECT 700.950 865.950 703.050 866.400 ;
        RECT 739.950 867.600 742.050 868.050 ;
        RECT 751.950 867.600 754.050 868.050 ;
        RECT 739.950 866.400 754.050 867.600 ;
        RECT 739.950 865.950 742.050 866.400 ;
        RECT 751.950 865.950 754.050 866.400 ;
        RECT 769.950 867.600 772.050 868.050 ;
        RECT 778.950 867.600 781.050 868.050 ;
        RECT 793.800 867.600 795.900 868.050 ;
        RECT 769.950 866.400 795.900 867.600 ;
        RECT 769.950 865.950 772.050 866.400 ;
        RECT 778.950 865.950 781.050 866.400 ;
        RECT 793.800 865.950 795.900 866.400 ;
        RECT 796.950 867.600 799.050 868.050 ;
        RECT 862.950 867.600 865.050 868.050 ;
        RECT 877.950 867.600 880.050 868.050 ;
        RECT 796.950 866.400 880.050 867.600 ;
        RECT 796.950 865.950 799.050 866.400 ;
        RECT 862.950 865.950 865.050 866.400 ;
        RECT 877.950 865.950 880.050 866.400 ;
        RECT 886.950 867.600 889.050 868.050 ;
        RECT 943.950 867.600 946.050 868.050 ;
        RECT 886.950 866.400 946.050 867.600 ;
        RECT 886.950 865.950 889.050 866.400 ;
        RECT 943.950 865.950 946.050 866.400 ;
        RECT 292.950 864.600 295.050 865.050 ;
        RECT 355.950 864.600 358.050 865.050 ;
        RECT 292.950 863.400 358.050 864.600 ;
        RECT 292.950 862.950 295.050 863.400 ;
        RECT 355.950 862.950 358.050 863.400 ;
        RECT 547.950 864.600 550.050 865.050 ;
        RECT 631.950 864.600 634.050 865.050 ;
        RECT 547.950 863.400 634.050 864.600 ;
        RECT 547.950 862.950 550.050 863.400 ;
        RECT 631.950 862.950 634.050 863.400 ;
        RECT 637.950 864.600 640.050 865.050 ;
        RECT 799.950 864.600 802.050 865.050 ;
        RECT 844.950 864.600 847.050 865.050 ;
        RECT 637.950 863.400 771.600 864.600 ;
        RECT 637.950 862.950 640.050 863.400 ;
        RECT 223.950 861.600 226.050 862.050 ;
        RECT 280.950 861.600 283.050 862.050 ;
        RECT 223.950 860.400 283.050 861.600 ;
        RECT 223.950 859.950 226.050 860.400 ;
        RECT 280.950 859.950 283.050 860.400 ;
        RECT 373.950 861.600 376.050 862.050 ;
        RECT 385.950 861.600 388.050 862.050 ;
        RECT 430.950 861.600 433.050 862.050 ;
        RECT 373.950 860.400 433.050 861.600 ;
        RECT 373.950 859.950 376.050 860.400 ;
        RECT 385.950 859.950 388.050 860.400 ;
        RECT 430.950 859.950 433.050 860.400 ;
        RECT 436.950 861.600 439.050 862.050 ;
        RECT 535.950 861.600 538.050 862.050 ;
        RECT 436.950 860.400 538.050 861.600 ;
        RECT 436.950 859.950 439.050 860.400 ;
        RECT 535.950 859.950 538.050 860.400 ;
        RECT 574.950 861.600 577.050 862.050 ;
        RECT 670.950 861.600 673.050 862.050 ;
        RECT 574.950 860.400 673.050 861.600 ;
        RECT 574.950 859.950 577.050 860.400 ;
        RECT 670.950 859.950 673.050 860.400 ;
        RECT 691.950 861.600 694.050 862.050 ;
        RECT 703.950 861.600 706.050 862.050 ;
        RECT 691.950 860.400 706.050 861.600 ;
        RECT 691.950 859.950 694.050 860.400 ;
        RECT 703.950 859.950 706.050 860.400 ;
        RECT 733.950 861.600 736.050 862.050 ;
        RECT 754.950 861.600 757.050 862.050 ;
        RECT 766.950 861.600 769.050 862.050 ;
        RECT 733.950 860.400 769.050 861.600 ;
        RECT 770.400 861.600 771.600 863.400 ;
        RECT 799.950 863.400 847.050 864.600 ;
        RECT 799.950 862.950 802.050 863.400 ;
        RECT 844.950 862.950 847.050 863.400 ;
        RECT 919.950 864.600 922.050 865.050 ;
        RECT 970.950 864.600 973.050 865.050 ;
        RECT 919.950 863.400 973.050 864.600 ;
        RECT 919.950 862.950 922.050 863.400 ;
        RECT 970.950 862.950 973.050 863.400 ;
        RECT 865.950 861.600 868.050 862.050 ;
        RECT 770.400 860.400 868.050 861.600 ;
        RECT 733.950 859.950 736.050 860.400 ;
        RECT 754.950 859.950 757.050 860.400 ;
        RECT 766.950 859.950 769.050 860.400 ;
        RECT 865.950 859.950 868.050 860.400 ;
        RECT 928.950 861.600 931.050 862.050 ;
        RECT 1021.950 861.600 1024.050 862.050 ;
        RECT 928.950 860.400 1024.050 861.600 ;
        RECT 928.950 859.950 931.050 860.400 ;
        RECT 1021.950 859.950 1024.050 860.400 ;
        RECT 7.950 858.600 10.050 859.050 ;
        RECT 28.950 858.600 31.050 859.050 ;
        RECT 145.950 858.600 148.050 859.050 ;
        RECT 169.950 858.600 172.050 859.050 ;
        RECT 7.950 857.400 172.050 858.600 ;
        RECT 7.950 856.950 10.050 857.400 ;
        RECT 28.950 856.950 31.050 857.400 ;
        RECT 145.950 856.950 148.050 857.400 ;
        RECT 169.950 856.950 172.050 857.400 ;
        RECT 286.950 858.600 289.050 859.050 ;
        RECT 313.950 858.600 316.050 859.050 ;
        RECT 322.950 858.600 325.050 859.050 ;
        RECT 286.950 857.400 325.050 858.600 ;
        RECT 286.950 856.950 289.050 857.400 ;
        RECT 313.950 856.950 316.050 857.400 ;
        RECT 322.950 856.950 325.050 857.400 ;
        RECT 343.950 858.600 346.050 859.050 ;
        RECT 394.950 858.600 397.050 859.050 ;
        RECT 343.950 857.400 397.050 858.600 ;
        RECT 343.950 856.950 346.050 857.400 ;
        RECT 394.950 856.950 397.050 857.400 ;
        RECT 565.950 858.600 568.050 859.050 ;
        RECT 643.950 858.600 646.050 859.050 ;
        RECT 913.950 858.600 916.050 859.050 ;
        RECT 565.950 857.400 916.050 858.600 ;
        RECT 565.950 856.950 568.050 857.400 ;
        RECT 643.950 856.950 646.050 857.400 ;
        RECT 913.950 856.950 916.050 857.400 ;
        RECT 175.950 855.600 178.050 856.050 ;
        RECT 244.950 855.600 247.050 856.050 ;
        RECT 175.950 854.400 247.050 855.600 ;
        RECT 175.950 853.950 178.050 854.400 ;
        RECT 244.950 853.950 247.050 854.400 ;
        RECT 334.950 855.600 337.050 856.050 ;
        RECT 400.950 855.600 403.050 856.050 ;
        RECT 334.950 854.400 403.050 855.600 ;
        RECT 334.950 853.950 337.050 854.400 ;
        RECT 400.950 853.950 403.050 854.400 ;
        RECT 571.950 855.600 574.050 856.050 ;
        RECT 613.950 855.600 616.050 856.050 ;
        RECT 571.950 854.400 616.050 855.600 ;
        RECT 571.950 853.950 574.050 854.400 ;
        RECT 613.950 853.950 616.050 854.400 ;
        RECT 619.950 855.600 622.050 856.050 ;
        RECT 628.950 855.600 631.050 856.050 ;
        RECT 793.950 855.600 796.050 856.050 ;
        RECT 619.950 854.400 631.050 855.600 ;
        RECT 619.950 853.950 622.050 854.400 ;
        RECT 628.950 853.950 631.050 854.400 ;
        RECT 632.400 854.400 796.050 855.600 ;
        RECT 142.950 852.600 145.050 853.050 ;
        RECT 271.950 852.600 274.050 853.050 ;
        RECT 316.950 852.600 319.050 853.050 ;
        RECT 142.950 851.400 267.600 852.600 ;
        RECT 142.950 850.950 145.050 851.400 ;
        RECT 266.400 850.050 267.600 851.400 ;
        RECT 271.950 851.400 319.050 852.600 ;
        RECT 271.950 850.950 274.050 851.400 ;
        RECT 316.950 850.950 319.050 851.400 ;
        RECT 442.950 852.600 445.050 853.050 ;
        RECT 538.950 852.600 541.050 853.050 ;
        RECT 442.950 851.400 541.050 852.600 ;
        RECT 442.950 850.950 445.050 851.400 ;
        RECT 538.950 850.950 541.050 851.400 ;
        RECT 616.950 852.600 619.050 853.050 ;
        RECT 632.400 852.600 633.600 854.400 ;
        RECT 793.950 853.950 796.050 854.400 ;
        RECT 838.950 855.600 841.050 856.050 ;
        RECT 868.950 855.600 871.050 856.050 ;
        RECT 838.950 854.400 871.050 855.600 ;
        RECT 838.950 853.950 841.050 854.400 ;
        RECT 868.950 853.950 871.050 854.400 ;
        RECT 922.950 855.600 925.050 856.050 ;
        RECT 946.950 855.600 949.050 856.050 ;
        RECT 922.950 854.400 949.050 855.600 ;
        RECT 922.950 853.950 925.050 854.400 ;
        RECT 946.950 853.950 949.050 854.400 ;
        RECT 616.950 851.400 633.600 852.600 ;
        RECT 661.950 852.600 664.050 853.050 ;
        RECT 823.950 852.600 826.050 853.050 ;
        RECT 892.950 852.600 895.050 853.050 ;
        RECT 661.950 851.400 765.600 852.600 ;
        RECT 616.950 850.950 619.050 851.400 ;
        RECT 661.950 850.950 664.050 851.400 ;
        RECT 265.950 849.600 268.050 850.050 ;
        RECT 334.950 849.600 337.050 850.050 ;
        RECT 265.950 848.400 337.050 849.600 ;
        RECT 265.950 847.950 268.050 848.400 ;
        RECT 334.950 847.950 337.050 848.400 ;
        RECT 400.950 849.600 403.050 850.050 ;
        RECT 457.950 849.600 460.050 850.050 ;
        RECT 400.950 848.400 460.050 849.600 ;
        RECT 400.950 847.950 403.050 848.400 ;
        RECT 457.950 847.950 460.050 848.400 ;
        RECT 592.950 849.600 595.050 850.050 ;
        RECT 646.950 849.600 649.050 850.050 ;
        RECT 712.950 849.600 715.050 850.050 ;
        RECT 592.950 848.400 715.050 849.600 ;
        RECT 592.950 847.950 595.050 848.400 ;
        RECT 646.950 847.950 649.050 848.400 ;
        RECT 712.950 847.950 715.050 848.400 ;
        RECT 742.950 849.600 745.050 850.050 ;
        RECT 757.950 849.600 760.050 850.050 ;
        RECT 742.950 848.400 760.050 849.600 ;
        RECT 764.400 849.600 765.600 851.400 ;
        RECT 823.950 851.400 895.050 852.600 ;
        RECT 823.950 850.950 826.050 851.400 ;
        RECT 892.950 850.950 895.050 851.400 ;
        RECT 913.950 852.600 916.050 853.050 ;
        RECT 994.950 852.600 997.050 853.050 ;
        RECT 1006.950 852.600 1009.050 853.050 ;
        RECT 913.950 851.400 1009.050 852.600 ;
        RECT 913.950 850.950 916.050 851.400 ;
        RECT 994.950 850.950 997.050 851.400 ;
        RECT 1006.950 850.950 1009.050 851.400 ;
        RECT 826.950 849.600 829.050 850.050 ;
        RECT 764.400 848.400 829.050 849.600 ;
        RECT 742.950 847.950 745.050 848.400 ;
        RECT 757.950 847.950 760.050 848.400 ;
        RECT 826.950 847.950 829.050 848.400 ;
        RECT 832.950 849.600 835.050 850.050 ;
        RECT 841.950 849.600 844.050 850.050 ;
        RECT 832.950 848.400 844.050 849.600 ;
        RECT 832.950 847.950 835.050 848.400 ;
        RECT 841.950 847.950 844.050 848.400 ;
        RECT 880.950 849.600 883.050 850.050 ;
        RECT 895.950 849.600 898.050 850.050 ;
        RECT 880.950 848.400 898.050 849.600 ;
        RECT 880.950 847.950 883.050 848.400 ;
        RECT 895.950 847.950 898.050 848.400 ;
        RECT 955.950 849.600 958.050 850.050 ;
        RECT 985.950 849.600 988.050 850.050 ;
        RECT 955.950 848.400 988.050 849.600 ;
        RECT 955.950 847.950 958.050 848.400 ;
        RECT 985.950 847.950 988.050 848.400 ;
        RECT 211.950 846.600 214.050 847.050 ;
        RECT 286.950 846.600 289.050 847.050 ;
        RECT 211.950 845.400 289.050 846.600 ;
        RECT 211.950 844.950 214.050 845.400 ;
        RECT 286.950 844.950 289.050 845.400 ;
        RECT 307.950 846.600 310.050 847.050 ;
        RECT 340.950 846.600 343.050 847.050 ;
        RECT 397.950 846.600 400.050 847.050 ;
        RECT 442.950 846.600 445.050 847.050 ;
        RECT 307.950 845.400 372.600 846.600 ;
        RECT 307.950 844.950 310.050 845.400 ;
        RECT 340.950 844.950 343.050 845.400 ;
        RECT 52.950 843.600 55.050 844.050 ;
        RECT 112.950 843.600 115.050 844.050 ;
        RECT 52.950 842.400 115.050 843.600 ;
        RECT 52.950 841.950 55.050 842.400 ;
        RECT 112.950 841.950 115.050 842.400 ;
        RECT 118.950 843.600 121.050 844.050 ;
        RECT 148.950 843.600 151.050 844.050 ;
        RECT 118.950 842.400 151.050 843.600 ;
        RECT 118.950 841.950 121.050 842.400 ;
        RECT 148.950 841.950 151.050 842.400 ;
        RECT 253.950 843.600 256.050 844.050 ;
        RECT 277.950 843.600 280.050 844.050 ;
        RECT 253.950 842.400 280.050 843.600 ;
        RECT 371.400 843.600 372.600 845.400 ;
        RECT 397.950 845.400 445.050 846.600 ;
        RECT 397.950 844.950 400.050 845.400 ;
        RECT 442.950 844.950 445.050 845.400 ;
        RECT 628.950 846.600 631.050 847.050 ;
        RECT 718.950 846.600 721.050 847.050 ;
        RECT 628.950 845.400 721.050 846.600 ;
        RECT 628.950 844.950 631.050 845.400 ;
        RECT 718.950 844.950 721.050 845.400 ;
        RECT 727.950 846.600 730.050 847.050 ;
        RECT 760.950 846.600 763.050 847.050 ;
        RECT 727.950 845.400 763.050 846.600 ;
        RECT 727.950 844.950 730.050 845.400 ;
        RECT 760.950 844.950 763.050 845.400 ;
        RECT 772.950 846.600 775.050 847.050 ;
        RECT 805.950 846.600 808.050 847.050 ;
        RECT 772.950 845.400 808.050 846.600 ;
        RECT 772.950 844.950 775.050 845.400 ;
        RECT 805.950 844.950 808.050 845.400 ;
        RECT 919.950 846.600 922.050 847.050 ;
        RECT 925.950 846.600 928.050 847.050 ;
        RECT 919.950 845.400 928.050 846.600 ;
        RECT 919.950 844.950 922.050 845.400 ;
        RECT 925.950 844.950 928.050 845.400 ;
        RECT 1018.950 846.600 1021.050 847.050 ;
        RECT 1033.950 846.600 1036.050 847.050 ;
        RECT 1018.950 845.400 1036.050 846.600 ;
        RECT 1018.950 844.950 1021.050 845.400 ;
        RECT 1033.950 844.950 1036.050 845.400 ;
        RECT 382.950 843.600 385.050 844.050 ;
        RECT 371.400 842.400 385.050 843.600 ;
        RECT 253.950 841.950 256.050 842.400 ;
        RECT 277.950 841.950 280.050 842.400 ;
        RECT 382.950 841.950 385.050 842.400 ;
        RECT 625.950 843.600 628.050 844.050 ;
        RECT 661.950 843.600 664.050 844.200 ;
        RECT 625.950 842.400 664.050 843.600 ;
        RECT 625.950 841.950 628.050 842.400 ;
        RECT 661.950 842.100 664.050 842.400 ;
        RECT 688.950 843.600 691.050 844.050 ;
        RECT 715.950 843.600 718.050 844.050 ;
        RECT 688.950 842.400 718.050 843.600 ;
        RECT 688.950 841.950 691.050 842.400 ;
        RECT 715.950 841.950 718.050 842.400 ;
        RECT 820.950 843.600 823.050 844.050 ;
        RECT 826.950 843.600 829.050 844.050 ;
        RECT 820.950 842.400 829.050 843.600 ;
        RECT 820.950 841.950 823.050 842.400 ;
        RECT 826.950 841.950 829.050 842.400 ;
        RECT 931.950 843.600 934.050 844.050 ;
        RECT 943.950 843.600 946.050 844.050 ;
        RECT 931.950 842.400 946.050 843.600 ;
        RECT 931.950 841.950 934.050 842.400 ;
        RECT 943.950 841.950 946.050 842.400 ;
        RECT 985.950 843.600 988.050 844.050 ;
        RECT 1012.950 843.600 1015.050 844.050 ;
        RECT 985.950 842.400 1015.050 843.600 ;
        RECT 985.950 841.950 988.050 842.400 ;
        RECT 1012.950 841.950 1015.050 842.400 ;
        RECT 124.950 840.600 127.050 841.050 ;
        RECT 136.950 840.600 139.050 841.200 ;
        RECT 124.950 839.400 139.050 840.600 ;
        RECT 124.950 838.950 127.050 839.400 ;
        RECT 136.950 839.100 139.050 839.400 ;
        RECT 157.950 840.750 160.050 841.200 ;
        RECT 172.950 840.750 175.050 841.200 ;
        RECT 157.950 839.550 175.050 840.750 ;
        RECT 157.950 839.100 160.050 839.550 ;
        RECT 172.950 839.100 175.050 839.550 ;
        RECT 187.950 840.600 190.050 841.200 ;
        RECT 193.950 840.600 196.050 841.050 ;
        RECT 187.950 839.400 196.050 840.600 ;
        RECT 187.950 839.100 190.050 839.400 ;
        RECT 193.950 838.950 196.050 839.400 ;
        RECT 199.950 840.600 202.050 841.050 ;
        RECT 217.950 840.600 220.050 841.200 ;
        RECT 238.950 840.600 241.050 841.200 ;
        RECT 250.950 840.750 253.050 841.200 ;
        RECT 259.950 840.750 262.050 841.200 ;
        RECT 199.950 839.400 249.600 840.600 ;
        RECT 199.950 838.950 202.050 839.400 ;
        RECT 217.950 839.100 220.050 839.400 ;
        RECT 238.950 839.100 241.050 839.400 ;
        RECT 88.950 837.600 91.050 837.900 ;
        RECT 248.400 837.600 249.600 839.400 ;
        RECT 250.950 839.550 262.050 840.750 ;
        RECT 250.950 839.100 253.050 839.550 ;
        RECT 259.950 839.100 262.050 839.550 ;
        RECT 274.950 840.750 277.050 841.200 ;
        RECT 286.950 840.750 289.050 841.200 ;
        RECT 274.950 840.600 289.050 840.750 ;
        RECT 307.800 840.600 309.900 841.050 ;
        RECT 274.950 839.550 309.900 840.600 ;
        RECT 274.950 839.100 277.050 839.550 ;
        RECT 286.950 839.400 309.900 839.550 ;
        RECT 286.950 839.100 289.050 839.400 ;
        RECT 307.800 838.950 309.900 839.400 ;
        RECT 310.950 840.750 313.050 841.200 ;
        RECT 319.950 840.750 322.050 841.200 ;
        RECT 310.950 839.550 322.050 840.750 ;
        RECT 310.950 839.100 313.050 839.550 ;
        RECT 319.950 839.100 322.050 839.550 ;
        RECT 334.950 839.100 337.050 841.200 ;
        RECT 340.950 840.600 343.050 841.200 ;
        RECT 364.950 840.600 367.050 841.200 ;
        RECT 409.950 840.600 412.050 841.200 ;
        RECT 340.950 839.400 367.050 840.600 ;
        RECT 340.950 839.100 343.050 839.400 ;
        RECT 364.950 839.100 367.050 839.400 ;
        RECT 377.400 839.400 412.050 840.600 ;
        RECT 335.400 837.600 336.600 839.100 ;
        RECT 88.950 836.400 132.600 837.600 ;
        RECT 248.400 836.400 336.600 837.600 ;
        RECT 352.950 837.600 355.050 838.050 ;
        RECT 377.400 837.600 378.600 839.400 ;
        RECT 409.950 839.100 412.050 839.400 ;
        RECT 421.950 840.750 424.050 841.200 ;
        RECT 427.950 840.750 430.050 841.200 ;
        RECT 421.950 839.550 430.050 840.750 ;
        RECT 421.950 839.100 424.050 839.550 ;
        RECT 427.950 839.100 430.050 839.550 ;
        RECT 457.950 840.600 460.050 841.200 ;
        RECT 463.950 840.600 466.050 841.050 ;
        RECT 457.950 839.400 466.050 840.600 ;
        RECT 457.950 839.100 460.050 839.400 ;
        RECT 463.950 838.950 466.050 839.400 ;
        RECT 481.950 839.100 484.050 841.200 ;
        RECT 535.950 839.100 538.050 841.200 ;
        RECT 541.950 840.750 544.050 841.200 ;
        RECT 550.950 840.750 553.050 841.200 ;
        RECT 541.950 839.550 553.050 840.750 ;
        RECT 541.950 839.100 544.050 839.550 ;
        RECT 550.950 839.100 553.050 839.550 ;
        RECT 559.950 840.750 562.050 841.200 ;
        RECT 571.950 840.750 574.050 841.200 ;
        RECT 559.950 839.550 574.050 840.750 ;
        RECT 559.950 839.100 562.050 839.550 ;
        RECT 571.950 839.100 574.050 839.550 ;
        RECT 586.950 840.600 589.050 841.200 ;
        RECT 613.950 840.600 616.050 841.200 ;
        RECT 628.950 840.600 631.050 841.050 ;
        RECT 586.950 839.400 631.050 840.600 ;
        RECT 586.950 839.100 589.050 839.400 ;
        RECT 613.950 839.100 616.050 839.400 ;
        RECT 352.950 836.400 378.600 837.600 ;
        RECT 88.950 835.800 91.050 836.400 ;
        RECT 115.950 834.450 118.050 834.900 ;
        RECT 124.950 834.450 127.050 834.900 ;
        RECT 115.950 833.250 127.050 834.450 ;
        RECT 131.400 834.600 132.600 836.400 ;
        RECT 352.950 835.950 355.050 836.400 ;
        RECT 133.950 834.600 136.050 834.900 ;
        RECT 131.400 834.450 136.050 834.600 ;
        RECT 139.950 834.450 142.050 834.900 ;
        RECT 131.400 833.400 142.050 834.450 ;
        RECT 115.950 832.800 118.050 833.250 ;
        RECT 124.950 832.800 127.050 833.250 ;
        RECT 133.950 833.250 142.050 833.400 ;
        RECT 133.950 832.800 136.050 833.250 ;
        RECT 139.950 832.800 142.050 833.250 ;
        RECT 148.950 834.600 151.050 835.050 ;
        RECT 154.950 834.600 157.050 834.900 ;
        RECT 148.950 833.400 157.050 834.600 ;
        RECT 148.950 832.950 151.050 833.400 ;
        RECT 154.950 832.800 157.050 833.400 ;
        RECT 166.950 834.450 169.050 834.900 ;
        RECT 175.950 834.450 178.050 834.900 ;
        RECT 166.950 833.250 178.050 834.450 ;
        RECT 166.950 832.800 169.050 833.250 ;
        RECT 175.950 832.800 178.050 833.250 ;
        RECT 190.950 834.450 193.050 834.900 ;
        RECT 199.950 834.450 202.050 834.900 ;
        RECT 190.950 833.250 202.050 834.450 ;
        RECT 190.950 832.800 193.050 833.250 ;
        RECT 199.950 832.800 202.050 833.250 ;
        RECT 235.950 834.450 238.050 834.900 ;
        RECT 244.950 834.450 247.050 834.900 ;
        RECT 235.950 833.250 247.050 834.450 ;
        RECT 235.950 832.800 238.050 833.250 ;
        RECT 244.950 832.800 247.050 833.250 ;
        RECT 262.950 834.450 265.050 834.900 ;
        RECT 271.950 834.450 274.050 834.900 ;
        RECT 262.950 833.250 274.050 834.450 ;
        RECT 262.950 832.800 265.050 833.250 ;
        RECT 271.950 832.800 274.050 833.250 ;
        RECT 277.950 834.600 280.050 835.050 ;
        RECT 283.950 834.600 286.050 834.900 ;
        RECT 277.950 833.400 286.050 834.600 ;
        RECT 277.950 832.950 280.050 833.400 ;
        RECT 283.950 832.800 286.050 833.400 ;
        RECT 289.950 834.600 292.050 834.900 ;
        RECT 313.950 834.600 316.050 834.900 ;
        RECT 289.950 833.400 316.050 834.600 ;
        RECT 289.950 832.800 292.050 833.400 ;
        RECT 313.950 832.800 316.050 833.400 ;
        RECT 319.950 834.600 322.050 835.050 ;
        RECT 328.950 834.600 331.050 835.050 ;
        RECT 319.950 833.400 331.050 834.600 ;
        RECT 319.950 832.950 322.050 833.400 ;
        RECT 328.950 832.950 331.050 833.400 ;
        RECT 343.950 834.450 346.050 834.900 ;
        RECT 373.950 834.450 376.050 834.900 ;
        RECT 343.950 833.250 376.050 834.450 ;
        RECT 343.950 832.800 346.050 833.250 ;
        RECT 373.950 832.800 376.050 833.250 ;
        RECT 388.950 834.450 391.050 834.900 ;
        RECT 394.950 834.450 397.050 834.900 ;
        RECT 388.950 833.250 397.050 834.450 ;
        RECT 388.950 832.800 391.050 833.250 ;
        RECT 394.950 832.800 397.050 833.250 ;
        RECT 460.950 834.450 463.050 834.900 ;
        RECT 469.950 834.450 472.050 834.900 ;
        RECT 460.950 833.250 472.050 834.450 ;
        RECT 460.950 832.800 463.050 833.250 ;
        RECT 469.950 832.800 472.050 833.250 ;
        RECT 475.950 834.600 478.050 835.050 ;
        RECT 482.400 834.600 483.600 839.100 ;
        RECT 536.400 837.600 537.600 839.100 ;
        RECT 628.950 838.950 631.050 839.400 ;
        RECT 637.950 840.600 640.050 841.200 ;
        RECT 661.950 840.600 664.050 841.050 ;
        RECT 637.950 839.400 664.050 840.600 ;
        RECT 637.950 839.100 640.050 839.400 ;
        RECT 661.950 838.950 664.050 839.400 ;
        RECT 667.950 840.750 670.050 841.200 ;
        RECT 673.950 840.750 676.050 841.200 ;
        RECT 667.950 839.550 676.050 840.750 ;
        RECT 667.950 839.100 670.050 839.550 ;
        RECT 673.950 839.100 676.050 839.550 ;
        RECT 685.950 840.600 688.050 841.200 ;
        RECT 685.950 839.400 708.600 840.600 ;
        RECT 685.950 839.100 688.050 839.400 ;
        RECT 536.400 836.400 543.600 837.600 ;
        RECT 542.400 835.050 543.600 836.400 ;
        RECT 475.950 833.400 483.600 834.600 ;
        RECT 490.950 834.600 493.050 834.900 ;
        RECT 538.950 834.600 541.050 834.900 ;
        RECT 490.950 833.400 541.050 834.600 ;
        RECT 542.400 833.400 547.050 835.050 ;
        RECT 475.950 832.950 478.050 833.400 ;
        RECT 490.950 832.800 493.050 833.400 ;
        RECT 538.950 832.800 541.050 833.400 ;
        RECT 543.000 832.950 547.050 833.400 ;
        RECT 550.950 834.600 553.050 835.050 ;
        RECT 562.950 834.600 565.050 834.900 ;
        RECT 550.950 833.400 565.050 834.600 ;
        RECT 550.950 832.950 553.050 833.400 ;
        RECT 562.950 832.800 565.050 833.400 ;
        RECT 595.950 834.600 598.050 835.050 ;
        RECT 604.950 834.600 607.050 834.900 ;
        RECT 595.950 834.450 607.050 834.600 ;
        RECT 610.950 834.450 613.050 834.900 ;
        RECT 595.950 833.400 613.050 834.450 ;
        RECT 595.950 832.950 598.050 833.400 ;
        RECT 604.950 833.250 613.050 833.400 ;
        RECT 604.950 832.800 607.050 833.250 ;
        RECT 610.950 832.800 613.050 833.250 ;
        RECT 628.950 834.450 631.050 834.900 ;
        RECT 634.950 834.450 637.050 834.900 ;
        RECT 628.950 833.250 637.050 834.450 ;
        RECT 628.950 832.800 631.050 833.250 ;
        RECT 634.950 832.800 637.050 833.250 ;
        RECT 640.950 834.450 643.050 834.900 ;
        RECT 646.950 834.450 649.050 834.900 ;
        RECT 640.950 833.250 649.050 834.450 ;
        RECT 640.950 832.800 643.050 833.250 ;
        RECT 646.950 832.800 649.050 833.250 ;
        RECT 664.950 834.600 667.050 834.900 ;
        RECT 688.950 834.600 691.050 834.900 ;
        RECT 664.950 833.400 691.050 834.600 ;
        RECT 707.400 834.600 708.600 839.400 ;
        RECT 718.950 837.600 721.050 841.050 ;
        RECT 730.950 840.600 733.050 841.050 ;
        RECT 742.950 840.600 745.050 841.200 ;
        RECT 730.950 839.400 745.050 840.600 ;
        RECT 730.950 838.950 733.050 839.400 ;
        RECT 742.950 839.100 745.050 839.400 ;
        RECT 766.950 840.750 769.050 841.200 ;
        RECT 778.950 840.750 781.050 841.200 ;
        RECT 766.950 840.600 781.050 840.750 ;
        RECT 799.950 840.600 802.050 841.200 ;
        RECT 766.950 839.550 802.050 840.600 ;
        RECT 766.950 839.100 769.050 839.550 ;
        RECT 778.950 839.400 802.050 839.550 ;
        RECT 778.950 839.100 781.050 839.400 ;
        RECT 799.950 839.100 802.050 839.400 ;
        RECT 805.950 840.750 808.050 841.200 ;
        RECT 814.950 840.750 817.050 841.200 ;
        RECT 805.950 839.550 817.050 840.750 ;
        RECT 805.950 839.100 808.050 839.550 ;
        RECT 814.950 839.100 817.050 839.550 ;
        RECT 832.950 839.100 835.050 841.200 ;
        RECT 856.950 840.600 859.050 841.200 ;
        RECT 871.950 840.600 874.050 841.050 ;
        RECT 880.950 840.600 883.050 841.200 ;
        RECT 856.950 839.400 883.050 840.600 ;
        RECT 856.950 839.100 859.050 839.400 ;
        RECT 743.400 837.600 744.600 839.100 ;
        RECT 760.950 837.600 763.050 838.050 ;
        RECT 718.950 837.000 738.600 837.600 ;
        RECT 719.400 836.400 738.600 837.000 ;
        RECT 743.400 836.400 763.050 837.600 ;
        RECT 737.400 834.900 738.600 836.400 ;
        RECT 760.950 835.950 763.050 836.400 ;
        RECT 790.950 837.600 795.000 838.050 ;
        RECT 833.400 837.600 834.600 839.100 ;
        RECT 871.950 838.950 874.050 839.400 ;
        RECT 880.950 839.100 883.050 839.400 ;
        RECT 907.950 839.100 910.050 841.200 ;
        RECT 913.950 840.750 916.050 841.200 ;
        RECT 925.950 840.750 928.050 841.200 ;
        RECT 913.950 839.550 928.050 840.750 ;
        RECT 913.950 839.100 916.050 839.550 ;
        RECT 925.950 839.100 928.050 839.550 ;
        RECT 937.950 839.100 940.050 841.200 ;
        RECT 955.950 840.600 958.050 841.200 ;
        RECT 953.400 839.400 958.050 840.600 ;
        RECT 790.950 835.950 795.600 837.600 ;
        RECT 833.400 836.400 846.600 837.600 ;
        RECT 709.950 834.600 712.050 834.900 ;
        RECT 707.400 833.400 712.050 834.600 ;
        RECT 664.950 832.800 667.050 833.400 ;
        RECT 688.950 832.800 691.050 833.400 ;
        RECT 709.950 832.800 712.050 833.400 ;
        RECT 715.950 834.450 718.050 834.900 ;
        RECT 721.950 834.450 724.050 834.900 ;
        RECT 715.950 833.250 724.050 834.450 ;
        RECT 715.950 832.800 718.050 833.250 ;
        RECT 721.950 832.800 724.050 833.250 ;
        RECT 736.950 834.450 739.050 834.900 ;
        RECT 769.950 834.450 772.050 834.900 ;
        RECT 775.950 834.600 778.050 834.900 ;
        RECT 736.950 833.250 772.050 834.450 ;
        RECT 736.950 832.800 739.050 833.250 ;
        RECT 769.950 832.800 772.050 833.250 ;
        RECT 773.400 833.400 778.050 834.600 ;
        RECT 794.400 834.600 795.600 835.950 ;
        RECT 808.950 834.600 811.050 834.900 ;
        RECT 794.400 833.400 811.050 834.600 ;
        RECT 196.950 831.600 199.050 832.050 ;
        RECT 214.950 831.600 217.050 832.050 ;
        RECT 196.950 830.400 217.050 831.600 ;
        RECT 196.950 829.950 199.050 830.400 ;
        RECT 214.950 829.950 217.050 830.400 ;
        RECT 229.950 831.600 232.050 832.050 ;
        RECT 328.950 831.600 331.050 831.900 ;
        RECT 229.950 830.400 331.050 831.600 ;
        RECT 229.950 829.950 232.050 830.400 ;
        RECT 328.950 829.800 331.050 830.400 ;
        RECT 361.950 831.600 364.050 832.050 ;
        RECT 376.950 831.600 379.050 832.050 ;
        RECT 361.950 830.400 379.050 831.600 ;
        RECT 361.950 829.950 364.050 830.400 ;
        RECT 376.950 829.950 379.050 830.400 ;
        RECT 430.950 831.600 433.050 832.050 ;
        RECT 442.950 831.600 445.050 832.050 ;
        RECT 430.950 830.400 445.050 831.600 ;
        RECT 430.950 829.950 433.050 830.400 ;
        RECT 442.950 829.950 445.050 830.400 ;
        RECT 691.950 831.600 694.050 832.050 ;
        RECT 703.950 831.600 706.050 832.050 ;
        RECT 691.950 830.400 706.050 831.600 ;
        RECT 691.950 829.950 694.050 830.400 ;
        RECT 703.950 829.950 706.050 830.400 ;
        RECT 748.950 831.600 751.050 832.050 ;
        RECT 773.400 831.600 774.600 833.400 ;
        RECT 775.950 832.800 778.050 833.400 ;
        RECT 808.950 832.800 811.050 833.400 ;
        RECT 829.950 834.600 832.050 834.900 ;
        RECT 841.950 834.600 844.050 835.050 ;
        RECT 829.950 833.400 844.050 834.600 ;
        RECT 829.950 832.800 832.050 833.400 ;
        RECT 841.950 832.950 844.050 833.400 ;
        RECT 748.950 830.400 774.600 831.600 ;
        RECT 781.950 831.600 784.050 832.050 ;
        RECT 787.800 831.600 789.900 832.050 ;
        RECT 781.950 830.400 789.900 831.600 ;
        RECT 748.950 829.950 751.050 830.400 ;
        RECT 781.950 829.950 784.050 830.400 ;
        RECT 787.800 829.950 789.900 830.400 ;
        RECT 790.950 831.600 793.050 832.050 ;
        RECT 826.950 831.600 829.050 832.050 ;
        RECT 790.950 830.400 829.050 831.600 ;
        RECT 845.400 831.600 846.600 836.400 ;
        RECT 865.950 834.600 870.000 835.050 ;
        RECT 883.950 834.600 886.050 834.900 ;
        RECT 895.950 834.600 898.050 835.050 ;
        RECT 865.950 832.950 870.600 834.600 ;
        RECT 853.950 831.600 856.050 832.050 ;
        RECT 845.400 830.400 856.050 831.600 ;
        RECT 869.400 831.600 870.600 832.950 ;
        RECT 883.950 833.400 898.050 834.600 ;
        RECT 883.950 832.800 886.050 833.400 ;
        RECT 895.950 832.950 898.050 833.400 ;
        RECT 880.950 831.600 883.050 832.050 ;
        RECT 869.400 830.400 883.050 831.600 ;
        RECT 790.950 829.950 793.050 830.400 ;
        RECT 826.950 829.950 829.050 830.400 ;
        RECT 853.950 829.950 856.050 830.400 ;
        RECT 880.950 829.950 883.050 830.400 ;
        RECT 889.950 831.600 892.050 832.050 ;
        RECT 908.400 831.600 909.600 839.100 ;
        RECT 938.400 835.050 939.600 839.100 ;
        RECT 953.400 835.050 954.600 839.400 ;
        RECT 955.950 839.100 958.050 839.400 ;
        RECT 961.950 839.100 964.050 841.200 ;
        RECT 973.950 840.600 976.050 841.050 ;
        RECT 982.950 840.600 985.050 841.050 ;
        RECT 973.950 839.400 985.050 840.600 ;
        RECT 925.950 834.600 928.050 835.050 ;
        RECT 934.950 834.600 937.050 834.900 ;
        RECT 925.950 833.400 937.050 834.600 ;
        RECT 938.400 833.400 943.050 835.050 ;
        RECT 925.950 832.950 928.050 833.400 ;
        RECT 934.950 832.800 937.050 833.400 ;
        RECT 939.000 832.950 943.050 833.400 ;
        RECT 952.950 832.950 955.050 835.050 ;
        RECT 962.400 832.050 963.600 839.100 ;
        RECT 973.950 838.950 976.050 839.400 ;
        RECT 982.950 838.950 985.050 839.400 ;
        RECT 988.950 839.100 991.050 841.200 ;
        RECT 989.400 835.050 990.600 839.100 ;
        RECT 1003.950 838.950 1006.050 841.050 ;
        RECT 1015.950 838.950 1018.050 841.050 ;
        RECT 1024.950 840.750 1027.050 841.200 ;
        RECT 1030.950 840.750 1033.050 841.200 ;
        RECT 1024.950 839.550 1033.050 840.750 ;
        RECT 1024.950 839.100 1027.050 839.550 ;
        RECT 1030.950 839.100 1033.050 839.550 ;
        RECT 1036.950 839.100 1039.050 841.200 ;
        RECT 1004.400 835.050 1005.600 838.950 ;
        RECT 964.950 834.600 967.050 834.900 ;
        RECT 973.950 834.600 976.050 835.050 ;
        RECT 964.950 833.400 976.050 834.600 ;
        RECT 989.400 833.400 994.050 835.050 ;
        RECT 964.950 832.800 967.050 833.400 ;
        RECT 973.950 832.950 976.050 833.400 ;
        RECT 990.000 832.950 994.050 833.400 ;
        RECT 1003.950 832.950 1006.050 835.050 ;
        RECT 1009.950 834.600 1012.050 834.900 ;
        RECT 1016.400 834.600 1017.600 838.950 ;
        RECT 1009.950 833.400 1017.600 834.600 ;
        RECT 1037.400 834.600 1038.600 839.100 ;
        RECT 1042.950 834.600 1045.050 835.050 ;
        RECT 1037.400 833.400 1045.050 834.600 ;
        RECT 1009.950 832.800 1012.050 833.400 ;
        RECT 1042.950 832.950 1045.050 833.400 ;
        RECT 889.950 830.400 909.600 831.600 ;
        RECT 943.950 831.600 946.050 832.050 ;
        RECT 958.800 831.600 960.900 832.050 ;
        RECT 943.950 830.400 960.900 831.600 ;
        RECT 889.950 829.950 892.050 830.400 ;
        RECT 943.950 829.950 946.050 830.400 ;
        RECT 958.800 829.950 960.900 830.400 ;
        RECT 961.950 829.950 964.050 832.050 ;
        RECT 109.950 828.600 112.050 829.050 ;
        RECT 127.950 828.600 130.050 829.050 ;
        RECT 109.950 827.400 130.050 828.600 ;
        RECT 109.950 826.950 112.050 827.400 ;
        RECT 127.950 826.950 130.050 827.400 ;
        RECT 133.950 828.600 136.050 829.050 ;
        RECT 184.950 828.600 187.050 829.050 ;
        RECT 133.950 827.400 187.050 828.600 ;
        RECT 133.950 826.950 136.050 827.400 ;
        RECT 184.950 826.950 187.050 827.400 ;
        RECT 232.950 828.600 235.050 829.050 ;
        RECT 256.950 828.600 259.050 829.050 ;
        RECT 232.950 827.400 259.050 828.600 ;
        RECT 232.950 826.950 235.050 827.400 ;
        RECT 256.950 826.950 259.050 827.400 ;
        RECT 307.950 828.600 310.050 829.050 ;
        RECT 325.950 828.600 328.050 829.050 ;
        RECT 307.950 827.400 328.050 828.600 ;
        RECT 307.950 826.950 310.050 827.400 ;
        RECT 325.950 826.950 328.050 827.400 ;
        RECT 424.950 828.600 427.050 829.050 ;
        RECT 454.950 828.600 457.050 829.050 ;
        RECT 466.950 828.600 469.050 829.050 ;
        RECT 424.950 827.400 469.050 828.600 ;
        RECT 424.950 826.950 427.050 827.400 ;
        RECT 454.950 826.950 457.050 827.400 ;
        RECT 466.950 826.950 469.050 827.400 ;
        RECT 496.950 828.600 499.050 829.050 ;
        RECT 532.950 828.600 535.050 829.050 ;
        RECT 496.950 827.400 535.050 828.600 ;
        RECT 496.950 826.950 499.050 827.400 ;
        RECT 532.950 826.950 535.050 827.400 ;
        RECT 556.950 828.600 559.050 829.050 ;
        RECT 604.950 828.600 607.050 829.050 ;
        RECT 556.950 827.400 607.050 828.600 ;
        RECT 556.950 826.950 559.050 827.400 ;
        RECT 604.950 826.950 607.050 827.400 ;
        RECT 670.950 828.600 673.050 829.050 ;
        RECT 769.950 828.600 772.050 829.050 ;
        RECT 670.950 827.400 772.050 828.600 ;
        RECT 670.950 826.950 673.050 827.400 ;
        RECT 769.950 826.950 772.050 827.400 ;
        RECT 775.950 828.600 778.050 829.050 ;
        RECT 793.950 828.600 796.050 829.050 ;
        RECT 802.950 828.600 805.050 829.050 ;
        RECT 775.950 827.400 805.050 828.600 ;
        RECT 775.950 826.950 778.050 827.400 ;
        RECT 793.950 826.950 796.050 827.400 ;
        RECT 802.950 826.950 805.050 827.400 ;
        RECT 844.950 828.600 847.050 829.050 ;
        RECT 859.950 828.600 862.050 829.050 ;
        RECT 844.950 827.400 862.050 828.600 ;
        RECT 844.950 826.950 847.050 827.400 ;
        RECT 859.950 826.950 862.050 827.400 ;
        RECT 886.950 828.600 889.050 829.050 ;
        RECT 922.950 828.600 925.050 829.050 ;
        RECT 886.950 827.400 925.050 828.600 ;
        RECT 886.950 826.950 889.050 827.400 ;
        RECT 922.950 826.950 925.050 827.400 ;
        RECT 970.950 828.600 973.050 829.050 ;
        RECT 985.950 828.600 988.050 829.050 ;
        RECT 970.950 827.400 988.050 828.600 ;
        RECT 970.950 826.950 973.050 827.400 ;
        RECT 985.950 826.950 988.050 827.400 ;
        RECT 1006.950 828.600 1009.050 829.050 ;
        RECT 1039.950 828.600 1042.050 829.050 ;
        RECT 1006.950 827.400 1042.050 828.600 ;
        RECT 1006.950 826.950 1009.050 827.400 ;
        RECT 1039.950 826.950 1042.050 827.400 ;
        RECT 22.950 825.600 25.050 826.050 ;
        RECT 76.950 825.600 79.050 826.050 ;
        RECT 22.950 824.400 79.050 825.600 ;
        RECT 22.950 823.950 25.050 824.400 ;
        RECT 76.950 823.950 79.050 824.400 ;
        RECT 130.950 825.600 133.050 826.050 ;
        RECT 199.950 825.600 202.050 826.050 ;
        RECT 130.950 824.400 202.050 825.600 ;
        RECT 130.950 823.950 133.050 824.400 ;
        RECT 199.950 823.950 202.050 824.400 ;
        RECT 316.950 825.600 319.050 826.050 ;
        RECT 361.950 825.600 364.050 826.050 ;
        RECT 316.950 824.400 364.050 825.600 ;
        RECT 316.950 823.950 319.050 824.400 ;
        RECT 361.950 823.950 364.050 824.400 ;
        RECT 394.950 825.600 397.050 826.050 ;
        RECT 400.950 825.600 403.050 826.050 ;
        RECT 394.950 824.400 403.050 825.600 ;
        RECT 394.950 823.950 397.050 824.400 ;
        RECT 400.950 823.950 403.050 824.400 ;
        RECT 418.950 825.600 421.050 826.050 ;
        RECT 445.950 825.600 448.050 826.050 ;
        RECT 469.950 825.600 472.050 826.050 ;
        RECT 484.950 825.600 487.050 826.050 ;
        RECT 418.950 824.400 468.600 825.600 ;
        RECT 418.950 823.950 421.050 824.400 ;
        RECT 445.950 823.950 448.050 824.400 ;
        RECT 37.950 822.600 40.050 823.050 ;
        RECT 58.950 822.600 61.050 823.050 ;
        RECT 37.950 821.400 61.050 822.600 ;
        RECT 37.950 820.950 40.050 821.400 ;
        RECT 58.950 820.950 61.050 821.400 ;
        RECT 94.950 822.600 97.050 823.050 ;
        RECT 157.950 822.600 160.050 823.050 ;
        RECT 94.950 821.400 160.050 822.600 ;
        RECT 94.950 820.950 97.050 821.400 ;
        RECT 157.950 820.950 160.050 821.400 ;
        RECT 172.950 822.600 175.050 823.050 ;
        RECT 193.950 822.600 196.050 823.050 ;
        RECT 232.950 822.600 235.050 823.050 ;
        RECT 172.950 821.400 235.050 822.600 ;
        RECT 172.950 820.950 175.050 821.400 ;
        RECT 193.950 820.950 196.050 821.400 ;
        RECT 232.950 820.950 235.050 821.400 ;
        RECT 328.950 822.600 331.050 823.050 ;
        RECT 352.950 822.600 355.050 823.050 ;
        RECT 328.950 821.400 355.050 822.600 ;
        RECT 328.950 820.950 331.050 821.400 ;
        RECT 352.950 820.950 355.050 821.400 ;
        RECT 367.950 822.600 370.050 823.050 ;
        RECT 460.950 822.600 463.050 823.050 ;
        RECT 367.950 821.400 463.050 822.600 ;
        RECT 467.400 822.600 468.600 824.400 ;
        RECT 469.950 824.400 487.050 825.600 ;
        RECT 469.950 823.950 472.050 824.400 ;
        RECT 484.950 823.950 487.050 824.400 ;
        RECT 544.950 825.600 547.050 826.050 ;
        RECT 598.950 825.600 601.050 826.050 ;
        RECT 658.950 825.600 661.050 826.050 ;
        RECT 544.950 824.400 597.600 825.600 ;
        RECT 544.950 823.950 547.050 824.400 ;
        RECT 478.950 822.600 481.050 823.050 ;
        RECT 484.950 822.600 487.050 822.900 ;
        RECT 467.400 821.400 487.050 822.600 ;
        RECT 367.950 820.950 370.050 821.400 ;
        RECT 460.950 820.950 463.050 821.400 ;
        RECT 478.950 820.950 481.050 821.400 ;
        RECT 484.950 820.800 487.050 821.400 ;
        RECT 502.950 822.600 505.050 823.050 ;
        RECT 514.950 822.600 517.050 823.050 ;
        RECT 541.950 822.600 544.050 823.050 ;
        RECT 502.950 821.400 544.050 822.600 ;
        RECT 502.950 820.950 505.050 821.400 ;
        RECT 514.950 820.950 517.050 821.400 ;
        RECT 541.950 820.950 544.050 821.400 ;
        RECT 574.950 822.600 577.050 823.050 ;
        RECT 589.950 822.600 592.050 823.050 ;
        RECT 574.950 821.400 592.050 822.600 ;
        RECT 596.400 822.600 597.600 824.400 ;
        RECT 598.950 824.400 661.050 825.600 ;
        RECT 598.950 823.950 601.050 824.400 ;
        RECT 658.950 823.950 661.050 824.400 ;
        RECT 700.950 825.600 703.050 826.050 ;
        RECT 721.950 825.600 724.050 826.050 ;
        RECT 700.950 824.400 724.050 825.600 ;
        RECT 700.950 823.950 703.050 824.400 ;
        RECT 721.950 823.950 724.050 824.400 ;
        RECT 733.950 825.600 736.050 826.050 ;
        RECT 742.950 825.600 745.050 826.050 ;
        RECT 766.950 825.600 769.050 826.050 ;
        RECT 733.950 824.400 769.050 825.600 ;
        RECT 733.950 823.950 736.050 824.400 ;
        RECT 742.950 823.950 745.050 824.400 ;
        RECT 766.950 823.950 769.050 824.400 ;
        RECT 799.950 825.600 802.050 826.050 ;
        RECT 820.950 825.600 823.050 826.050 ;
        RECT 799.950 824.400 823.050 825.600 ;
        RECT 799.950 823.950 802.050 824.400 ;
        RECT 820.950 823.950 823.050 824.400 ;
        RECT 850.950 825.600 853.050 826.050 ;
        RECT 856.950 825.600 859.050 826.050 ;
        RECT 850.950 824.400 859.050 825.600 ;
        RECT 850.950 823.950 853.050 824.400 ;
        RECT 856.950 823.950 859.050 824.400 ;
        RECT 868.950 825.600 871.050 826.050 ;
        RECT 940.950 825.600 943.050 826.050 ;
        RECT 961.950 825.600 964.050 826.050 ;
        RECT 868.950 824.400 964.050 825.600 ;
        RECT 868.950 823.950 871.050 824.400 ;
        RECT 940.950 823.950 943.050 824.400 ;
        RECT 961.950 823.950 964.050 824.400 ;
        RECT 1021.950 825.600 1024.050 826.050 ;
        RECT 1033.950 825.600 1036.050 826.050 ;
        RECT 1021.950 824.400 1036.050 825.600 ;
        RECT 1021.950 823.950 1024.050 824.400 ;
        RECT 1033.950 823.950 1036.050 824.400 ;
        RECT 613.950 822.600 616.050 823.050 ;
        RECT 596.400 821.400 616.050 822.600 ;
        RECT 574.950 820.950 577.050 821.400 ;
        RECT 589.950 820.950 592.050 821.400 ;
        RECT 613.950 820.950 616.050 821.400 ;
        RECT 622.950 822.600 625.050 823.050 ;
        RECT 637.950 822.600 640.050 823.050 ;
        RECT 622.950 821.400 640.050 822.600 ;
        RECT 622.950 820.950 625.050 821.400 ;
        RECT 637.950 820.950 640.050 821.400 ;
        RECT 685.950 822.600 688.050 823.050 ;
        RECT 781.950 822.600 784.050 823.050 ;
        RECT 817.950 822.600 820.050 823.050 ;
        RECT 685.950 821.400 820.050 822.600 ;
        RECT 685.950 820.950 688.050 821.400 ;
        RECT 781.950 820.950 784.050 821.400 ;
        RECT 817.950 820.950 820.050 821.400 ;
        RECT 847.950 822.600 850.050 823.050 ;
        RECT 865.950 822.600 868.050 823.050 ;
        RECT 847.950 821.400 868.050 822.600 ;
        RECT 847.950 820.950 850.050 821.400 ;
        RECT 865.950 820.950 868.050 821.400 ;
        RECT 871.950 822.600 874.050 823.050 ;
        RECT 904.950 822.600 907.050 823.050 ;
        RECT 871.950 821.400 907.050 822.600 ;
        RECT 871.950 820.950 874.050 821.400 ;
        RECT 904.950 820.950 907.050 821.400 ;
        RECT 997.950 822.600 1000.050 823.050 ;
        RECT 1039.950 822.600 1042.050 823.050 ;
        RECT 997.950 821.400 1042.050 822.600 ;
        RECT 997.950 820.950 1000.050 821.400 ;
        RECT 1039.950 820.950 1042.050 821.400 ;
        RECT 235.950 819.600 238.050 820.050 ;
        RECT 280.950 819.600 283.050 820.050 ;
        RECT 319.950 819.600 322.050 820.050 ;
        RECT 235.950 818.400 322.050 819.600 ;
        RECT 235.950 817.950 238.050 818.400 ;
        RECT 280.950 817.950 283.050 818.400 ;
        RECT 319.950 817.950 322.050 818.400 ;
        RECT 355.950 819.600 358.050 820.050 ;
        RECT 361.950 819.600 364.050 820.050 ;
        RECT 355.950 818.400 364.050 819.600 ;
        RECT 355.950 817.950 358.050 818.400 ;
        RECT 361.950 817.950 364.050 818.400 ;
        RECT 670.950 819.600 673.050 820.050 ;
        RECT 727.950 819.600 730.050 820.050 ;
        RECT 670.950 818.400 730.050 819.600 ;
        RECT 670.950 817.950 673.050 818.400 ;
        RECT 727.950 817.950 730.050 818.400 ;
        RECT 802.950 819.600 805.050 820.050 ;
        RECT 814.950 819.600 817.050 820.050 ;
        RECT 802.950 818.400 817.050 819.600 ;
        RECT 802.950 817.950 805.050 818.400 ;
        RECT 814.950 817.950 817.050 818.400 ;
        RECT 820.950 819.600 823.050 820.050 ;
        RECT 829.950 819.600 832.050 820.050 ;
        RECT 844.950 819.600 847.050 820.050 ;
        RECT 820.950 818.400 847.050 819.600 ;
        RECT 820.950 817.950 823.050 818.400 ;
        RECT 829.950 817.950 832.050 818.400 ;
        RECT 844.950 817.950 847.050 818.400 ;
        RECT 850.950 819.600 853.050 820.050 ;
        RECT 862.950 819.600 865.050 820.050 ;
        RECT 889.950 819.600 892.050 820.050 ;
        RECT 850.950 818.400 865.050 819.600 ;
        RECT 850.950 817.950 853.050 818.400 ;
        RECT 862.950 817.950 865.050 818.400 ;
        RECT 878.400 818.400 892.050 819.600 ;
        RECT 878.400 817.050 879.600 818.400 ;
        RECT 889.950 817.950 892.050 818.400 ;
        RECT 928.950 819.600 931.050 820.050 ;
        RECT 952.950 819.600 955.050 820.050 ;
        RECT 928.950 818.400 955.050 819.600 ;
        RECT 928.950 817.950 931.050 818.400 ;
        RECT 952.950 817.950 955.050 818.400 ;
        RECT 115.950 816.600 118.050 817.050 ;
        RECT 127.950 816.600 130.050 817.050 ;
        RECT 115.950 815.400 130.050 816.600 ;
        RECT 115.950 814.950 118.050 815.400 ;
        RECT 127.950 814.950 130.050 815.400 ;
        RECT 139.950 816.600 142.050 817.050 ;
        RECT 229.950 816.600 232.050 817.050 ;
        RECT 139.950 815.400 232.050 816.600 ;
        RECT 139.950 814.950 142.050 815.400 ;
        RECT 229.950 814.950 232.050 815.400 ;
        RECT 400.950 816.600 403.050 817.050 ;
        RECT 406.950 816.600 409.050 817.050 ;
        RECT 400.950 815.400 409.050 816.600 ;
        RECT 400.950 814.950 403.050 815.400 ;
        RECT 406.950 814.950 409.050 815.400 ;
        RECT 475.950 816.600 478.050 817.050 ;
        RECT 556.950 816.600 559.050 817.050 ;
        RECT 475.950 815.400 559.050 816.600 ;
        RECT 475.950 814.950 478.050 815.400 ;
        RECT 556.950 814.950 559.050 815.400 ;
        RECT 568.950 816.600 571.050 817.050 ;
        RECT 583.950 816.600 586.050 817.050 ;
        RECT 568.950 815.400 586.050 816.600 ;
        RECT 568.950 814.950 571.050 815.400 ;
        RECT 583.950 814.950 586.050 815.400 ;
        RECT 592.950 816.600 595.050 817.050 ;
        RECT 622.950 816.600 625.050 817.050 ;
        RECT 592.950 815.400 625.050 816.600 ;
        RECT 592.950 814.950 595.050 815.400 ;
        RECT 622.950 814.950 625.050 815.400 ;
        RECT 628.950 816.600 631.050 817.050 ;
        RECT 643.950 816.600 646.050 817.050 ;
        RECT 703.950 816.600 706.050 817.050 ;
        RECT 628.950 815.400 706.050 816.600 ;
        RECT 628.950 814.950 631.050 815.400 ;
        RECT 643.950 814.950 646.050 815.400 ;
        RECT 703.950 814.950 706.050 815.400 ;
        RECT 739.950 816.600 742.050 817.050 ;
        RECT 757.950 816.600 760.050 817.050 ;
        RECT 739.950 815.400 760.050 816.600 ;
        RECT 739.950 814.950 742.050 815.400 ;
        RECT 757.950 814.950 760.050 815.400 ;
        RECT 772.950 816.600 775.050 817.050 ;
        RECT 799.950 816.600 802.050 817.050 ;
        RECT 772.950 815.400 802.050 816.600 ;
        RECT 772.950 814.950 775.050 815.400 ;
        RECT 799.950 814.950 802.050 815.400 ;
        RECT 817.950 816.600 820.050 817.050 ;
        RECT 844.950 816.600 847.050 816.900 ;
        RECT 877.950 816.600 880.050 817.050 ;
        RECT 817.950 815.400 840.600 816.600 ;
        RECT 817.950 814.950 820.050 815.400 ;
        RECT 70.950 813.600 73.050 814.050 ;
        RECT 88.950 813.600 91.050 814.050 ;
        RECT 70.950 812.400 91.050 813.600 ;
        RECT 70.950 811.950 73.050 812.400 ;
        RECT 88.950 811.950 91.050 812.400 ;
        RECT 154.950 813.600 157.050 814.050 ;
        RECT 208.950 813.600 211.050 814.050 ;
        RECT 154.950 812.400 211.050 813.600 ;
        RECT 154.950 811.950 157.050 812.400 ;
        RECT 208.950 811.950 211.050 812.400 ;
        RECT 346.950 813.600 349.050 814.050 ;
        RECT 367.950 813.600 370.050 814.050 ;
        RECT 346.950 812.400 370.050 813.600 ;
        RECT 346.950 811.950 349.050 812.400 ;
        RECT 367.950 811.950 370.050 812.400 ;
        RECT 409.950 813.600 412.050 814.050 ;
        RECT 433.950 813.600 436.050 814.050 ;
        RECT 409.950 812.400 436.050 813.600 ;
        RECT 409.950 811.950 412.050 812.400 ;
        RECT 433.950 811.950 436.050 812.400 ;
        RECT 508.950 813.600 511.050 814.050 ;
        RECT 601.950 813.600 604.050 814.050 ;
        RECT 673.950 813.600 676.050 814.050 ;
        RECT 508.950 812.400 552.600 813.600 ;
        RECT 508.950 811.950 511.050 812.400 ;
        RECT 79.950 810.600 82.050 811.050 ;
        RECT 112.950 810.600 115.050 811.050 ;
        RECT 79.950 809.400 115.050 810.600 ;
        RECT 79.950 808.950 82.050 809.400 ;
        RECT 112.950 808.950 115.050 809.400 ;
        RECT 373.950 810.600 376.050 811.050 ;
        RECT 382.950 810.600 385.050 811.050 ;
        RECT 373.950 809.400 385.050 810.600 ;
        RECT 373.950 808.950 376.050 809.400 ;
        RECT 382.950 808.950 385.050 809.400 ;
        RECT 388.950 810.600 391.050 811.050 ;
        RECT 397.950 810.600 400.050 810.900 ;
        RECT 388.950 809.400 400.050 810.600 ;
        RECT 388.950 808.950 391.050 809.400 ;
        RECT 397.950 808.800 400.050 809.400 ;
        RECT 451.950 810.600 454.050 811.050 ;
        RECT 457.950 810.600 460.050 811.050 ;
        RECT 451.950 809.400 460.050 810.600 ;
        RECT 551.400 810.600 552.600 812.400 ;
        RECT 601.950 812.400 676.050 813.600 ;
        RECT 601.950 811.950 604.050 812.400 ;
        RECT 673.950 811.950 676.050 812.400 ;
        RECT 760.950 813.600 763.050 814.050 ;
        RECT 790.950 813.600 793.050 814.050 ;
        RECT 760.950 812.400 793.050 813.600 ;
        RECT 760.950 811.950 763.050 812.400 ;
        RECT 790.950 811.950 793.050 812.400 ;
        RECT 826.950 813.600 829.050 814.050 ;
        RECT 835.950 813.600 838.050 814.050 ;
        RECT 826.950 812.400 838.050 813.600 ;
        RECT 839.400 813.600 840.600 815.400 ;
        RECT 844.950 815.400 880.050 816.600 ;
        RECT 844.950 814.800 847.050 815.400 ;
        RECT 877.950 814.950 880.050 815.400 ;
        RECT 892.950 816.600 895.050 817.050 ;
        RECT 904.950 816.600 907.050 817.050 ;
        RECT 892.950 815.400 907.050 816.600 ;
        RECT 892.950 814.950 895.050 815.400 ;
        RECT 904.950 814.950 907.050 815.400 ;
        RECT 922.950 816.600 925.050 817.050 ;
        RECT 943.950 816.600 946.050 817.050 ;
        RECT 922.950 815.400 946.050 816.600 ;
        RECT 922.950 814.950 925.050 815.400 ;
        RECT 943.950 814.950 946.050 815.400 ;
        RECT 955.950 816.600 958.050 817.050 ;
        RECT 967.950 816.600 970.050 817.050 ;
        RECT 955.950 815.400 970.050 816.600 ;
        RECT 955.950 814.950 958.050 815.400 ;
        RECT 967.950 814.950 970.050 815.400 ;
        RECT 886.950 813.600 889.050 814.050 ;
        RECT 839.400 812.400 889.050 813.600 ;
        RECT 826.950 811.950 829.050 812.400 ;
        RECT 835.950 811.950 838.050 812.400 ;
        RECT 886.950 811.950 889.050 812.400 ;
        RECT 958.950 813.600 961.050 814.050 ;
        RECT 967.950 813.600 970.050 813.900 ;
        RECT 958.950 812.400 970.050 813.600 ;
        RECT 958.950 811.950 961.050 812.400 ;
        RECT 967.950 811.800 970.050 812.400 ;
        RECT 1009.950 813.600 1012.050 814.050 ;
        RECT 1018.950 813.600 1021.050 814.050 ;
        RECT 1009.950 812.400 1021.050 813.600 ;
        RECT 1009.950 811.950 1012.050 812.400 ;
        RECT 1018.950 811.950 1021.050 812.400 ;
        RECT 562.950 810.600 565.050 811.050 ;
        RECT 551.400 809.400 565.050 810.600 ;
        RECT 451.950 808.950 454.050 809.400 ;
        RECT 457.950 808.950 460.050 809.400 ;
        RECT 562.950 808.950 565.050 809.400 ;
        RECT 604.950 810.600 607.050 811.050 ;
        RECT 652.950 810.600 655.050 811.050 ;
        RECT 604.950 809.400 655.050 810.600 ;
        RECT 604.950 808.950 607.050 809.400 ;
        RECT 652.950 808.950 655.050 809.400 ;
        RECT 682.950 810.600 685.050 811.050 ;
        RECT 718.950 810.600 721.050 811.050 ;
        RECT 754.950 810.600 757.050 811.050 ;
        RECT 682.950 809.400 693.600 810.600 ;
        RECT 682.950 808.950 685.050 809.400 ;
        RECT 103.950 807.600 106.050 808.050 ;
        RECT 118.950 807.600 121.050 808.200 ;
        RECT 139.950 807.600 142.050 808.200 ;
        RECT 103.950 806.400 121.050 807.600 ;
        RECT 103.950 805.950 106.050 806.400 ;
        RECT 118.950 806.100 121.050 806.400 ;
        RECT 134.400 806.400 142.050 807.600 ;
        RECT 6.000 804.600 10.050 805.050 ;
        RECT 5.400 802.950 10.050 804.600 ;
        RECT 55.950 804.750 58.050 805.200 ;
        RECT 73.950 804.750 76.050 805.200 ;
        RECT 55.950 804.600 76.050 804.750 ;
        RECT 130.950 804.600 133.050 805.050 ;
        RECT 55.950 803.550 133.050 804.600 ;
        RECT 55.950 803.100 58.050 803.550 ;
        RECT 73.950 803.400 133.050 803.550 ;
        RECT 73.950 803.100 76.050 803.400 ;
        RECT 130.950 802.950 133.050 803.400 ;
        RECT 5.400 798.900 6.600 802.950 ;
        RECT 79.950 801.450 82.050 801.900 ;
        RECT 85.950 801.450 88.050 801.900 ;
        RECT 79.950 800.250 88.050 801.450 ;
        RECT 79.950 799.800 82.050 800.250 ;
        RECT 85.950 799.800 88.050 800.250 ;
        RECT 91.950 801.450 94.050 801.900 ;
        RECT 103.950 801.450 106.050 801.900 ;
        RECT 91.950 800.250 106.050 801.450 ;
        RECT 91.950 799.800 94.050 800.250 ;
        RECT 103.950 799.800 106.050 800.250 ;
        RECT 109.950 801.600 112.050 802.050 ;
        RECT 121.950 801.600 124.050 801.900 ;
        RECT 109.950 800.400 124.050 801.600 ;
        RECT 109.950 799.950 112.050 800.400 ;
        RECT 121.950 799.800 124.050 800.400 ;
        RECT 134.400 799.050 135.600 806.400 ;
        RECT 139.950 806.100 142.050 806.400 ;
        RECT 145.950 807.600 150.000 808.050 ;
        RECT 154.950 807.600 157.050 808.050 ;
        RECT 214.950 807.600 217.050 808.050 ;
        RECT 229.950 807.600 232.050 808.200 ;
        RECT 145.950 805.950 150.600 807.600 ;
        RECT 154.950 807.000 171.600 807.600 ;
        RECT 154.950 806.400 172.050 807.000 ;
        RECT 154.950 805.950 157.050 806.400 ;
        RECT 4.950 796.800 7.050 798.900 ;
        RECT 133.950 796.950 136.050 799.050 ;
        RECT 149.400 798.900 150.600 805.950 ;
        RECT 169.950 802.950 172.050 806.400 ;
        RECT 214.950 806.400 232.050 807.600 ;
        RECT 214.950 805.950 217.050 806.400 ;
        RECT 229.950 806.100 232.050 806.400 ;
        RECT 250.950 807.750 253.050 808.200 ;
        RECT 259.950 807.750 262.050 808.200 ;
        RECT 250.950 806.550 262.050 807.750 ;
        RECT 250.950 806.100 253.050 806.550 ;
        RECT 259.950 806.100 262.050 806.550 ;
        RECT 292.950 807.750 295.050 808.200 ;
        RECT 301.950 807.750 304.050 808.200 ;
        RECT 292.950 806.550 304.050 807.750 ;
        RECT 292.950 806.100 295.050 806.550 ;
        RECT 301.950 806.100 304.050 806.550 ;
        RECT 355.950 806.100 358.050 808.200 ;
        RECT 390.000 807.600 394.050 808.050 ;
        RECT 356.400 804.600 357.600 806.100 ;
        RECT 389.400 805.950 394.050 807.600 ;
        RECT 415.950 807.750 418.050 808.200 ;
        RECT 427.950 807.750 430.050 808.200 ;
        RECT 415.950 806.550 430.050 807.750 ;
        RECT 415.950 806.100 418.050 806.550 ;
        RECT 427.950 806.100 430.050 806.550 ;
        RECT 448.950 807.750 451.050 808.200 ;
        RECT 490.950 807.750 493.050 808.200 ;
        RECT 448.950 806.550 493.050 807.750 ;
        RECT 448.950 806.100 451.050 806.550 ;
        RECT 490.950 806.100 493.050 806.550 ;
        RECT 499.950 807.600 502.050 808.050 ;
        RECT 505.950 807.600 508.050 808.050 ;
        RECT 499.950 806.400 508.050 807.600 ;
        RECT 499.950 805.950 502.050 806.400 ;
        RECT 505.950 805.950 508.050 806.400 ;
        RECT 514.950 807.600 517.050 808.200 ;
        RECT 526.950 807.600 529.050 808.050 ;
        RECT 514.950 806.400 529.050 807.600 ;
        RECT 514.950 806.100 517.050 806.400 ;
        RECT 526.950 805.950 529.050 806.400 ;
        RECT 535.950 806.100 538.050 808.200 ;
        RECT 541.950 807.600 544.050 808.050 ;
        RECT 565.950 807.600 568.050 808.050 ;
        RECT 574.950 807.600 577.050 808.200 ;
        RECT 541.950 806.400 577.050 807.600 ;
        RECT 389.400 804.600 390.600 805.950 ;
        RECT 311.400 803.400 363.600 804.600 ;
        RECT 262.950 801.450 265.050 801.900 ;
        RECT 277.950 801.600 280.050 801.900 ;
        RECT 311.400 801.600 312.600 803.400 ;
        RECT 277.950 801.450 312.600 801.600 ;
        RECT 262.950 800.400 312.600 801.450 ;
        RECT 322.950 801.600 325.050 802.050 ;
        RECT 358.950 801.600 361.050 801.900 ;
        RECT 322.950 800.400 361.050 801.600 ;
        RECT 262.950 800.250 280.050 800.400 ;
        RECT 262.950 799.800 265.050 800.250 ;
        RECT 277.950 799.800 280.050 800.250 ;
        RECT 322.950 799.950 325.050 800.400 ;
        RECT 358.950 799.800 361.050 800.400 ;
        RECT 362.400 799.050 363.600 803.400 ;
        RECT 386.400 803.400 390.600 804.600 ;
        RECT 386.400 801.900 387.600 803.400 ;
        RECT 536.400 802.050 537.600 806.100 ;
        RECT 541.950 805.950 544.050 806.400 ;
        RECT 565.950 805.950 568.050 806.400 ;
        RECT 574.950 806.100 577.050 806.400 ;
        RECT 580.950 807.600 583.050 808.200 ;
        RECT 595.950 807.600 600.000 808.050 ;
        RECT 613.950 807.600 616.050 808.050 ;
        RECT 679.950 807.750 682.050 808.200 ;
        RECT 688.950 807.750 691.050 808.200 ;
        RECT 580.950 806.400 585.600 807.600 ;
        RECT 580.950 806.100 583.050 806.400 ;
        RECT 584.400 802.050 585.600 806.400 ;
        RECT 595.950 805.950 600.600 807.600 ;
        RECT 613.950 806.400 627.600 807.600 ;
        RECT 613.950 805.950 616.050 806.400 ;
        RECT 367.950 801.450 370.050 801.900 ;
        RECT 379.950 801.450 382.050 801.900 ;
        RECT 367.950 800.250 382.050 801.450 ;
        RECT 367.950 799.800 370.050 800.250 ;
        RECT 379.950 799.800 382.050 800.250 ;
        RECT 385.950 799.800 388.050 801.900 ;
        RECT 397.950 801.450 400.050 801.900 ;
        RECT 406.950 801.450 409.050 801.900 ;
        RECT 397.950 800.250 409.050 801.450 ;
        RECT 397.950 799.800 400.050 800.250 ;
        RECT 406.950 799.800 409.050 800.250 ;
        RECT 421.950 801.600 424.050 802.050 ;
        RECT 430.950 801.600 433.050 802.050 ;
        RECT 421.950 800.400 433.050 801.600 ;
        RECT 421.950 799.950 424.050 800.400 ;
        RECT 430.950 799.950 433.050 800.400 ;
        RECT 466.950 801.600 469.050 801.900 ;
        RECT 487.950 801.600 490.050 801.900 ;
        RECT 466.950 800.400 490.050 801.600 ;
        RECT 466.950 799.800 469.050 800.400 ;
        RECT 487.950 799.800 490.050 800.400 ;
        RECT 526.950 801.450 529.050 801.900 ;
        RECT 532.950 801.450 535.050 801.900 ;
        RECT 526.950 800.250 535.050 801.450 ;
        RECT 536.400 800.400 541.050 802.050 ;
        RECT 526.950 799.800 529.050 800.250 ;
        RECT 532.950 799.800 535.050 800.250 ;
        RECT 537.000 799.950 541.050 800.400 ;
        RECT 544.950 801.600 547.050 802.050 ;
        RECT 553.950 801.600 556.050 801.900 ;
        RECT 544.950 800.400 556.050 801.600 ;
        RECT 544.950 799.950 547.050 800.400 ;
        RECT 553.950 799.800 556.050 800.400 ;
        RECT 562.950 801.600 565.050 802.050 ;
        RECT 571.950 801.600 574.050 802.050 ;
        RECT 562.950 800.400 574.050 801.600 ;
        RECT 562.950 799.950 565.050 800.400 ;
        RECT 571.950 799.950 574.050 800.400 ;
        RECT 583.950 799.950 586.050 802.050 ;
        RECT 599.400 801.900 600.600 805.950 ;
        RECT 626.400 804.600 627.600 806.400 ;
        RECT 679.950 806.550 691.050 807.750 ;
        RECT 679.950 806.100 682.050 806.550 ;
        RECT 688.950 806.100 691.050 806.550 ;
        RECT 667.950 804.600 670.050 805.050 ;
        RECT 626.400 803.400 670.050 804.600 ;
        RECT 692.400 804.600 693.600 809.400 ;
        RECT 718.950 809.400 757.050 810.600 ;
        RECT 718.950 808.950 721.050 809.400 ;
        RECT 754.950 808.950 757.050 809.400 ;
        RECT 865.950 810.600 868.050 811.050 ;
        RECT 877.950 810.600 880.050 811.050 ;
        RECT 865.950 809.400 880.050 810.600 ;
        RECT 865.950 808.950 868.050 809.400 ;
        RECT 877.950 808.950 880.050 809.400 ;
        RECT 925.950 810.600 928.050 811.050 ;
        RECT 946.950 810.600 949.050 811.050 ;
        RECT 925.950 809.400 949.050 810.600 ;
        RECT 925.950 808.950 928.050 809.400 ;
        RECT 946.950 808.950 949.050 809.400 ;
        RECT 982.950 810.600 985.050 811.050 ;
        RECT 994.950 810.600 997.050 811.050 ;
        RECT 982.950 809.400 997.050 810.600 ;
        RECT 982.950 808.950 985.050 809.400 ;
        RECT 994.950 808.950 997.050 809.400 ;
        RECT 709.950 807.750 712.050 808.200 ;
        RECT 715.950 807.750 718.050 808.200 ;
        RECT 709.950 806.550 718.050 807.750 ;
        RECT 709.950 806.100 712.050 806.550 ;
        RECT 715.950 806.100 718.050 806.550 ;
        RECT 745.950 807.750 748.050 808.200 ;
        RECT 760.950 807.750 763.050 808.200 ;
        RECT 745.950 806.550 763.050 807.750 ;
        RECT 745.950 806.100 748.050 806.550 ;
        RECT 760.950 806.100 763.050 806.550 ;
        RECT 775.950 807.750 778.050 808.200 ;
        RECT 787.950 807.750 790.050 808.200 ;
        RECT 775.950 806.550 790.050 807.750 ;
        RECT 775.950 806.100 778.050 806.550 ;
        RECT 787.950 806.100 790.050 806.550 ;
        RECT 802.950 807.750 805.050 808.200 ;
        RECT 811.950 807.750 814.050 808.200 ;
        RECT 802.950 807.600 814.050 807.750 ;
        RECT 823.950 807.600 826.050 808.050 ;
        RECT 802.950 806.550 826.050 807.600 ;
        RECT 802.950 806.100 805.050 806.550 ;
        RECT 811.950 806.400 826.050 806.550 ;
        RECT 811.950 806.100 814.050 806.400 ;
        RECT 823.950 805.950 826.050 806.400 ;
        RECT 769.950 804.600 772.050 805.050 ;
        RECT 847.950 804.600 850.050 808.050 ;
        RECT 856.950 807.750 859.050 808.200 ;
        RECT 862.950 807.750 865.050 808.200 ;
        RECT 856.950 806.550 865.050 807.750 ;
        RECT 856.950 806.100 859.050 806.550 ;
        RECT 862.950 806.100 865.050 806.550 ;
        RECT 889.950 807.600 892.050 808.200 ;
        RECT 907.950 807.600 910.050 808.050 ;
        RECT 889.950 806.400 910.050 807.600 ;
        RECT 889.950 806.100 892.050 806.400 ;
        RECT 907.950 805.950 910.050 806.400 ;
        RECT 916.950 807.600 919.050 808.200 ;
        RECT 937.950 807.600 940.050 808.200 ;
        RECT 961.950 807.600 964.050 808.200 ;
        RECT 979.950 807.600 982.050 808.050 ;
        RECT 916.950 806.400 924.600 807.600 ;
        RECT 916.950 806.100 919.050 806.400 ;
        RECT 692.400 803.400 705.600 804.600 ;
        RECT 667.950 802.950 670.050 803.400 ;
        RECT 598.950 799.800 601.050 801.900 ;
        RECT 604.950 801.450 607.050 801.900 ;
        RECT 616.950 801.450 619.050 801.900 ;
        RECT 604.950 800.250 619.050 801.450 ;
        RECT 604.950 799.800 607.050 800.250 ;
        RECT 616.950 799.800 619.050 800.250 ;
        RECT 643.950 801.450 646.050 801.900 ;
        RECT 655.950 801.450 658.050 801.900 ;
        RECT 643.950 800.250 658.050 801.450 ;
        RECT 643.950 799.800 646.050 800.250 ;
        RECT 655.950 799.800 658.050 800.250 ;
        RECT 688.950 801.600 691.050 802.050 ;
        RECT 700.950 801.600 703.050 801.900 ;
        RECT 688.950 800.400 703.050 801.600 ;
        RECT 704.400 801.600 705.600 803.400 ;
        RECT 769.950 804.000 850.050 804.600 ;
        RECT 923.400 804.600 924.600 806.400 ;
        RECT 937.950 806.400 948.600 807.600 ;
        RECT 937.950 806.100 940.050 806.400 ;
        RECT 769.950 803.400 849.600 804.000 ;
        RECT 923.400 803.400 936.600 804.600 ;
        RECT 769.950 802.950 772.050 803.400 ;
        RECT 727.950 801.600 730.050 801.900 ;
        RECT 704.400 800.400 730.050 801.600 ;
        RECT 688.950 799.950 691.050 800.400 ;
        RECT 700.950 799.800 703.050 800.400 ;
        RECT 727.950 799.800 730.050 800.400 ;
        RECT 736.950 801.600 739.050 801.900 ;
        RECT 745.950 801.600 748.050 802.050 ;
        RECT 736.950 800.400 748.050 801.600 ;
        RECT 736.950 799.800 739.050 800.400 ;
        RECT 745.950 799.950 748.050 800.400 ;
        RECT 757.950 801.600 760.050 801.900 ;
        RECT 784.950 801.600 787.050 801.900 ;
        RECT 757.950 800.400 787.050 801.600 ;
        RECT 148.950 796.800 151.050 798.900 ;
        RECT 238.950 798.600 241.050 799.050 ;
        RECT 256.950 798.600 259.050 799.050 ;
        RECT 238.950 797.400 259.050 798.600 ;
        RECT 362.400 797.400 367.050 799.050 ;
        RECT 238.950 796.950 241.050 797.400 ;
        RECT 256.950 796.950 259.050 797.400 ;
        RECT 363.000 796.950 367.050 797.400 ;
        RECT 412.950 798.600 415.050 799.050 ;
        RECT 496.950 798.600 499.050 799.050 ;
        RECT 412.950 797.400 499.050 798.600 ;
        RECT 412.950 796.950 415.050 797.400 ;
        RECT 496.950 796.950 499.050 797.400 ;
        RECT 508.950 798.600 511.050 799.050 ;
        RECT 520.950 798.600 523.050 799.050 ;
        RECT 508.950 797.400 523.050 798.600 ;
        RECT 746.400 798.600 747.600 799.950 ;
        RECT 757.950 799.800 760.050 800.400 ;
        RECT 784.950 799.800 787.050 800.400 ;
        RECT 814.950 801.600 817.050 801.900 ;
        RECT 859.950 801.600 862.050 802.050 ;
        RECT 814.950 800.400 862.050 801.600 ;
        RECT 814.950 799.800 817.050 800.400 ;
        RECT 859.950 799.950 862.050 800.400 ;
        RECT 886.950 801.600 889.050 802.050 ;
        RECT 935.400 801.900 936.600 803.400 ;
        RECT 947.400 802.050 948.600 806.400 ;
        RECT 961.950 806.400 982.050 807.600 ;
        RECT 961.950 806.100 964.050 806.400 ;
        RECT 979.950 805.950 982.050 806.400 ;
        RECT 1003.950 807.600 1006.050 807.900 ;
        RECT 1015.950 807.600 1018.050 808.200 ;
        RECT 1003.950 806.400 1018.050 807.600 ;
        RECT 1003.950 805.800 1006.050 806.400 ;
        RECT 1015.950 806.100 1018.050 806.400 ;
        RECT 1021.950 807.750 1024.050 808.200 ;
        RECT 1027.950 807.750 1030.050 808.200 ;
        RECT 1021.950 806.550 1030.050 807.750 ;
        RECT 1021.950 806.100 1024.050 806.550 ;
        RECT 1027.950 806.100 1030.050 806.550 ;
        RECT 1033.950 805.950 1036.050 808.050 ;
        RECT 1042.950 805.950 1045.050 808.050 ;
        RECT 1034.400 802.050 1035.600 805.950 ;
        RECT 1043.400 802.050 1044.600 805.950 ;
        RECT 892.950 801.600 895.050 801.900 ;
        RECT 886.950 800.400 895.050 801.600 ;
        RECT 886.950 799.950 889.050 800.400 ;
        RECT 892.950 799.800 895.050 800.400 ;
        RECT 934.950 799.800 937.050 801.900 ;
        RECT 946.950 799.950 949.050 802.050 ;
        RECT 958.950 801.450 961.050 801.900 ;
        RECT 964.950 801.450 967.050 801.900 ;
        RECT 958.950 800.250 967.050 801.450 ;
        RECT 958.950 799.800 961.050 800.250 ;
        RECT 964.950 799.800 967.050 800.250 ;
        RECT 982.950 801.450 985.050 801.900 ;
        RECT 988.950 801.450 991.050 801.900 ;
        RECT 982.950 800.250 991.050 801.450 ;
        RECT 982.950 799.800 985.050 800.250 ;
        RECT 988.950 799.800 991.050 800.250 ;
        RECT 1033.950 799.950 1036.050 802.050 ;
        RECT 1042.950 799.950 1045.050 802.050 ;
        RECT 790.950 798.600 793.050 799.050 ;
        RECT 802.950 798.600 805.050 799.050 ;
        RECT 746.400 797.400 805.050 798.600 ;
        RECT 508.950 796.950 511.050 797.400 ;
        RECT 520.950 796.950 523.050 797.400 ;
        RECT 790.950 796.950 793.050 797.400 ;
        RECT 802.950 796.950 805.050 797.400 ;
        RECT 850.950 798.600 853.050 799.050 ;
        RECT 868.950 798.600 871.050 799.050 ;
        RECT 850.950 797.400 871.050 798.600 ;
        RECT 850.950 796.950 853.050 797.400 ;
        RECT 868.950 796.950 871.050 797.400 ;
        RECT 907.950 798.600 910.050 799.050 ;
        RECT 913.950 798.600 916.050 799.050 ;
        RECT 907.950 797.400 916.050 798.600 ;
        RECT 907.950 796.950 910.050 797.400 ;
        RECT 913.950 796.950 916.050 797.400 ;
        RECT 922.950 798.600 925.050 799.050 ;
        RECT 949.950 798.600 952.050 799.050 ;
        RECT 922.950 797.400 952.050 798.600 ;
        RECT 922.950 796.950 925.050 797.400 ;
        RECT 949.950 796.950 952.050 797.400 ;
        RECT 970.950 798.600 973.050 799.050 ;
        RECT 994.950 798.600 997.050 799.050 ;
        RECT 970.950 797.400 997.050 798.600 ;
        RECT 970.950 796.950 973.050 797.400 ;
        RECT 994.950 796.950 997.050 797.400 ;
        RECT 28.950 795.600 31.050 796.050 ;
        RECT 70.950 795.600 73.050 796.050 ;
        RECT 28.950 794.400 73.050 795.600 ;
        RECT 28.950 793.950 31.050 794.400 ;
        RECT 70.950 793.950 73.050 794.400 ;
        RECT 151.950 795.600 154.050 796.050 ;
        RECT 169.950 795.600 172.050 796.050 ;
        RECT 151.950 794.400 172.050 795.600 ;
        RECT 151.950 793.950 154.050 794.400 ;
        RECT 169.950 793.950 172.050 794.400 ;
        RECT 259.950 795.600 262.050 796.050 ;
        RECT 310.950 795.600 313.050 796.050 ;
        RECT 259.950 794.400 313.050 795.600 ;
        RECT 259.950 793.950 262.050 794.400 ;
        RECT 310.950 793.950 313.050 794.400 ;
        RECT 403.950 795.600 406.050 796.050 ;
        RECT 499.950 795.600 502.050 796.050 ;
        RECT 529.950 795.600 532.050 796.050 ;
        RECT 403.950 794.400 532.050 795.600 ;
        RECT 403.950 793.950 406.050 794.400 ;
        RECT 499.950 793.950 502.050 794.400 ;
        RECT 529.950 793.950 532.050 794.400 ;
        RECT 631.950 795.600 634.050 796.050 ;
        RECT 649.950 795.600 652.050 796.050 ;
        RECT 673.950 795.600 676.050 796.050 ;
        RECT 631.950 794.400 676.050 795.600 ;
        RECT 631.950 793.950 634.050 794.400 ;
        RECT 649.950 793.950 652.050 794.400 ;
        RECT 673.950 793.950 676.050 794.400 ;
        RECT 700.950 795.600 703.050 796.050 ;
        RECT 709.950 795.600 712.050 796.050 ;
        RECT 700.950 794.400 712.050 795.600 ;
        RECT 700.950 793.950 703.050 794.400 ;
        RECT 709.950 793.950 712.050 794.400 ;
        RECT 718.950 795.600 721.050 795.900 ;
        RECT 727.950 795.600 730.050 796.050 ;
        RECT 718.950 794.400 730.050 795.600 ;
        RECT 718.950 793.800 721.050 794.400 ;
        RECT 727.950 793.950 730.050 794.400 ;
        RECT 775.950 795.600 778.050 796.050 ;
        RECT 787.950 795.600 790.050 796.050 ;
        RECT 775.950 794.400 790.050 795.600 ;
        RECT 775.950 793.950 778.050 794.400 ;
        RECT 787.950 793.950 790.050 794.400 ;
        RECT 829.950 795.600 832.050 796.050 ;
        RECT 847.950 795.600 850.050 796.050 ;
        RECT 829.950 794.400 850.050 795.600 ;
        RECT 829.950 793.950 832.050 794.400 ;
        RECT 847.950 793.950 850.050 794.400 ;
        RECT 856.950 795.600 859.050 796.050 ;
        RECT 877.950 795.600 880.050 796.050 ;
        RECT 856.950 794.400 880.050 795.600 ;
        RECT 856.950 793.950 859.050 794.400 ;
        RECT 877.950 793.950 880.050 794.400 ;
        RECT 901.950 795.600 904.050 796.050 ;
        RECT 943.950 795.600 946.050 796.050 ;
        RECT 901.950 794.400 946.050 795.600 ;
        RECT 901.950 793.950 904.050 794.400 ;
        RECT 943.950 793.950 946.050 794.400 ;
        RECT 58.950 792.600 61.050 793.050 ;
        RECT 64.950 792.600 67.050 793.050 ;
        RECT 58.950 791.400 67.050 792.600 ;
        RECT 58.950 790.950 61.050 791.400 ;
        RECT 64.950 790.950 67.050 791.400 ;
        RECT 142.950 792.600 145.050 793.050 ;
        RECT 157.950 792.600 160.050 793.050 ;
        RECT 142.950 791.400 160.050 792.600 ;
        RECT 142.950 790.950 145.050 791.400 ;
        RECT 157.950 790.950 160.050 791.400 ;
        RECT 400.950 792.600 403.050 793.050 ;
        RECT 406.950 792.600 409.050 793.050 ;
        RECT 412.950 792.600 415.050 793.050 ;
        RECT 400.950 791.400 415.050 792.600 ;
        RECT 400.950 790.950 403.050 791.400 ;
        RECT 406.950 790.950 409.050 791.400 ;
        RECT 412.950 790.950 415.050 791.400 ;
        RECT 460.950 792.600 463.050 793.050 ;
        RECT 511.950 792.600 514.050 793.050 ;
        RECT 460.950 791.400 514.050 792.600 ;
        RECT 460.950 790.950 463.050 791.400 ;
        RECT 511.950 790.950 514.050 791.400 ;
        RECT 736.950 792.600 739.050 793.050 ;
        RECT 742.950 792.600 745.050 793.050 ;
        RECT 766.950 792.600 769.050 793.050 ;
        RECT 736.950 791.400 769.050 792.600 ;
        RECT 736.950 790.950 739.050 791.400 ;
        RECT 742.950 790.950 745.050 791.400 ;
        RECT 766.950 790.950 769.050 791.400 ;
        RECT 793.950 792.600 796.050 793.050 ;
        RECT 799.950 792.600 802.050 792.900 ;
        RECT 793.950 791.400 802.050 792.600 ;
        RECT 793.950 790.950 796.050 791.400 ;
        RECT 799.950 790.800 802.050 791.400 ;
        RECT 856.950 792.600 859.050 792.900 ;
        RECT 898.800 792.600 900.900 793.050 ;
        RECT 856.950 791.400 900.900 792.600 ;
        RECT 856.950 790.800 859.050 791.400 ;
        RECT 898.800 790.950 900.900 791.400 ;
        RECT 901.950 792.600 904.050 792.900 ;
        RECT 979.950 792.600 982.050 793.050 ;
        RECT 1009.950 792.600 1012.050 793.050 ;
        RECT 901.950 791.400 933.600 792.600 ;
        RECT 901.950 790.800 904.050 791.400 ;
        RECT 286.950 789.600 289.050 790.050 ;
        RECT 352.950 789.600 355.050 790.050 ;
        RECT 286.950 788.400 355.050 789.600 ;
        RECT 286.950 787.950 289.050 788.400 ;
        RECT 352.950 787.950 355.050 788.400 ;
        RECT 364.950 789.600 367.050 790.050 ;
        RECT 448.950 789.600 451.050 790.050 ;
        RECT 364.950 788.400 451.050 789.600 ;
        RECT 364.950 787.950 367.050 788.400 ;
        RECT 448.950 787.950 451.050 788.400 ;
        RECT 514.950 789.600 517.050 790.050 ;
        RECT 592.950 789.600 595.050 790.050 ;
        RECT 748.950 789.600 751.050 790.050 ;
        RECT 757.950 789.600 760.050 790.050 ;
        RECT 514.950 788.400 595.050 789.600 ;
        RECT 514.950 787.950 517.050 788.400 ;
        RECT 592.950 787.950 595.050 788.400 ;
        RECT 728.400 788.400 735.600 789.600 ;
        RECT 157.950 786.600 160.050 787.050 ;
        RECT 193.950 786.600 196.050 787.050 ;
        RECT 223.950 786.600 226.050 787.050 ;
        RECT 304.950 786.600 307.050 787.050 ;
        RECT 157.950 785.400 196.050 786.600 ;
        RECT 157.950 784.950 160.050 785.400 ;
        RECT 193.950 784.950 196.050 785.400 ;
        RECT 215.400 785.400 307.050 786.600 ;
        RECT 115.950 783.600 118.050 784.050 ;
        RECT 136.950 783.600 139.050 784.050 ;
        RECT 215.400 783.600 216.600 785.400 ;
        RECT 223.950 784.950 226.050 785.400 ;
        RECT 304.950 784.950 307.050 785.400 ;
        RECT 361.950 786.600 364.050 787.050 ;
        RECT 400.950 786.600 403.050 787.050 ;
        RECT 424.950 786.600 427.050 787.050 ;
        RECT 361.950 785.400 427.050 786.600 ;
        RECT 361.950 784.950 364.050 785.400 ;
        RECT 400.950 784.950 403.050 785.400 ;
        RECT 424.950 784.950 427.050 785.400 ;
        RECT 439.950 786.600 442.050 787.050 ;
        RECT 451.950 786.600 454.050 787.050 ;
        RECT 439.950 785.400 454.050 786.600 ;
        RECT 439.950 784.950 442.050 785.400 ;
        RECT 451.950 784.950 454.050 785.400 ;
        RECT 487.950 786.600 490.050 787.050 ;
        RECT 538.950 786.600 541.050 787.050 ;
        RECT 487.950 785.400 541.050 786.600 ;
        RECT 487.950 784.950 490.050 785.400 ;
        RECT 538.950 784.950 541.050 785.400 ;
        RECT 583.950 786.600 586.050 787.050 ;
        RECT 728.400 786.600 729.600 788.400 ;
        RECT 583.950 785.400 729.600 786.600 ;
        RECT 734.400 786.600 735.600 788.400 ;
        RECT 748.950 788.400 760.050 789.600 ;
        RECT 748.950 787.950 751.050 788.400 ;
        RECT 757.950 787.950 760.050 788.400 ;
        RECT 784.950 789.600 787.050 790.050 ;
        RECT 805.950 789.600 808.050 790.050 ;
        RECT 784.950 788.400 808.050 789.600 ;
        RECT 784.950 787.950 787.050 788.400 ;
        RECT 805.950 787.950 808.050 788.400 ;
        RECT 850.950 789.600 853.050 790.050 ;
        RECT 928.950 789.600 931.050 790.050 ;
        RECT 850.950 788.400 931.050 789.600 ;
        RECT 932.400 789.600 933.600 791.400 ;
        RECT 979.950 791.400 1012.050 792.600 ;
        RECT 979.950 790.950 982.050 791.400 ;
        RECT 1009.950 790.950 1012.050 791.400 ;
        RECT 955.950 789.600 958.050 790.050 ;
        RECT 932.400 788.400 958.050 789.600 ;
        RECT 850.950 787.950 853.050 788.400 ;
        RECT 928.950 787.950 931.050 788.400 ;
        RECT 955.950 787.950 958.050 788.400 ;
        RECT 769.950 786.600 772.050 787.050 ;
        RECT 734.400 785.400 772.050 786.600 ;
        RECT 583.950 784.950 586.050 785.400 ;
        RECT 769.950 784.950 772.050 785.400 ;
        RECT 847.950 786.600 850.050 787.050 ;
        RECT 919.950 786.600 922.050 787.050 ;
        RECT 847.950 785.400 922.050 786.600 ;
        RECT 847.950 784.950 850.050 785.400 ;
        RECT 919.950 784.950 922.050 785.400 ;
        RECT 991.950 786.600 994.050 787.050 ;
        RECT 1000.950 786.600 1003.050 787.050 ;
        RECT 991.950 785.400 1003.050 786.600 ;
        RECT 991.950 784.950 994.050 785.400 ;
        RECT 1000.950 784.950 1003.050 785.400 ;
        RECT 115.950 782.400 216.600 783.600 ;
        RECT 427.950 783.600 430.050 784.050 ;
        RECT 457.950 783.600 460.050 784.050 ;
        RECT 427.950 782.400 460.050 783.600 ;
        RECT 115.950 781.950 118.050 782.400 ;
        RECT 136.950 781.950 139.050 782.400 ;
        RECT 427.950 781.950 430.050 782.400 ;
        RECT 457.950 781.950 460.050 782.400 ;
        RECT 601.950 783.600 604.050 784.050 ;
        RECT 634.950 783.600 637.050 784.050 ;
        RECT 697.950 783.600 700.050 784.050 ;
        RECT 601.950 782.400 700.050 783.600 ;
        RECT 601.950 781.950 604.050 782.400 ;
        RECT 634.950 781.950 637.050 782.400 ;
        RECT 697.950 781.950 700.050 782.400 ;
        RECT 730.950 783.600 733.050 784.050 ;
        RECT 772.950 783.600 775.050 784.050 ;
        RECT 730.950 782.400 775.050 783.600 ;
        RECT 730.950 781.950 733.050 782.400 ;
        RECT 772.950 781.950 775.050 782.400 ;
        RECT 778.950 783.600 781.050 784.050 ;
        RECT 796.950 783.600 799.050 784.050 ;
        RECT 778.950 782.400 799.050 783.600 ;
        RECT 778.950 781.950 781.050 782.400 ;
        RECT 796.950 781.950 799.050 782.400 ;
        RECT 805.950 783.600 808.050 784.050 ;
        RECT 820.950 783.600 823.050 784.050 ;
        RECT 805.950 782.400 823.050 783.600 ;
        RECT 805.950 781.950 808.050 782.400 ;
        RECT 820.950 781.950 823.050 782.400 ;
        RECT 841.950 783.600 844.050 784.050 ;
        RECT 859.950 783.600 862.050 784.050 ;
        RECT 841.950 782.400 862.050 783.600 ;
        RECT 841.950 781.950 844.050 782.400 ;
        RECT 859.950 781.950 862.050 782.400 ;
        RECT 943.950 783.600 946.050 784.050 ;
        RECT 961.950 783.600 964.050 784.050 ;
        RECT 943.950 782.400 964.050 783.600 ;
        RECT 943.950 781.950 946.050 782.400 ;
        RECT 961.950 781.950 964.050 782.400 ;
        RECT 976.950 783.600 979.050 784.050 ;
        RECT 988.950 783.600 991.050 784.050 ;
        RECT 976.950 782.400 991.050 783.600 ;
        RECT 976.950 781.950 979.050 782.400 ;
        RECT 988.950 781.950 991.050 782.400 ;
        RECT 1003.950 783.600 1006.050 784.050 ;
        RECT 1039.950 783.600 1042.050 784.050 ;
        RECT 1003.950 782.400 1042.050 783.600 ;
        RECT 1003.950 781.950 1006.050 782.400 ;
        RECT 1039.950 781.950 1042.050 782.400 ;
        RECT 121.950 780.600 124.050 781.050 ;
        RECT 160.950 780.600 163.050 781.050 ;
        RECT 121.950 779.400 163.050 780.600 ;
        RECT 121.950 778.950 124.050 779.400 ;
        RECT 160.950 778.950 163.050 779.400 ;
        RECT 172.950 780.600 175.050 781.050 ;
        RECT 184.950 780.600 187.050 781.050 ;
        RECT 172.950 779.400 187.050 780.600 ;
        RECT 172.950 778.950 175.050 779.400 ;
        RECT 184.950 778.950 187.050 779.400 ;
        RECT 217.950 780.600 220.050 781.050 ;
        RECT 295.950 780.600 298.050 781.050 ;
        RECT 217.950 779.400 298.050 780.600 ;
        RECT 217.950 778.950 220.050 779.400 ;
        RECT 295.950 778.950 298.050 779.400 ;
        RECT 484.950 780.600 487.050 781.050 ;
        RECT 514.950 780.600 517.050 781.050 ;
        RECT 484.950 779.400 517.050 780.600 ;
        RECT 484.950 778.950 487.050 779.400 ;
        RECT 514.950 778.950 517.050 779.400 ;
        RECT 559.950 780.600 562.050 781.050 ;
        RECT 568.950 780.600 571.050 781.050 ;
        RECT 559.950 779.400 571.050 780.600 ;
        RECT 559.950 778.950 562.050 779.400 ;
        RECT 568.950 778.950 571.050 779.400 ;
        RECT 823.950 780.600 826.050 781.050 ;
        RECT 856.950 780.600 859.050 781.050 ;
        RECT 823.950 779.400 859.050 780.600 ;
        RECT 823.950 778.950 826.050 779.400 ;
        RECT 856.950 778.950 859.050 779.400 ;
        RECT 862.950 780.600 865.050 781.050 ;
        RECT 880.950 780.600 883.050 781.050 ;
        RECT 895.950 780.600 898.050 781.050 ;
        RECT 862.950 779.400 898.050 780.600 ;
        RECT 862.950 778.950 865.050 779.400 ;
        RECT 880.950 778.950 883.050 779.400 ;
        RECT 895.950 778.950 898.050 779.400 ;
        RECT 919.950 780.600 922.050 781.050 ;
        RECT 970.950 780.600 973.050 781.050 ;
        RECT 919.950 779.400 973.050 780.600 ;
        RECT 919.950 778.950 922.050 779.400 ;
        RECT 970.950 778.950 973.050 779.400 ;
        RECT 334.950 777.600 337.050 778.050 ;
        RECT 373.950 777.600 376.050 778.050 ;
        RECT 334.950 776.400 376.050 777.600 ;
        RECT 334.950 775.950 337.050 776.400 ;
        RECT 373.950 775.950 376.050 776.400 ;
        RECT 445.950 777.600 448.050 778.050 ;
        RECT 499.950 777.600 502.050 778.050 ;
        RECT 445.950 776.400 502.050 777.600 ;
        RECT 445.950 775.950 448.050 776.400 ;
        RECT 499.950 775.950 502.050 776.400 ;
        RECT 577.950 777.600 580.050 778.050 ;
        RECT 595.950 777.600 598.050 778.050 ;
        RECT 577.950 776.400 598.050 777.600 ;
        RECT 577.950 775.950 580.050 776.400 ;
        RECT 595.950 775.950 598.050 776.400 ;
        RECT 625.950 777.600 628.050 778.050 ;
        RECT 631.950 777.600 634.050 778.050 ;
        RECT 625.950 776.400 634.050 777.600 ;
        RECT 625.950 775.950 628.050 776.400 ;
        RECT 631.950 775.950 634.050 776.400 ;
        RECT 670.950 777.600 673.050 778.050 ;
        RECT 703.950 777.600 706.050 778.050 ;
        RECT 670.950 776.400 706.050 777.600 ;
        RECT 670.950 775.950 673.050 776.400 ;
        RECT 703.950 775.950 706.050 776.400 ;
        RECT 712.950 777.600 715.050 778.050 ;
        RECT 796.950 777.600 799.050 778.050 ;
        RECT 712.950 776.400 799.050 777.600 ;
        RECT 712.950 775.950 715.050 776.400 ;
        RECT 796.950 775.950 799.050 776.400 ;
        RECT 805.950 777.600 808.050 778.050 ;
        RECT 847.950 777.600 850.050 778.050 ;
        RECT 805.950 776.400 850.050 777.600 ;
        RECT 805.950 775.950 808.050 776.400 ;
        RECT 847.950 775.950 850.050 776.400 ;
        RECT 898.950 777.600 901.050 778.050 ;
        RECT 937.950 777.600 940.050 778.050 ;
        RECT 898.950 776.400 940.050 777.600 ;
        RECT 898.950 775.950 901.050 776.400 ;
        RECT 937.950 775.950 940.050 776.400 ;
        RECT 952.950 777.600 955.050 778.050 ;
        RECT 967.950 777.600 970.050 778.050 ;
        RECT 952.950 776.400 970.050 777.600 ;
        RECT 952.950 775.950 955.050 776.400 ;
        RECT 967.950 775.950 970.050 776.400 ;
        RECT 67.950 774.600 70.050 775.050 ;
        RECT 163.950 774.600 166.050 775.050 ;
        RECT 67.950 773.400 166.050 774.600 ;
        RECT 67.950 772.950 70.050 773.400 ;
        RECT 163.950 772.950 166.050 773.400 ;
        RECT 244.950 774.600 247.050 775.050 ;
        RECT 379.950 774.600 382.050 775.050 ;
        RECT 502.950 774.600 505.050 775.050 ;
        RECT 244.950 773.400 505.050 774.600 ;
        RECT 244.950 772.950 247.050 773.400 ;
        RECT 379.950 772.950 382.050 773.400 ;
        RECT 502.950 772.950 505.050 773.400 ;
        RECT 571.950 774.600 574.050 775.050 ;
        RECT 607.950 774.600 610.050 775.050 ;
        RECT 571.950 773.400 610.050 774.600 ;
        RECT 571.950 772.950 574.050 773.400 ;
        RECT 607.950 772.950 610.050 773.400 ;
        RECT 688.950 774.600 691.050 775.050 ;
        RECT 718.800 774.600 720.900 775.050 ;
        RECT 688.950 773.400 720.900 774.600 ;
        RECT 688.950 772.950 691.050 773.400 ;
        RECT 718.800 772.950 720.900 773.400 ;
        RECT 721.950 774.600 724.050 775.050 ;
        RECT 748.950 774.600 751.050 775.050 ;
        RECT 721.950 773.400 751.050 774.600 ;
        RECT 797.400 774.600 798.600 775.950 ;
        RECT 871.950 774.600 874.050 775.050 ;
        RECT 797.400 773.400 874.050 774.600 ;
        RECT 721.950 772.950 724.050 773.400 ;
        RECT 748.950 772.950 751.050 773.400 ;
        RECT 871.950 772.950 874.050 773.400 ;
        RECT 883.950 774.600 886.050 775.050 ;
        RECT 943.950 774.600 946.050 775.050 ;
        RECT 994.950 774.600 997.050 775.050 ;
        RECT 1033.950 774.600 1036.050 775.050 ;
        RECT 883.950 773.400 936.600 774.600 ;
        RECT 883.950 772.950 886.050 773.400 ;
        RECT 103.950 771.600 106.050 772.050 ;
        RECT 130.950 771.600 133.050 772.050 ;
        RECT 103.950 770.400 133.050 771.600 ;
        RECT 103.950 769.950 106.050 770.400 ;
        RECT 130.950 769.950 133.050 770.400 ;
        RECT 382.950 771.600 385.050 772.050 ;
        RECT 394.950 771.600 397.050 772.050 ;
        RECT 382.950 770.400 397.050 771.600 ;
        RECT 382.950 769.950 385.050 770.400 ;
        RECT 394.950 769.950 397.050 770.400 ;
        RECT 409.950 771.600 412.050 772.050 ;
        RECT 472.950 771.600 475.050 772.050 ;
        RECT 409.950 770.400 475.050 771.600 ;
        RECT 409.950 769.950 412.050 770.400 ;
        RECT 472.950 769.950 475.050 770.400 ;
        RECT 499.950 771.600 502.050 772.050 ;
        RECT 544.950 771.600 547.050 772.050 ;
        RECT 499.950 770.400 547.050 771.600 ;
        RECT 499.950 769.950 502.050 770.400 ;
        RECT 544.950 769.950 547.050 770.400 ;
        RECT 589.950 771.600 592.050 772.050 ;
        RECT 610.950 771.600 613.050 772.050 ;
        RECT 676.950 771.600 679.050 772.050 ;
        RECT 685.950 771.600 688.050 772.050 ;
        RECT 763.950 771.600 766.050 772.050 ;
        RECT 841.950 771.600 844.050 772.050 ;
        RECT 589.950 770.400 688.050 771.600 ;
        RECT 589.950 769.950 592.050 770.400 ;
        RECT 610.950 769.950 613.050 770.400 ;
        RECT 676.950 769.950 679.050 770.400 ;
        RECT 685.950 769.950 688.050 770.400 ;
        RECT 755.400 770.400 844.050 771.600 ;
        RECT 52.950 768.600 55.050 769.050 ;
        RECT 91.950 768.600 94.050 769.050 ;
        RECT 133.950 768.600 136.050 769.050 ;
        RECT 52.950 767.400 136.050 768.600 ;
        RECT 52.950 766.950 55.050 767.400 ;
        RECT 91.950 766.950 94.050 767.400 ;
        RECT 133.950 766.950 136.050 767.400 ;
        RECT 232.950 768.600 235.050 769.050 ;
        RECT 271.950 768.600 274.050 769.050 ;
        RECT 277.950 768.600 280.050 769.050 ;
        RECT 331.950 768.600 334.050 769.050 ;
        RECT 232.950 767.400 334.050 768.600 ;
        RECT 232.950 766.950 235.050 767.400 ;
        RECT 271.950 766.950 274.050 767.400 ;
        RECT 277.950 766.950 280.050 767.400 ;
        RECT 331.950 766.950 334.050 767.400 ;
        RECT 388.950 768.600 391.050 769.050 ;
        RECT 490.950 768.600 493.050 769.050 ;
        RECT 388.950 767.400 493.050 768.600 ;
        RECT 388.950 766.950 391.050 767.400 ;
        RECT 490.950 766.950 493.050 767.400 ;
        RECT 565.950 768.600 568.050 769.050 ;
        RECT 580.950 768.600 583.050 769.050 ;
        RECT 565.950 767.400 583.050 768.600 ;
        RECT 565.950 766.950 568.050 767.400 ;
        RECT 580.950 766.950 583.050 767.400 ;
        RECT 637.950 768.600 640.050 769.050 ;
        RECT 706.950 768.600 709.050 769.050 ;
        RECT 755.400 768.600 756.600 770.400 ;
        RECT 763.950 769.950 766.050 770.400 ;
        RECT 841.950 769.950 844.050 770.400 ;
        RECT 874.950 771.600 877.050 772.050 ;
        RECT 913.950 771.600 916.050 772.050 ;
        RECT 874.950 770.400 916.050 771.600 ;
        RECT 874.950 769.950 877.050 770.400 ;
        RECT 913.950 769.950 916.050 770.400 ;
        RECT 919.950 771.600 922.050 772.050 ;
        RECT 931.950 771.600 934.050 772.050 ;
        RECT 919.950 770.400 934.050 771.600 ;
        RECT 935.400 771.600 936.600 773.400 ;
        RECT 943.950 773.400 987.600 774.600 ;
        RECT 943.950 772.950 946.050 773.400 ;
        RECT 964.800 771.600 966.900 772.050 ;
        RECT 935.400 770.400 966.900 771.600 ;
        RECT 919.950 769.950 922.050 770.400 ;
        RECT 931.950 769.950 934.050 770.400 ;
        RECT 964.800 769.950 966.900 770.400 ;
        RECT 967.950 771.600 970.050 772.050 ;
        RECT 986.400 771.600 987.600 773.400 ;
        RECT 994.950 773.400 1036.050 774.600 ;
        RECT 994.950 772.950 997.050 773.400 ;
        RECT 1033.950 772.950 1036.050 773.400 ;
        RECT 1036.950 771.600 1039.050 772.050 ;
        RECT 967.950 770.400 981.600 771.600 ;
        RECT 986.400 770.400 1039.050 771.600 ;
        RECT 967.950 769.950 970.050 770.400 ;
        RECT 637.950 767.400 756.600 768.600 ;
        RECT 757.950 768.600 760.050 769.050 ;
        RECT 814.950 768.600 817.050 769.050 ;
        RECT 853.950 768.600 856.050 769.050 ;
        RECT 865.950 768.600 868.050 769.050 ;
        RECT 757.950 767.400 868.050 768.600 ;
        RECT 637.950 766.950 640.050 767.400 ;
        RECT 706.950 766.950 709.050 767.400 ;
        RECT 757.950 766.950 760.050 767.400 ;
        RECT 814.950 766.950 817.050 767.400 ;
        RECT 853.950 766.950 856.050 767.400 ;
        RECT 865.950 766.950 868.050 767.400 ;
        RECT 886.950 768.600 889.050 769.050 ;
        RECT 898.950 768.600 901.050 769.050 ;
        RECT 886.950 767.400 901.050 768.600 ;
        RECT 886.950 766.950 889.050 767.400 ;
        RECT 898.950 766.950 901.050 767.400 ;
        RECT 937.950 768.600 940.050 769.050 ;
        RECT 973.950 768.600 976.050 769.050 ;
        RECT 937.950 767.400 976.050 768.600 ;
        RECT 980.400 768.600 981.600 770.400 ;
        RECT 1036.950 769.950 1039.050 770.400 ;
        RECT 1027.950 768.600 1030.050 769.050 ;
        RECT 980.400 767.400 1030.050 768.600 ;
        RECT 937.950 766.950 940.050 767.400 ;
        RECT 973.950 766.950 976.050 767.400 ;
        RECT 1027.950 766.950 1030.050 767.400 ;
        RECT 1042.950 768.600 1047.000 769.050 ;
        RECT 1042.950 766.950 1047.600 768.600 ;
        RECT 109.950 765.600 112.050 766.050 ;
        RECT 139.950 765.600 142.050 766.050 ;
        RECT 109.950 764.400 142.050 765.600 ;
        RECT 109.950 763.950 112.050 764.400 ;
        RECT 139.950 763.950 142.050 764.400 ;
        RECT 193.950 765.600 196.050 766.050 ;
        RECT 214.950 765.600 217.050 766.050 ;
        RECT 193.950 764.400 217.050 765.600 ;
        RECT 193.950 763.950 196.050 764.400 ;
        RECT 214.950 763.950 217.050 764.400 ;
        RECT 337.950 765.600 340.050 766.050 ;
        RECT 355.950 765.600 358.050 766.050 ;
        RECT 337.950 764.400 358.050 765.600 ;
        RECT 337.950 763.950 340.050 764.400 ;
        RECT 355.950 763.950 358.050 764.400 ;
        RECT 535.950 765.600 538.050 766.050 ;
        RECT 547.950 765.600 550.050 766.050 ;
        RECT 535.950 764.400 550.050 765.600 ;
        RECT 535.950 763.950 538.050 764.400 ;
        RECT 547.950 763.950 550.050 764.400 ;
        RECT 682.950 765.600 685.050 766.050 ;
        RECT 694.950 765.600 697.050 766.050 ;
        RECT 682.950 764.400 697.050 765.600 ;
        RECT 682.950 763.950 685.050 764.400 ;
        RECT 694.950 763.950 697.050 764.400 ;
        RECT 733.950 765.600 736.050 766.050 ;
        RECT 739.950 765.600 742.050 766.050 ;
        RECT 733.950 764.400 742.050 765.600 ;
        RECT 733.950 763.950 736.050 764.400 ;
        RECT 739.950 763.950 742.050 764.400 ;
        RECT 769.950 765.600 772.050 766.050 ;
        RECT 805.950 765.600 808.050 766.050 ;
        RECT 769.950 764.400 808.050 765.600 ;
        RECT 769.950 763.950 772.050 764.400 ;
        RECT 805.950 763.950 808.050 764.400 ;
        RECT 871.950 765.600 874.050 766.050 ;
        RECT 883.950 765.600 886.050 766.050 ;
        RECT 871.950 764.400 886.050 765.600 ;
        RECT 871.950 763.950 874.050 764.400 ;
        RECT 883.950 763.950 886.050 764.400 ;
        RECT 892.950 765.600 895.050 766.050 ;
        RECT 907.950 765.600 910.050 766.050 ;
        RECT 892.950 764.400 910.050 765.600 ;
        RECT 892.950 763.950 895.050 764.400 ;
        RECT 907.950 763.950 910.050 764.400 ;
        RECT 913.950 765.600 916.050 766.050 ;
        RECT 919.950 765.600 922.050 765.900 ;
        RECT 913.950 764.400 922.050 765.600 ;
        RECT 913.950 763.950 916.050 764.400 ;
        RECT 919.950 763.800 922.050 764.400 ;
        RECT 928.950 765.600 931.050 766.050 ;
        RECT 928.950 764.400 942.600 765.600 ;
        RECT 928.950 763.950 931.050 764.400 ;
        RECT 25.950 762.750 28.050 763.200 ;
        RECT 43.950 762.750 46.050 763.200 ;
        RECT 25.950 761.550 46.050 762.750 ;
        RECT 82.950 762.600 85.050 763.200 ;
        RECT 25.950 761.100 28.050 761.550 ;
        RECT 43.950 761.100 46.050 761.550 ;
        RECT 62.400 761.400 85.050 762.600 ;
        RECT 62.400 759.600 63.600 761.400 ;
        RECT 82.950 761.100 85.050 761.400 ;
        RECT 112.950 762.750 115.050 763.200 ;
        RECT 121.950 762.750 124.050 763.200 ;
        RECT 112.950 761.550 124.050 762.750 ;
        RECT 112.950 761.100 115.050 761.550 ;
        RECT 121.950 761.100 124.050 761.550 ;
        RECT 160.950 762.600 163.050 763.050 ;
        RECT 172.950 762.600 175.050 763.200 ;
        RECT 160.950 761.400 175.050 762.600 ;
        RECT 160.950 760.950 163.050 761.400 ;
        RECT 172.950 761.100 175.050 761.400 ;
        RECT 199.950 762.750 202.050 763.200 ;
        RECT 205.950 762.750 208.050 763.200 ;
        RECT 199.950 761.550 208.050 762.750 ;
        RECT 199.950 761.100 202.050 761.550 ;
        RECT 205.950 761.100 208.050 761.550 ;
        RECT 211.950 762.600 214.050 763.050 ;
        RECT 217.950 762.750 220.050 763.200 ;
        RECT 232.950 762.750 235.050 763.200 ;
        RECT 217.950 762.600 235.050 762.750 ;
        RECT 211.950 761.550 235.050 762.600 ;
        RECT 211.950 761.400 220.050 761.550 ;
        RECT 211.950 760.950 214.050 761.400 ;
        RECT 217.950 761.100 220.050 761.400 ;
        RECT 232.950 761.100 235.050 761.550 ;
        RECT 256.950 762.750 259.050 763.200 ;
        RECT 271.950 762.750 274.050 763.200 ;
        RECT 256.950 761.550 274.050 762.750 ;
        RECT 256.950 761.100 259.050 761.550 ;
        RECT 271.950 761.100 274.050 761.550 ;
        RECT 346.950 762.750 349.050 763.200 ;
        RECT 352.950 762.750 355.050 763.200 ;
        RECT 346.950 761.550 355.050 762.750 ;
        RECT 346.950 761.100 349.050 761.550 ;
        RECT 352.950 761.100 355.050 761.550 ;
        RECT 397.950 762.600 400.050 763.200 ;
        RECT 418.950 762.600 421.050 763.200 ;
        RECT 397.950 761.400 421.050 762.600 ;
        RECT 397.950 761.100 400.050 761.400 ;
        RECT 418.950 761.100 421.050 761.400 ;
        RECT 424.950 762.750 427.050 763.200 ;
        RECT 433.950 762.750 436.050 763.200 ;
        RECT 424.950 761.550 436.050 762.750 ;
        RECT 424.950 761.100 427.050 761.550 ;
        RECT 433.950 761.100 436.050 761.550 ;
        RECT 451.950 762.600 454.050 763.200 ;
        RECT 469.950 762.600 472.050 763.200 ;
        RECT 451.950 761.400 472.050 762.600 ;
        RECT 451.950 761.100 454.050 761.400 ;
        RECT 469.950 761.100 472.050 761.400 ;
        RECT 481.950 762.600 484.050 763.050 ;
        RECT 520.950 762.600 523.050 763.200 ;
        RECT 481.950 761.400 523.050 762.600 ;
        RECT 481.950 760.950 484.050 761.400 ;
        RECT 520.950 761.100 523.050 761.400 ;
        RECT 553.950 762.750 556.050 763.200 ;
        RECT 568.950 762.750 571.050 763.200 ;
        RECT 553.950 761.550 571.050 762.750 ;
        RECT 553.950 761.100 556.050 761.550 ;
        RECT 568.950 761.100 571.050 761.550 ;
        RECT 574.950 762.750 577.050 763.200 ;
        RECT 583.950 762.750 586.050 762.900 ;
        RECT 574.950 761.550 586.050 762.750 ;
        RECT 574.950 761.100 577.050 761.550 ;
        RECT 583.950 760.800 586.050 761.550 ;
        RECT 56.400 758.400 63.600 759.600 ;
        RECT 589.950 759.600 592.050 763.050 ;
        RECT 595.950 762.600 598.050 763.200 ;
        RECT 613.950 762.600 616.050 763.050 ;
        RECT 595.950 761.400 616.050 762.600 ;
        RECT 595.950 761.100 598.050 761.400 ;
        RECT 613.950 760.950 616.050 761.400 ;
        RECT 622.950 762.600 625.050 763.200 ;
        RECT 646.950 762.600 649.050 763.200 ;
        RECT 622.950 761.400 649.050 762.600 ;
        RECT 622.950 761.100 625.050 761.400 ;
        RECT 646.950 761.100 649.050 761.400 ;
        RECT 652.950 761.100 655.050 763.200 ;
        RECT 637.950 759.600 640.050 760.050 ;
        RECT 653.400 759.600 654.600 761.100 ;
        RECT 589.950 759.000 603.600 759.600 ;
        RECT 590.400 758.400 603.600 759.000 ;
        RECT 22.950 756.600 25.050 756.900 ;
        RECT 56.400 756.600 57.600 758.400 ;
        RECT 602.400 757.050 603.600 758.400 ;
        RECT 637.950 758.400 654.600 759.600 ;
        RECT 691.950 759.600 694.050 763.050 ;
        RECT 736.950 760.950 739.050 763.050 ;
        RECT 742.950 762.600 745.050 763.200 ;
        RECT 751.950 762.600 754.050 763.050 ;
        RECT 742.950 761.400 754.050 762.600 ;
        RECT 742.950 761.100 745.050 761.400 ;
        RECT 751.950 760.950 754.050 761.400 ;
        RECT 808.950 762.600 811.050 763.200 ;
        RECT 826.950 762.750 829.050 763.200 ;
        RECT 835.950 762.750 838.050 763.200 ;
        RECT 826.950 762.600 838.050 762.750 ;
        RECT 808.950 761.550 838.050 762.600 ;
        RECT 808.950 761.400 829.050 761.550 ;
        RECT 808.950 761.100 811.050 761.400 ;
        RECT 826.950 761.100 829.050 761.400 ;
        RECT 835.950 761.100 838.050 761.550 ;
        RECT 841.950 762.750 844.050 763.200 ;
        RECT 853.800 762.750 855.900 763.200 ;
        RECT 841.950 761.550 855.900 762.750 ;
        RECT 841.950 761.100 844.050 761.550 ;
        RECT 853.800 761.100 855.900 761.550 ;
        RECT 856.950 762.600 859.050 763.050 ;
        RECT 889.950 762.600 892.050 763.200 ;
        RECT 925.950 762.600 928.050 763.050 ;
        RECT 856.950 761.400 892.050 762.600 ;
        RECT 856.950 760.950 859.050 761.400 ;
        RECT 889.950 761.100 892.050 761.400 ;
        RECT 893.400 761.400 928.050 762.600 ;
        RECT 691.950 759.000 702.600 759.600 ;
        RECT 692.400 758.400 702.600 759.000 ;
        RECT 637.950 757.950 640.050 758.400 ;
        RECT 22.950 755.400 57.600 756.600 ;
        RECT 97.950 756.450 100.050 756.900 ;
        RECT 103.950 756.450 106.050 756.900 ;
        RECT 22.950 754.800 25.050 755.400 ;
        RECT 97.950 755.250 106.050 756.450 ;
        RECT 97.950 754.800 100.050 755.250 ;
        RECT 103.950 754.800 106.050 755.250 ;
        RECT 124.950 756.450 127.050 756.900 ;
        RECT 133.950 756.450 136.050 756.900 ;
        RECT 124.950 755.250 136.050 756.450 ;
        RECT 124.950 754.800 127.050 755.250 ;
        RECT 133.950 754.800 136.050 755.250 ;
        RECT 151.950 756.450 154.050 756.900 ;
        RECT 157.950 756.450 160.050 756.900 ;
        RECT 151.950 755.250 160.050 756.450 ;
        RECT 151.950 754.800 154.050 755.250 ;
        RECT 157.950 754.800 160.050 755.250 ;
        RECT 163.950 756.600 166.050 757.050 ;
        RECT 169.950 756.600 172.050 756.900 ;
        RECT 163.950 755.400 172.050 756.600 ;
        RECT 163.950 754.950 166.050 755.400 ;
        RECT 169.950 754.800 172.050 755.400 ;
        RECT 205.950 756.600 208.050 757.050 ;
        RECT 220.950 756.600 223.050 756.900 ;
        RECT 205.950 755.400 223.050 756.600 ;
        RECT 205.950 754.950 208.050 755.400 ;
        RECT 220.950 754.800 223.050 755.400 ;
        RECT 232.950 756.600 235.050 757.050 ;
        RECT 244.950 756.600 247.050 756.900 ;
        RECT 262.950 756.600 265.050 757.050 ;
        RECT 232.950 755.400 265.050 756.600 ;
        RECT 232.950 754.950 235.050 755.400 ;
        RECT 244.950 754.800 247.050 755.400 ;
        RECT 262.950 754.950 265.050 755.400 ;
        RECT 355.950 756.450 358.050 756.900 ;
        RECT 364.950 756.450 367.050 756.900 ;
        RECT 355.950 755.250 367.050 756.450 ;
        RECT 355.950 754.800 358.050 755.250 ;
        RECT 364.950 754.800 367.050 755.250 ;
        RECT 370.950 756.450 373.050 756.900 ;
        RECT 385.950 756.450 388.050 756.900 ;
        RECT 370.950 755.250 388.050 756.450 ;
        RECT 370.950 754.800 373.050 755.250 ;
        RECT 385.950 754.800 388.050 755.250 ;
        RECT 421.950 756.600 424.050 756.900 ;
        RECT 430.800 756.600 432.900 757.050 ;
        RECT 421.950 755.400 432.900 756.600 ;
        RECT 421.950 754.800 424.050 755.400 ;
        RECT 430.800 754.950 432.900 755.400 ;
        RECT 433.950 756.600 436.050 757.050 ;
        RECT 442.950 756.600 445.050 756.900 ;
        RECT 433.950 755.400 445.050 756.600 ;
        RECT 433.950 754.950 436.050 755.400 ;
        RECT 442.950 754.800 445.050 755.400 ;
        RECT 472.950 756.600 475.050 756.900 ;
        RECT 496.950 756.600 499.050 756.900 ;
        RECT 472.950 755.400 499.050 756.600 ;
        RECT 472.950 754.800 475.050 755.400 ;
        RECT 496.950 754.800 499.050 755.400 ;
        RECT 535.950 756.450 538.050 756.900 ;
        RECT 547.950 756.450 550.050 756.900 ;
        RECT 535.950 755.250 550.050 756.450 ;
        RECT 535.950 754.800 538.050 755.250 ;
        RECT 547.950 754.800 550.050 755.250 ;
        RECT 559.950 756.450 562.050 756.900 ;
        RECT 565.950 756.450 568.050 756.900 ;
        RECT 559.950 755.250 568.050 756.450 ;
        RECT 602.400 755.400 607.050 757.050 ;
        RECT 559.950 754.800 562.050 755.250 ;
        RECT 565.950 754.800 568.050 755.250 ;
        RECT 603.000 754.950 607.050 755.400 ;
        RECT 613.950 756.450 616.050 756.900 ;
        RECT 619.950 756.450 622.050 756.900 ;
        RECT 613.950 755.250 622.050 756.450 ;
        RECT 613.950 754.800 616.050 755.250 ;
        RECT 619.950 754.800 622.050 755.250 ;
        RECT 625.950 756.450 628.050 756.900 ;
        RECT 634.950 756.450 637.050 756.900 ;
        RECT 625.950 755.250 637.050 756.450 ;
        RECT 625.950 754.800 628.050 755.250 ;
        RECT 634.950 754.800 637.050 755.250 ;
        RECT 649.950 756.600 652.050 756.900 ;
        RECT 673.950 756.600 676.050 756.900 ;
        RECT 649.950 755.400 676.050 756.600 ;
        RECT 649.950 754.800 652.050 755.400 ;
        RECT 673.950 754.800 676.050 755.400 ;
        RECT 685.950 756.450 688.050 756.900 ;
        RECT 694.950 756.450 697.050 756.900 ;
        RECT 685.950 755.250 697.050 756.450 ;
        RECT 701.400 756.600 702.600 758.400 ;
        RECT 721.950 756.600 724.050 756.900 ;
        RECT 737.400 756.600 738.600 760.950 ;
        RECT 754.950 759.600 757.050 760.050 ;
        RECT 874.950 759.600 877.050 760.050 ;
        RECT 893.400 759.600 894.600 761.400 ;
        RECT 925.950 760.950 928.050 761.400 ;
        RECT 754.950 758.400 777.600 759.600 ;
        RECT 754.950 757.950 757.050 758.400 ;
        RECT 739.950 756.600 742.050 756.900 ;
        RECT 701.400 755.400 724.050 756.600 ;
        RECT 685.950 754.800 688.050 755.250 ;
        RECT 694.950 754.800 697.050 755.250 ;
        RECT 721.950 754.800 724.050 755.400 ;
        RECT 725.400 755.400 742.050 756.600 ;
        RECT 106.950 753.600 109.050 754.050 ;
        RECT 148.950 753.600 151.050 754.050 ;
        RECT 106.950 752.400 151.050 753.600 ;
        RECT 106.950 751.950 109.050 752.400 ;
        RECT 148.950 751.950 151.050 752.400 ;
        RECT 364.950 753.600 367.050 754.050 ;
        RECT 391.950 753.600 394.050 754.050 ;
        RECT 364.950 752.400 394.050 753.600 ;
        RECT 364.950 751.950 367.050 752.400 ;
        RECT 391.950 751.950 394.050 752.400 ;
        RECT 583.950 753.600 586.050 754.050 ;
        RECT 592.950 753.600 595.050 754.050 ;
        RECT 583.950 752.400 595.050 753.600 ;
        RECT 583.950 751.950 586.050 752.400 ;
        RECT 592.950 751.950 595.050 752.400 ;
        RECT 601.950 753.600 604.050 754.050 ;
        RECT 670.950 753.600 673.050 754.050 ;
        RECT 601.950 752.400 673.050 753.600 ;
        RECT 601.950 751.950 604.050 752.400 ;
        RECT 670.950 751.950 673.050 752.400 ;
        RECT 715.950 753.600 718.050 754.050 ;
        RECT 725.400 753.600 726.600 755.400 ;
        RECT 739.950 754.800 742.050 755.400 ;
        RECT 763.950 756.600 766.050 756.900 ;
        RECT 772.950 756.600 775.050 757.050 ;
        RECT 763.950 755.400 775.050 756.600 ;
        RECT 776.400 756.600 777.600 758.400 ;
        RECT 874.950 758.400 894.600 759.600 ;
        RECT 941.400 759.600 942.600 764.400 ;
        RECT 1006.950 763.950 1009.050 766.050 ;
        RECT 1030.950 765.600 1033.050 766.050 ;
        RECT 1042.950 765.600 1045.050 765.900 ;
        RECT 1030.950 764.400 1045.050 765.600 ;
        RECT 1030.950 763.950 1033.050 764.400 ;
        RECT 955.950 762.600 958.050 763.200 ;
        RECT 964.950 762.600 967.050 763.050 ;
        RECT 955.950 761.400 967.050 762.600 ;
        RECT 955.950 761.100 958.050 761.400 ;
        RECT 964.950 760.950 967.050 761.400 ;
        RECT 973.950 762.750 976.050 763.200 ;
        RECT 982.950 762.750 985.050 763.200 ;
        RECT 973.950 761.550 985.050 762.750 ;
        RECT 973.950 761.100 976.050 761.550 ;
        RECT 982.950 761.100 985.050 761.550 ;
        RECT 1003.950 761.100 1006.050 763.200 ;
        RECT 1004.400 759.600 1005.600 761.100 ;
        RECT 941.400 758.400 954.600 759.600 ;
        RECT 874.950 757.950 877.050 758.400 ;
        RECT 781.950 756.600 784.050 757.050 ;
        RECT 776.400 755.400 784.050 756.600 ;
        RECT 763.950 754.800 766.050 755.400 ;
        RECT 772.950 754.950 775.050 755.400 ;
        RECT 781.950 754.950 784.050 755.400 ;
        RECT 790.950 756.450 793.050 756.900 ;
        RECT 796.950 756.450 799.050 756.900 ;
        RECT 790.950 755.250 799.050 756.450 ;
        RECT 790.950 754.800 793.050 755.250 ;
        RECT 796.950 754.800 799.050 755.250 ;
        RECT 820.950 756.600 823.050 757.050 ;
        RECT 832.950 756.600 835.050 756.900 ;
        RECT 820.950 755.400 835.050 756.600 ;
        RECT 820.950 754.950 823.050 755.400 ;
        RECT 832.950 754.800 835.050 755.400 ;
        RECT 838.950 754.800 841.050 756.900 ;
        RECT 844.950 756.600 847.050 757.050 ;
        RECT 862.950 756.600 865.050 756.900 ;
        RECT 877.950 756.600 880.050 757.050 ;
        RECT 953.400 756.900 954.600 758.400 ;
        RECT 989.400 758.400 1005.600 759.600 ;
        RECT 844.950 755.400 880.050 756.600 ;
        RECT 844.950 754.950 847.050 755.400 ;
        RECT 862.950 754.800 865.050 755.400 ;
        RECT 877.950 754.950 880.050 755.400 ;
        RECT 952.950 754.800 955.050 756.900 ;
        RECT 967.950 756.600 970.050 756.900 ;
        RECT 989.400 756.600 990.600 758.400 ;
        RECT 967.950 755.400 990.600 756.600 ;
        RECT 1007.400 756.600 1008.600 763.950 ;
        RECT 1042.950 763.800 1045.050 764.400 ;
        RECT 1009.950 762.750 1012.050 763.200 ;
        RECT 1018.950 762.750 1021.050 762.900 ;
        RECT 1009.950 761.550 1021.050 762.750 ;
        RECT 1009.950 761.100 1012.050 761.550 ;
        RECT 1018.950 760.800 1021.050 761.550 ;
        RECT 1012.950 756.600 1015.050 757.050 ;
        RECT 1007.400 755.400 1015.050 756.600 ;
        RECT 967.950 754.800 970.050 755.400 ;
        RECT 1012.950 754.950 1015.050 755.400 ;
        RECT 715.950 752.400 726.600 753.600 ;
        RECT 808.950 753.600 811.050 754.050 ;
        RECT 839.400 753.600 840.600 754.800 ;
        RECT 808.950 752.400 840.600 753.600 ;
        RECT 868.950 753.600 871.050 754.050 ;
        RECT 991.950 753.600 994.050 754.050 ;
        RECT 1006.800 753.600 1008.900 754.050 ;
        RECT 868.950 752.400 876.600 753.600 ;
        RECT 715.950 751.950 718.050 752.400 ;
        RECT 808.950 751.950 811.050 752.400 ;
        RECT 868.950 751.950 871.050 752.400 ;
        RECT 34.950 750.600 37.050 751.050 ;
        RECT 49.950 750.600 52.050 751.050 ;
        RECT 34.950 749.400 52.050 750.600 ;
        RECT 34.950 748.950 37.050 749.400 ;
        RECT 49.950 748.950 52.050 749.400 ;
        RECT 58.950 750.600 61.050 751.050 ;
        RECT 97.950 750.600 100.050 751.050 ;
        RECT 58.950 749.400 100.050 750.600 ;
        RECT 58.950 748.950 61.050 749.400 ;
        RECT 97.950 748.950 100.050 749.400 ;
        RECT 115.950 750.600 118.050 751.050 ;
        RECT 145.950 750.600 148.050 751.050 ;
        RECT 115.950 749.400 148.050 750.600 ;
        RECT 115.950 748.950 118.050 749.400 ;
        RECT 145.950 748.950 148.050 749.400 ;
        RECT 184.950 750.600 187.050 751.050 ;
        RECT 196.950 750.600 199.050 751.050 ;
        RECT 184.950 749.400 199.050 750.600 ;
        RECT 184.950 748.950 187.050 749.400 ;
        RECT 196.950 748.950 199.050 749.400 ;
        RECT 388.950 750.600 391.050 751.050 ;
        RECT 415.950 750.600 418.050 751.050 ;
        RECT 388.950 749.400 418.050 750.600 ;
        RECT 388.950 748.950 391.050 749.400 ;
        RECT 415.950 748.950 418.050 749.400 ;
        RECT 523.950 750.600 526.050 751.050 ;
        RECT 577.950 750.600 580.050 751.050 ;
        RECT 523.950 749.400 580.050 750.600 ;
        RECT 523.950 748.950 526.050 749.400 ;
        RECT 577.950 748.950 580.050 749.400 ;
        RECT 592.950 750.600 595.050 750.900 ;
        RECT 598.950 750.600 601.050 751.050 ;
        RECT 637.950 750.600 640.050 751.050 ;
        RECT 592.950 749.400 640.050 750.600 ;
        RECT 592.950 748.800 595.050 749.400 ;
        RECT 598.950 748.950 601.050 749.400 ;
        RECT 637.950 748.950 640.050 749.400 ;
        RECT 667.950 750.600 670.050 751.050 ;
        RECT 754.950 750.600 757.050 751.050 ;
        RECT 667.950 749.400 757.050 750.600 ;
        RECT 667.950 748.950 670.050 749.400 ;
        RECT 754.950 748.950 757.050 749.400 ;
        RECT 781.950 750.600 784.050 751.050 ;
        RECT 871.950 750.600 874.050 751.050 ;
        RECT 781.950 749.400 874.050 750.600 ;
        RECT 875.400 750.600 876.600 752.400 ;
        RECT 991.950 752.400 1008.900 753.600 ;
        RECT 991.950 751.950 994.050 752.400 ;
        RECT 1006.800 751.950 1008.900 752.400 ;
        RECT 1009.950 753.600 1012.050 754.050 ;
        RECT 1021.950 753.600 1024.050 754.050 ;
        RECT 1009.950 752.400 1024.050 753.600 ;
        RECT 1009.950 751.950 1012.050 752.400 ;
        RECT 1021.950 751.950 1024.050 752.400 ;
        RECT 1027.950 753.600 1030.050 754.050 ;
        RECT 1046.400 753.600 1047.600 766.950 ;
        RECT 1027.950 752.400 1047.600 753.600 ;
        RECT 1027.950 751.950 1030.050 752.400 ;
        RECT 886.950 750.600 889.050 751.050 ;
        RECT 910.950 750.600 913.050 751.050 ;
        RECT 875.400 749.400 913.050 750.600 ;
        RECT 781.950 748.950 784.050 749.400 ;
        RECT 871.950 748.950 874.050 749.400 ;
        RECT 886.950 748.950 889.050 749.400 ;
        RECT 910.950 748.950 913.050 749.400 ;
        RECT 925.950 750.600 928.050 751.050 ;
        RECT 931.950 750.600 934.050 751.050 ;
        RECT 925.950 749.400 934.050 750.600 ;
        RECT 925.950 748.950 928.050 749.400 ;
        RECT 931.950 748.950 934.050 749.400 ;
        RECT 940.950 750.600 943.050 751.050 ;
        RECT 958.950 750.600 961.050 751.050 ;
        RECT 985.950 750.600 988.050 751.050 ;
        RECT 940.950 749.400 988.050 750.600 ;
        RECT 940.950 748.950 943.050 749.400 ;
        RECT 958.950 748.950 961.050 749.400 ;
        RECT 985.950 748.950 988.050 749.400 ;
        RECT 1015.950 750.600 1020.000 751.050 ;
        RECT 1015.950 748.950 1020.600 750.600 ;
        RECT 232.950 747.600 235.050 748.050 ;
        RECT 250.950 747.600 253.050 748.050 ;
        RECT 286.950 747.600 289.050 748.050 ;
        RECT 232.950 746.400 289.050 747.600 ;
        RECT 232.950 745.950 235.050 746.400 ;
        RECT 250.950 745.950 253.050 746.400 ;
        RECT 286.950 745.950 289.050 746.400 ;
        RECT 352.950 747.600 355.050 748.050 ;
        RECT 385.950 747.600 388.050 748.050 ;
        RECT 448.950 747.600 451.050 748.050 ;
        RECT 481.950 747.600 484.050 748.050 ;
        RECT 352.950 746.400 484.050 747.600 ;
        RECT 352.950 745.950 355.050 746.400 ;
        RECT 385.950 745.950 388.050 746.400 ;
        RECT 448.950 745.950 451.050 746.400 ;
        RECT 481.950 745.950 484.050 746.400 ;
        RECT 505.950 747.600 508.050 748.050 ;
        RECT 601.950 747.600 604.050 748.050 ;
        RECT 505.950 746.400 604.050 747.600 ;
        RECT 505.950 745.950 508.050 746.400 ;
        RECT 601.950 745.950 604.050 746.400 ;
        RECT 661.950 747.600 664.050 748.050 ;
        RECT 712.950 747.600 715.050 748.050 ;
        RECT 661.950 746.400 715.050 747.600 ;
        RECT 661.950 745.950 664.050 746.400 ;
        RECT 712.950 745.950 715.050 746.400 ;
        RECT 799.950 747.600 802.050 748.050 ;
        RECT 823.950 747.600 826.050 748.050 ;
        RECT 799.950 746.400 826.050 747.600 ;
        RECT 799.950 745.950 802.050 746.400 ;
        RECT 823.950 745.950 826.050 746.400 ;
        RECT 865.950 747.600 868.050 748.050 ;
        RECT 895.950 747.600 898.050 748.050 ;
        RECT 865.950 746.400 898.050 747.600 ;
        RECT 865.950 745.950 868.050 746.400 ;
        RECT 895.950 745.950 898.050 746.400 ;
        RECT 928.950 747.600 931.050 748.050 ;
        RECT 967.950 747.600 970.050 748.050 ;
        RECT 928.950 746.400 970.050 747.600 ;
        RECT 928.950 745.950 931.050 746.400 ;
        RECT 967.950 745.950 970.050 746.400 ;
        RECT 1006.950 747.600 1009.050 748.050 ;
        RECT 1012.950 747.600 1015.050 748.050 ;
        RECT 1006.950 746.400 1015.050 747.600 ;
        RECT 1019.400 747.600 1020.600 748.950 ;
        RECT 1036.950 747.600 1039.050 748.050 ;
        RECT 1019.400 746.400 1039.050 747.600 ;
        RECT 1006.950 745.950 1009.050 746.400 ;
        RECT 1012.950 745.950 1015.050 746.400 ;
        RECT 1036.950 745.950 1039.050 746.400 ;
        RECT 151.950 744.600 154.050 745.050 ;
        RECT 190.950 744.600 193.050 745.050 ;
        RECT 151.950 743.400 193.050 744.600 ;
        RECT 151.950 742.950 154.050 743.400 ;
        RECT 190.950 742.950 193.050 743.400 ;
        RECT 208.950 744.600 211.050 745.050 ;
        RECT 223.950 744.600 226.050 745.050 ;
        RECT 208.950 743.400 226.050 744.600 ;
        RECT 208.950 742.950 211.050 743.400 ;
        RECT 223.950 742.950 226.050 743.400 ;
        RECT 343.950 744.600 346.050 745.050 ;
        RECT 367.950 744.600 370.050 745.050 ;
        RECT 343.950 743.400 370.050 744.600 ;
        RECT 343.950 742.950 346.050 743.400 ;
        RECT 367.950 742.950 370.050 743.400 ;
        RECT 400.950 744.600 403.050 745.050 ;
        RECT 433.950 744.600 436.050 745.050 ;
        RECT 703.950 744.600 706.050 745.050 ;
        RECT 400.950 743.400 436.050 744.600 ;
        RECT 400.950 742.950 403.050 743.400 ;
        RECT 433.950 742.950 436.050 743.400 ;
        RECT 605.400 743.400 706.050 744.600 ;
        RECT 191.400 741.600 192.600 742.950 ;
        RECT 220.950 741.600 223.050 742.050 ;
        RECT 191.400 740.400 223.050 741.600 ;
        RECT 220.950 739.950 223.050 740.400 ;
        RECT 226.950 741.600 229.050 742.050 ;
        RECT 352.950 741.600 355.050 742.050 ;
        RECT 388.950 741.600 391.050 742.050 ;
        RECT 226.950 740.400 276.600 741.600 ;
        RECT 226.950 739.950 229.050 740.400 ;
        RECT 112.950 738.600 115.050 739.050 ;
        RECT 181.950 738.600 184.050 739.050 ;
        RECT 112.950 737.400 184.050 738.600 ;
        RECT 275.400 738.600 276.600 740.400 ;
        RECT 352.950 740.400 391.050 741.600 ;
        RECT 434.400 741.600 435.600 742.950 ;
        RECT 605.400 742.050 606.600 743.400 ;
        RECT 703.950 742.950 706.050 743.400 ;
        RECT 721.950 744.600 724.050 745.050 ;
        RECT 736.950 744.600 739.050 745.050 ;
        RECT 721.950 743.400 739.050 744.600 ;
        RECT 721.950 742.950 724.050 743.400 ;
        RECT 736.950 742.950 739.050 743.400 ;
        RECT 784.950 744.600 787.050 745.050 ;
        RECT 829.950 744.600 832.050 745.050 ;
        RECT 784.950 743.400 832.050 744.600 ;
        RECT 784.950 742.950 787.050 743.400 ;
        RECT 829.950 742.950 832.050 743.400 ;
        RECT 841.950 744.600 844.050 745.050 ;
        RECT 850.950 744.600 853.050 745.050 ;
        RECT 841.950 743.400 853.050 744.600 ;
        RECT 841.950 742.950 844.050 743.400 ;
        RECT 850.950 742.950 853.050 743.400 ;
        RECT 859.950 744.600 862.050 745.050 ;
        RECT 874.950 744.600 877.050 745.050 ;
        RECT 859.950 743.400 877.050 744.600 ;
        RECT 859.950 742.950 862.050 743.400 ;
        RECT 874.950 742.950 877.050 743.400 ;
        RECT 898.950 744.600 901.050 745.050 ;
        RECT 910.950 744.600 913.050 745.050 ;
        RECT 898.950 743.400 913.050 744.600 ;
        RECT 898.950 742.950 901.050 743.400 ;
        RECT 910.950 742.950 913.050 743.400 ;
        RECT 925.950 744.600 928.050 745.050 ;
        RECT 982.950 744.600 985.050 745.050 ;
        RECT 925.950 743.400 985.050 744.600 ;
        RECT 925.950 742.950 928.050 743.400 ;
        RECT 982.950 742.950 985.050 743.400 ;
        RECT 517.950 741.600 520.050 742.050 ;
        RECT 434.400 740.400 520.050 741.600 ;
        RECT 352.950 739.950 355.050 740.400 ;
        RECT 388.950 739.950 391.050 740.400 ;
        RECT 517.950 739.950 520.050 740.400 ;
        RECT 532.950 741.600 535.050 742.050 ;
        RECT 550.950 741.600 553.050 742.050 ;
        RECT 532.950 740.400 553.050 741.600 ;
        RECT 532.950 739.950 535.050 740.400 ;
        RECT 550.950 739.950 553.050 740.400 ;
        RECT 571.950 741.600 574.050 742.050 ;
        RECT 580.950 741.600 583.050 742.050 ;
        RECT 571.950 740.400 583.050 741.600 ;
        RECT 571.950 739.950 574.050 740.400 ;
        RECT 580.950 739.950 583.050 740.400 ;
        RECT 601.950 740.400 606.600 742.050 ;
        RECT 607.950 741.600 610.050 742.050 ;
        RECT 661.950 741.600 664.050 742.050 ;
        RECT 607.950 740.400 664.050 741.600 ;
        RECT 601.950 739.950 606.000 740.400 ;
        RECT 607.950 739.950 610.050 740.400 ;
        RECT 661.950 739.950 664.050 740.400 ;
        RECT 670.950 741.600 673.050 742.050 ;
        RECT 739.950 741.600 742.050 742.050 ;
        RECT 670.950 740.400 742.050 741.600 ;
        RECT 670.950 739.950 673.050 740.400 ;
        RECT 739.950 739.950 742.050 740.400 ;
        RECT 853.950 741.600 856.050 742.050 ;
        RECT 985.950 741.600 988.050 742.050 ;
        RECT 1024.950 741.600 1027.050 742.050 ;
        RECT 853.950 740.400 1027.050 741.600 ;
        RECT 853.950 739.950 856.050 740.400 ;
        RECT 985.950 739.950 988.050 740.400 ;
        RECT 1024.950 739.950 1027.050 740.400 ;
        RECT 292.950 738.600 295.050 739.050 ;
        RECT 275.400 737.400 295.050 738.600 ;
        RECT 112.950 736.950 115.050 737.400 ;
        RECT 181.950 736.950 184.050 737.400 ;
        RECT 292.950 736.950 295.050 737.400 ;
        RECT 553.950 738.600 556.050 739.050 ;
        RECT 571.950 738.600 574.050 738.900 ;
        RECT 643.950 738.600 646.050 739.050 ;
        RECT 553.950 737.400 646.050 738.600 ;
        RECT 553.950 736.950 556.050 737.400 ;
        RECT 571.950 736.800 574.050 737.400 ;
        RECT 643.950 736.950 646.050 737.400 ;
        RECT 664.950 738.600 667.050 739.050 ;
        RECT 727.950 738.600 730.050 739.050 ;
        RECT 745.950 738.600 748.050 739.050 ;
        RECT 664.950 737.400 748.050 738.600 ;
        RECT 664.950 736.950 667.050 737.400 ;
        RECT 727.950 736.950 730.050 737.400 ;
        RECT 745.950 736.950 748.050 737.400 ;
        RECT 766.950 738.600 769.050 739.050 ;
        RECT 790.950 738.600 793.050 739.050 ;
        RECT 766.950 737.400 793.050 738.600 ;
        RECT 766.950 736.950 769.050 737.400 ;
        RECT 790.950 736.950 793.050 737.400 ;
        RECT 829.950 738.600 832.050 739.050 ;
        RECT 844.950 738.600 847.050 739.050 ;
        RECT 829.950 737.400 847.050 738.600 ;
        RECT 829.950 736.950 832.050 737.400 ;
        RECT 844.950 736.950 847.050 737.400 ;
        RECT 862.950 738.600 865.050 739.050 ;
        RECT 925.950 738.600 928.050 739.050 ;
        RECT 862.950 737.400 928.050 738.600 ;
        RECT 862.950 736.950 865.050 737.400 ;
        RECT 925.950 736.950 928.050 737.400 ;
        RECT 946.950 738.600 949.050 739.050 ;
        RECT 976.950 738.600 979.050 739.050 ;
        RECT 946.950 737.400 979.050 738.600 ;
        RECT 946.950 736.950 949.050 737.400 ;
        RECT 976.950 736.950 979.050 737.400 ;
        RECT 217.950 735.600 220.050 736.050 ;
        RECT 262.950 735.600 265.050 736.050 ;
        RECT 217.950 734.400 265.050 735.600 ;
        RECT 217.950 733.950 220.050 734.400 ;
        RECT 262.950 733.950 265.050 734.400 ;
        RECT 340.950 735.600 343.050 736.050 ;
        RECT 349.950 735.600 352.050 736.050 ;
        RECT 340.950 734.400 352.050 735.600 ;
        RECT 340.950 733.950 343.050 734.400 ;
        RECT 349.950 733.950 352.050 734.400 ;
        RECT 409.950 735.600 412.050 736.050 ;
        RECT 436.950 735.600 439.050 736.050 ;
        RECT 409.950 734.400 439.050 735.600 ;
        RECT 409.950 733.950 412.050 734.400 ;
        RECT 436.950 733.950 439.050 734.400 ;
        RECT 454.950 735.600 457.050 736.050 ;
        RECT 487.950 735.600 490.050 736.050 ;
        RECT 454.950 734.400 490.050 735.600 ;
        RECT 454.950 733.950 457.050 734.400 ;
        RECT 487.950 733.950 490.050 734.400 ;
        RECT 565.950 735.600 568.050 736.050 ;
        RECT 586.950 735.600 589.050 736.050 ;
        RECT 565.950 734.400 589.050 735.600 ;
        RECT 565.950 733.950 568.050 734.400 ;
        RECT 586.950 733.950 589.050 734.400 ;
        RECT 703.950 735.600 706.050 736.050 ;
        RECT 757.950 735.600 760.050 736.050 ;
        RECT 703.950 734.400 760.050 735.600 ;
        RECT 703.950 733.950 706.050 734.400 ;
        RECT 757.950 733.950 760.050 734.400 ;
        RECT 847.950 735.600 850.050 736.050 ;
        RECT 853.950 735.600 856.050 736.050 ;
        RECT 847.950 734.400 856.050 735.600 ;
        RECT 847.950 733.950 850.050 734.400 ;
        RECT 853.950 733.950 856.050 734.400 ;
        RECT 874.950 735.600 877.050 736.050 ;
        RECT 883.950 735.600 886.050 736.050 ;
        RECT 874.950 734.400 886.050 735.600 ;
        RECT 874.950 733.950 877.050 734.400 ;
        RECT 883.950 733.950 886.050 734.400 ;
        RECT 901.950 735.600 904.050 736.050 ;
        RECT 907.950 735.600 910.050 736.050 ;
        RECT 901.950 734.400 910.050 735.600 ;
        RECT 901.950 733.950 904.050 734.400 ;
        RECT 907.950 733.950 910.050 734.400 ;
        RECT 949.950 735.600 952.050 736.050 ;
        RECT 979.950 735.600 982.050 736.050 ;
        RECT 949.950 734.400 982.050 735.600 ;
        RECT 949.950 733.950 952.050 734.400 ;
        RECT 979.950 733.950 982.050 734.400 ;
        RECT 136.950 730.950 139.050 733.050 ;
        RECT 280.950 732.600 283.050 733.050 ;
        RECT 286.950 732.600 289.050 733.050 ;
        RECT 280.950 731.400 289.050 732.600 ;
        RECT 280.950 730.950 283.050 731.400 ;
        RECT 286.950 730.950 289.050 731.400 ;
        RECT 361.950 732.600 364.050 733.050 ;
        RECT 379.950 732.600 382.050 733.050 ;
        RECT 361.950 731.400 382.050 732.600 ;
        RECT 361.950 730.950 364.050 731.400 ;
        RECT 379.950 730.950 382.050 731.400 ;
        RECT 496.950 732.600 499.050 733.050 ;
        RECT 514.950 732.600 517.050 733.050 ;
        RECT 532.950 732.600 535.050 733.050 ;
        RECT 496.950 731.400 510.600 732.600 ;
        RECT 496.950 730.950 499.050 731.400 ;
        RECT 40.950 729.600 43.050 730.200 ;
        RECT 64.950 729.600 67.050 730.200 ;
        RECT 40.950 728.400 67.050 729.600 ;
        RECT 40.950 728.100 43.050 728.400 ;
        RECT 64.950 728.100 67.050 728.400 ;
        RECT 124.950 729.750 127.050 730.200 ;
        RECT 133.950 729.750 136.050 730.200 ;
        RECT 124.950 728.550 136.050 729.750 ;
        RECT 124.950 728.100 127.050 728.550 ;
        RECT 133.950 728.100 136.050 728.550 ;
        RECT 137.400 723.900 138.600 730.950 ;
        RECT 139.950 729.750 142.050 730.200 ;
        RECT 145.950 729.750 148.050 730.200 ;
        RECT 139.950 728.550 148.050 729.750 ;
        RECT 139.950 728.100 142.050 728.550 ;
        RECT 145.950 728.100 148.050 728.550 ;
        RECT 163.950 728.100 166.050 730.200 ;
        RECT 136.950 721.800 139.050 723.900 ;
        RECT 164.400 721.050 165.600 728.100 ;
        RECT 169.950 727.950 172.050 730.050 ;
        RECT 220.950 729.750 223.050 730.200 ;
        RECT 256.950 729.750 259.050 730.200 ;
        RECT 220.950 728.550 259.050 729.750 ;
        RECT 220.950 728.100 223.050 728.550 ;
        RECT 256.950 728.100 259.050 728.550 ;
        RECT 274.950 729.600 277.050 730.050 ;
        RECT 304.950 729.600 307.050 730.200 ;
        RECT 319.950 729.600 322.050 730.050 ;
        RECT 274.950 728.400 322.050 729.600 ;
        RECT 274.950 727.950 277.050 728.400 ;
        RECT 304.950 728.100 307.050 728.400 ;
        RECT 319.950 727.950 322.050 728.400 ;
        RECT 337.950 729.750 340.050 730.200 ;
        RECT 346.950 729.750 349.050 730.200 ;
        RECT 337.950 728.550 349.050 729.750 ;
        RECT 337.950 728.100 340.050 728.550 ;
        RECT 346.950 728.100 349.050 728.550 ;
        RECT 170.400 723.600 171.600 727.950 ;
        RECT 196.950 726.450 199.050 726.900 ;
        RECT 217.950 726.450 220.050 726.900 ;
        RECT 196.950 725.250 220.050 726.450 ;
        RECT 358.950 726.600 361.050 730.050 ;
        RECT 364.950 729.600 367.050 730.050 ;
        RECT 376.950 729.600 379.050 730.200 ;
        RECT 364.950 728.400 379.050 729.600 ;
        RECT 364.950 727.950 367.050 728.400 ;
        RECT 376.950 728.100 379.050 728.400 ;
        RECT 388.950 729.600 391.050 730.050 ;
        RECT 421.950 729.600 424.050 730.200 ;
        RECT 388.950 728.400 424.050 729.600 ;
        RECT 388.950 727.950 391.050 728.400 ;
        RECT 421.950 728.100 424.050 728.400 ;
        RECT 436.950 729.750 439.050 730.200 ;
        RECT 445.950 729.750 448.050 730.200 ;
        RECT 436.950 728.550 448.050 729.750 ;
        RECT 436.950 728.100 439.050 728.550 ;
        RECT 445.950 728.100 448.050 728.550 ;
        RECT 451.950 729.600 454.050 730.050 ;
        RECT 460.950 729.600 463.050 730.050 ;
        RECT 451.950 728.400 463.050 729.600 ;
        RECT 451.950 727.950 454.050 728.400 ;
        RECT 460.950 727.950 463.050 728.400 ;
        RECT 466.950 728.100 469.050 730.200 ;
        RECT 478.950 729.600 481.050 730.050 ;
        RECT 493.950 729.600 496.050 730.200 ;
        RECT 502.950 729.600 505.050 730.050 ;
        RECT 478.950 728.400 505.050 729.600 ;
        RECT 467.400 726.600 468.600 728.100 ;
        RECT 478.950 727.950 481.050 728.400 ;
        RECT 493.950 728.100 496.050 728.400 ;
        RECT 502.950 727.950 505.050 728.400 ;
        RECT 484.950 726.600 487.050 727.050 ;
        RECT 358.950 726.000 369.600 726.600 ;
        RECT 359.400 725.400 369.600 726.000 ;
        RECT 467.400 725.400 487.050 726.600 ;
        RECT 196.950 724.800 199.050 725.250 ;
        RECT 217.950 724.800 220.050 725.250 ;
        RECT 170.400 723.000 177.600 723.600 ;
        RECT 259.950 723.450 262.050 723.900 ;
        RECT 268.950 723.450 271.050 723.900 ;
        RECT 170.400 722.400 178.050 723.000 ;
        RECT 73.950 720.600 76.050 721.050 ;
        RECT 91.950 720.600 94.050 721.050 ;
        RECT 73.950 719.400 94.050 720.600 ;
        RECT 73.950 718.950 76.050 719.400 ;
        RECT 91.950 718.950 94.050 719.400 ;
        RECT 97.950 720.600 100.050 721.050 ;
        RECT 106.950 720.600 109.050 721.050 ;
        RECT 112.950 720.600 115.050 721.050 ;
        RECT 97.950 719.400 115.050 720.600 ;
        RECT 97.950 718.950 100.050 719.400 ;
        RECT 106.950 718.950 109.050 719.400 ;
        RECT 112.950 718.950 115.050 719.400 ;
        RECT 163.950 718.950 166.050 721.050 ;
        RECT 175.950 718.950 178.050 722.400 ;
        RECT 259.950 722.250 271.050 723.450 ;
        RECT 259.950 721.800 262.050 722.250 ;
        RECT 268.950 721.800 271.050 722.250 ;
        RECT 328.950 723.600 331.050 723.900 ;
        RECT 349.950 723.600 352.050 723.900 ;
        RECT 328.950 722.400 352.050 723.600 ;
        RECT 328.950 721.800 331.050 722.400 ;
        RECT 349.950 721.800 352.050 722.400 ;
        RECT 355.950 723.450 358.050 723.900 ;
        RECT 364.950 723.450 367.050 723.900 ;
        RECT 355.950 722.250 367.050 723.450 ;
        RECT 368.400 723.600 369.600 725.400 ;
        RECT 484.950 724.950 487.050 725.400 ;
        RECT 418.950 723.600 421.050 723.900 ;
        RECT 368.400 722.400 421.050 723.600 ;
        RECT 355.950 721.800 358.050 722.250 ;
        RECT 364.950 721.800 367.050 722.250 ;
        RECT 418.950 721.800 421.050 722.400 ;
        RECT 460.950 723.450 463.050 723.900 ;
        RECT 469.950 723.450 472.050 723.900 ;
        RECT 460.950 722.250 472.050 723.450 ;
        RECT 460.950 721.800 463.050 722.250 ;
        RECT 469.950 721.800 472.050 722.250 ;
        RECT 490.950 723.450 493.050 723.900 ;
        RECT 505.950 723.450 508.050 723.900 ;
        RECT 490.950 722.250 508.050 723.450 ;
        RECT 509.400 723.600 510.600 731.400 ;
        RECT 514.950 731.400 535.050 732.600 ;
        RECT 514.950 730.950 517.050 731.400 ;
        RECT 532.950 730.950 535.050 731.400 ;
        RECT 541.950 732.600 544.050 733.050 ;
        RECT 616.950 732.600 619.050 733.050 ;
        RECT 541.950 731.400 619.050 732.600 ;
        RECT 541.950 730.950 544.050 731.400 ;
        RECT 616.950 730.950 619.050 731.400 ;
        RECT 643.950 732.600 646.050 733.200 ;
        RECT 685.950 732.600 688.050 733.050 ;
        RECT 643.950 731.400 688.050 732.600 ;
        RECT 643.950 731.100 646.050 731.400 ;
        RECT 685.950 730.950 688.050 731.400 ;
        RECT 700.950 732.600 703.050 733.050 ;
        RECT 721.950 732.600 724.050 733.050 ;
        RECT 700.950 731.400 724.050 732.600 ;
        RECT 700.950 730.950 703.050 731.400 ;
        RECT 721.950 730.950 724.050 731.400 ;
        RECT 742.950 732.600 745.050 733.050 ;
        RECT 763.950 732.600 766.050 733.050 ;
        RECT 742.950 731.400 766.050 732.600 ;
        RECT 742.950 730.950 745.050 731.400 ;
        RECT 763.950 730.950 766.050 731.400 ;
        RECT 973.950 732.600 976.050 733.050 ;
        RECT 979.950 732.600 982.050 732.900 ;
        RECT 973.950 731.400 982.050 732.600 ;
        RECT 973.950 730.950 976.050 731.400 ;
        RECT 979.950 730.800 982.050 731.400 ;
        RECT 994.950 732.600 997.050 733.050 ;
        RECT 1030.950 732.600 1033.050 733.050 ;
        RECT 994.950 731.400 1033.050 732.600 ;
        RECT 994.950 730.950 997.050 731.400 ;
        RECT 1030.950 730.950 1033.050 731.400 ;
        RECT 520.950 729.750 523.050 730.200 ;
        RECT 526.950 729.750 529.050 730.200 ;
        RECT 520.950 728.550 529.050 729.750 ;
        RECT 520.950 728.100 523.050 728.550 ;
        RECT 526.950 728.100 529.050 728.550 ;
        RECT 544.950 729.600 547.050 730.200 ;
        RECT 601.950 729.600 604.050 730.050 ;
        RECT 544.950 728.400 604.050 729.600 ;
        RECT 544.950 728.100 547.050 728.400 ;
        RECT 601.950 727.950 604.050 728.400 ;
        RECT 619.950 728.100 622.050 730.200 ;
        RECT 625.950 729.600 628.050 730.050 ;
        RECT 640.950 729.600 643.050 730.050 ;
        RECT 646.950 729.600 649.050 730.200 ;
        RECT 625.950 728.400 643.050 729.600 ;
        RECT 620.400 726.600 621.600 728.100 ;
        RECT 625.950 727.950 628.050 728.400 ;
        RECT 640.950 727.950 643.050 728.400 ;
        RECT 644.400 728.400 649.050 729.600 ;
        RECT 644.400 726.600 645.600 728.400 ;
        RECT 646.950 728.100 649.050 728.400 ;
        RECT 673.950 729.600 676.050 730.200 ;
        RECT 694.950 729.600 697.050 730.200 ;
        RECT 673.950 728.400 697.050 729.600 ;
        RECT 673.950 728.100 676.050 728.400 ;
        RECT 694.950 728.100 697.050 728.400 ;
        RECT 739.950 729.600 742.050 730.050 ;
        RECT 757.950 729.600 760.050 730.050 ;
        RECT 739.950 728.400 760.050 729.600 ;
        RECT 739.950 727.950 742.050 728.400 ;
        RECT 757.950 727.950 760.050 728.400 ;
        RECT 772.950 729.750 775.050 730.200 ;
        RECT 784.950 729.750 787.050 730.200 ;
        RECT 772.950 728.550 787.050 729.750 ;
        RECT 772.950 728.100 775.050 728.550 ;
        RECT 784.950 728.100 787.050 728.550 ;
        RECT 793.950 729.600 796.050 730.050 ;
        RECT 811.950 729.750 814.050 730.200 ;
        RECT 823.950 729.750 826.050 730.200 ;
        RECT 811.950 729.600 826.050 729.750 ;
        RECT 793.950 728.550 826.050 729.600 ;
        RECT 793.950 728.400 814.050 728.550 ;
        RECT 793.950 727.950 796.050 728.400 ;
        RECT 811.950 728.100 814.050 728.400 ;
        RECT 823.950 728.100 826.050 728.550 ;
        RECT 829.950 729.600 832.050 730.200 ;
        RECT 838.950 729.600 841.050 730.050 ;
        RECT 829.950 728.400 841.050 729.600 ;
        RECT 829.950 728.100 832.050 728.400 ;
        RECT 838.950 727.950 841.050 728.400 ;
        RECT 847.950 728.100 850.050 730.200 ;
        RECT 620.400 725.400 645.600 726.600 ;
        RECT 517.950 723.600 520.050 723.900 ;
        RECT 509.400 722.400 520.050 723.600 ;
        RECT 490.950 721.800 493.050 722.250 ;
        RECT 505.950 721.800 508.050 722.250 ;
        RECT 517.950 721.800 520.050 722.400 ;
        RECT 556.950 723.600 559.050 724.050 ;
        RECT 568.950 723.600 571.050 723.900 ;
        RECT 556.950 722.400 571.050 723.600 ;
        RECT 556.950 721.950 559.050 722.400 ;
        RECT 568.950 721.800 571.050 722.400 ;
        RECT 583.950 723.450 586.050 723.900 ;
        RECT 589.950 723.450 592.050 723.900 ;
        RECT 583.950 722.250 592.050 723.450 ;
        RECT 583.950 721.800 586.050 722.250 ;
        RECT 589.950 721.800 592.050 722.250 ;
        RECT 595.950 723.450 598.050 723.900 ;
        RECT 604.950 723.450 607.050 723.900 ;
        RECT 595.950 722.250 607.050 723.450 ;
        RECT 595.950 721.800 598.050 722.250 ;
        RECT 604.950 721.800 607.050 722.250 ;
        RECT 634.950 723.600 637.050 724.050 ;
        RECT 649.950 723.600 652.050 723.900 ;
        RECT 634.950 722.400 652.050 723.600 ;
        RECT 634.950 721.950 637.050 722.400 ;
        RECT 649.950 721.800 652.050 722.400 ;
        RECT 670.950 723.600 673.050 723.900 ;
        RECT 709.950 723.600 712.050 724.050 ;
        RECT 670.950 722.400 712.050 723.600 ;
        RECT 670.950 721.800 673.050 722.400 ;
        RECT 709.950 721.950 712.050 722.400 ;
        RECT 718.950 723.450 721.050 723.900 ;
        RECT 736.800 723.450 738.900 723.900 ;
        RECT 718.950 722.250 738.900 723.450 ;
        RECT 718.950 721.800 721.050 722.250 ;
        RECT 736.800 721.800 738.900 722.250 ;
        RECT 739.950 723.450 742.050 723.900 ;
        RECT 745.950 723.450 748.050 723.900 ;
        RECT 739.950 722.250 748.050 723.450 ;
        RECT 739.950 721.800 742.050 722.250 ;
        RECT 745.950 721.800 748.050 722.250 ;
        RECT 775.950 723.450 778.050 723.900 ;
        RECT 805.950 723.450 808.050 723.900 ;
        RECT 775.950 722.250 808.050 723.450 ;
        RECT 775.950 721.800 778.050 722.250 ;
        RECT 805.950 721.800 808.050 722.250 ;
        RECT 848.400 721.050 849.600 728.100 ;
        RECT 892.950 727.950 895.050 730.050 ;
        RECT 903.000 729.600 907.050 730.050 ;
        RECT 902.400 727.950 907.050 729.600 ;
        RECT 916.950 729.600 919.050 730.050 ;
        RECT 937.950 729.600 940.050 730.050 ;
        RECT 916.950 728.400 940.050 729.600 ;
        RECT 916.950 727.950 919.050 728.400 ;
        RECT 937.950 727.950 940.050 728.400 ;
        RECT 970.950 727.950 973.050 730.050 ;
        RECT 982.950 729.600 985.050 729.900 ;
        RECT 988.950 729.600 991.050 730.050 ;
        RECT 982.950 728.400 991.050 729.600 ;
        RECT 861.000 726.600 865.050 727.050 ;
        RECT 860.400 724.950 865.050 726.600 ;
        RECT 850.950 723.600 853.050 723.900 ;
        RECT 860.400 723.600 861.600 724.950 ;
        RECT 893.400 724.050 894.600 727.950 ;
        RECT 850.950 722.400 861.600 723.600 ;
        RECT 850.950 721.800 853.050 722.400 ;
        RECT 892.950 721.950 895.050 724.050 ;
        RECT 898.950 723.600 901.050 723.900 ;
        RECT 902.400 723.600 903.600 727.950 ;
        RECT 898.950 722.400 903.600 723.600 ;
        RECT 940.950 723.450 943.050 723.900 ;
        RECT 946.950 723.450 949.050 723.900 ;
        RECT 898.950 721.800 901.050 722.400 ;
        RECT 940.950 722.250 949.050 723.450 ;
        RECT 940.950 721.800 943.050 722.250 ;
        RECT 946.950 721.800 949.050 722.250 ;
        RECT 952.950 723.600 955.050 723.900 ;
        RECT 971.400 723.600 972.600 727.950 ;
        RECT 982.950 727.800 985.050 728.400 ;
        RECT 988.950 727.950 991.050 728.400 ;
        RECT 997.950 728.100 1000.050 730.200 ;
        RECT 1003.950 729.600 1006.050 730.050 ;
        RECT 1033.950 729.600 1036.050 730.050 ;
        RECT 1003.950 728.400 1036.050 729.600 ;
        RECT 952.950 722.400 972.600 723.600 ;
        RECT 973.950 723.600 976.050 723.900 ;
        RECT 998.400 723.600 999.600 728.100 ;
        RECT 1003.950 727.950 1006.050 728.400 ;
        RECT 1033.950 727.950 1036.050 728.400 ;
        RECT 973.950 722.400 999.600 723.600 ;
        RECT 952.950 721.800 955.050 722.400 ;
        RECT 973.950 721.800 976.050 722.400 ;
        RECT 253.950 720.600 256.050 721.050 ;
        RECT 271.950 720.600 274.050 721.050 ;
        RECT 283.950 720.600 286.050 721.050 ;
        RECT 253.950 719.400 286.050 720.600 ;
        RECT 253.950 718.950 256.050 719.400 ;
        RECT 271.950 718.950 274.050 719.400 ;
        RECT 283.950 718.950 286.050 719.400 ;
        RECT 379.950 720.600 382.050 721.050 ;
        RECT 400.950 720.600 403.050 721.050 ;
        RECT 379.950 719.400 403.050 720.600 ;
        RECT 379.950 718.950 382.050 719.400 ;
        RECT 400.950 718.950 403.050 719.400 ;
        RECT 502.950 720.600 505.050 721.050 ;
        RECT 541.950 720.600 544.050 721.050 ;
        RECT 502.950 719.400 544.050 720.600 ;
        RECT 502.950 718.950 505.050 719.400 ;
        RECT 541.950 718.950 544.050 719.400 ;
        RECT 718.950 720.600 721.050 720.750 ;
        RECT 775.950 720.600 778.050 721.050 ;
        RECT 718.950 719.400 778.050 720.600 ;
        RECT 718.950 718.650 721.050 719.400 ;
        RECT 775.950 718.950 778.050 719.400 ;
        RECT 790.950 720.600 793.050 721.050 ;
        RECT 802.950 720.600 805.050 721.050 ;
        RECT 790.950 719.400 805.050 720.600 ;
        RECT 790.950 718.950 793.050 719.400 ;
        RECT 802.950 718.950 805.050 719.400 ;
        RECT 814.950 720.600 817.050 721.050 ;
        RECT 847.950 720.600 850.050 721.050 ;
        RECT 814.950 719.400 850.050 720.600 ;
        RECT 814.950 718.950 817.050 719.400 ;
        RECT 847.950 718.950 850.050 719.400 ;
        RECT 865.950 720.600 868.050 721.050 ;
        RECT 871.950 720.600 874.050 721.050 ;
        RECT 865.950 719.400 874.050 720.600 ;
        RECT 865.950 718.950 868.050 719.400 ;
        RECT 871.950 718.950 874.050 719.400 ;
        RECT 919.950 720.600 922.050 721.050 ;
        RECT 928.950 720.600 931.050 721.050 ;
        RECT 919.950 719.400 931.050 720.600 ;
        RECT 919.950 718.950 922.050 719.400 ;
        RECT 928.950 718.950 931.050 719.400 ;
        RECT 994.950 720.600 997.050 721.050 ;
        RECT 1015.950 720.600 1018.050 721.050 ;
        RECT 994.950 719.400 1018.050 720.600 ;
        RECT 994.950 718.950 997.050 719.400 ;
        RECT 1015.950 718.950 1018.050 719.400 ;
        RECT 1021.950 720.600 1024.050 721.050 ;
        RECT 1042.950 720.600 1045.050 721.050 ;
        RECT 1021.950 719.400 1045.050 720.600 ;
        RECT 1021.950 718.950 1024.050 719.400 ;
        RECT 1042.950 718.950 1045.050 719.400 ;
        RECT 70.950 717.600 73.050 718.050 ;
        RECT 94.950 717.600 97.050 718.050 ;
        RECT 172.950 717.600 175.050 718.050 ;
        RECT 70.950 716.400 175.050 717.600 ;
        RECT 70.950 715.950 73.050 716.400 ;
        RECT 94.950 715.950 97.050 716.400 ;
        RECT 172.950 715.950 175.050 716.400 ;
        RECT 301.950 717.600 304.050 718.050 ;
        RECT 355.950 717.600 358.050 718.050 ;
        RECT 301.950 716.400 358.050 717.600 ;
        RECT 301.950 715.950 304.050 716.400 ;
        RECT 355.950 715.950 358.050 716.400 ;
        RECT 463.950 717.600 466.050 718.050 ;
        RECT 478.950 717.600 481.050 718.050 ;
        RECT 463.950 716.400 481.050 717.600 ;
        RECT 463.950 715.950 466.050 716.400 ;
        RECT 478.950 715.950 481.050 716.400 ;
        RECT 496.950 717.600 499.050 718.050 ;
        RECT 505.950 717.600 508.050 718.050 ;
        RECT 550.950 717.600 553.050 718.050 ;
        RECT 496.950 716.400 553.050 717.600 ;
        RECT 496.950 715.950 499.050 716.400 ;
        RECT 505.950 715.950 508.050 716.400 ;
        RECT 550.950 715.950 553.050 716.400 ;
        RECT 643.950 717.600 646.050 718.050 ;
        RECT 655.950 717.600 658.050 718.050 ;
        RECT 643.950 716.400 658.050 717.600 ;
        RECT 643.950 715.950 646.050 716.400 ;
        RECT 655.950 715.950 658.050 716.400 ;
        RECT 661.950 717.600 664.050 718.050 ;
        RECT 676.950 717.600 679.050 718.050 ;
        RECT 661.950 716.400 679.050 717.600 ;
        RECT 661.950 715.950 664.050 716.400 ;
        RECT 676.950 715.950 679.050 716.400 ;
        RECT 694.950 717.600 697.050 718.050 ;
        RECT 781.950 717.600 784.050 718.050 ;
        RECT 694.950 716.400 784.050 717.600 ;
        RECT 694.950 715.950 697.050 716.400 ;
        RECT 781.950 715.950 784.050 716.400 ;
        RECT 802.950 717.600 805.050 717.900 ;
        RECT 877.950 717.600 880.050 717.900 ;
        RECT 916.950 717.600 919.050 718.050 ;
        RECT 802.950 716.400 816.600 717.600 ;
        RECT 802.950 715.800 805.050 716.400 ;
        RECT 10.950 714.600 13.050 715.050 ;
        RECT 88.950 714.600 91.050 715.050 ;
        RECT 10.950 713.400 91.050 714.600 ;
        RECT 10.950 712.950 13.050 713.400 ;
        RECT 88.950 712.950 91.050 713.400 ;
        RECT 136.950 714.600 139.050 715.050 ;
        RECT 145.950 714.600 148.050 715.050 ;
        RECT 136.950 713.400 148.050 714.600 ;
        RECT 136.950 712.950 139.050 713.400 ;
        RECT 145.950 712.950 148.050 713.400 ;
        RECT 247.950 714.600 250.050 715.050 ;
        RECT 373.950 714.600 376.050 715.050 ;
        RECT 421.950 714.600 424.050 715.050 ;
        RECT 247.950 713.400 424.050 714.600 ;
        RECT 247.950 712.950 250.050 713.400 ;
        RECT 373.950 712.950 376.050 713.400 ;
        RECT 421.950 712.950 424.050 713.400 ;
        RECT 604.950 714.600 607.050 715.050 ;
        RECT 631.950 714.600 634.050 715.050 ;
        RECT 739.950 714.600 742.050 715.050 ;
        RECT 604.950 713.400 742.050 714.600 ;
        RECT 604.950 712.950 607.050 713.400 ;
        RECT 631.950 712.950 634.050 713.400 ;
        RECT 739.950 712.950 742.050 713.400 ;
        RECT 745.950 714.600 748.050 715.050 ;
        RECT 784.950 714.600 787.050 715.050 ;
        RECT 811.950 714.600 814.050 715.050 ;
        RECT 745.950 713.400 814.050 714.600 ;
        RECT 815.400 714.600 816.600 716.400 ;
        RECT 877.950 716.400 919.050 717.600 ;
        RECT 877.950 715.800 880.050 716.400 ;
        RECT 916.950 715.950 919.050 716.400 ;
        RECT 874.950 714.600 877.050 715.050 ;
        RECT 815.400 713.400 877.050 714.600 ;
        RECT 745.950 712.950 748.050 713.400 ;
        RECT 784.950 712.950 787.050 713.400 ;
        RECT 811.950 712.950 814.050 713.400 ;
        RECT 874.950 712.950 877.050 713.400 ;
        RECT 880.950 714.600 883.050 715.050 ;
        RECT 910.950 714.600 913.050 715.050 ;
        RECT 880.950 713.400 913.050 714.600 ;
        RECT 880.950 712.950 883.050 713.400 ;
        RECT 910.950 712.950 913.050 713.400 ;
        RECT 919.950 714.600 922.050 715.050 ;
        RECT 931.950 714.600 934.050 715.050 ;
        RECT 919.950 713.400 934.050 714.600 ;
        RECT 919.950 712.950 922.050 713.400 ;
        RECT 931.950 712.950 934.050 713.400 ;
        RECT 337.950 711.600 340.050 712.050 ;
        RECT 388.950 711.600 391.050 712.050 ;
        RECT 337.950 710.400 391.050 711.600 ;
        RECT 337.950 709.950 340.050 710.400 ;
        RECT 388.950 709.950 391.050 710.400 ;
        RECT 400.950 711.600 403.050 712.050 ;
        RECT 433.950 711.600 436.050 712.050 ;
        RECT 490.950 711.600 493.050 712.050 ;
        RECT 400.950 710.400 493.050 711.600 ;
        RECT 400.950 709.950 403.050 710.400 ;
        RECT 433.950 709.950 436.050 710.400 ;
        RECT 490.950 709.950 493.050 710.400 ;
        RECT 502.950 711.600 505.050 712.050 ;
        RECT 526.950 711.600 529.050 712.050 ;
        RECT 559.950 711.600 562.050 712.050 ;
        RECT 613.950 711.600 616.050 712.050 ;
        RECT 502.950 710.400 558.600 711.600 ;
        RECT 502.950 709.950 505.050 710.400 ;
        RECT 526.950 709.950 529.050 710.400 ;
        RECT 103.950 708.600 106.050 709.050 ;
        RECT 160.950 708.600 163.050 709.050 ;
        RECT 226.950 708.600 229.050 709.050 ;
        RECT 103.950 707.400 229.050 708.600 ;
        RECT 103.950 706.950 106.050 707.400 ;
        RECT 160.950 706.950 163.050 707.400 ;
        RECT 226.950 706.950 229.050 707.400 ;
        RECT 418.950 708.600 421.050 709.050 ;
        RECT 454.950 708.600 457.050 709.050 ;
        RECT 418.950 707.400 457.050 708.600 ;
        RECT 557.400 708.600 558.600 710.400 ;
        RECT 559.950 710.400 616.050 711.600 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 613.950 709.950 616.050 710.400 ;
        RECT 622.950 711.600 625.050 712.050 ;
        RECT 679.950 711.600 682.050 712.050 ;
        RECT 622.950 710.400 682.050 711.600 ;
        RECT 622.950 709.950 625.050 710.400 ;
        RECT 679.950 709.950 682.050 710.400 ;
        RECT 697.950 711.600 700.050 712.050 ;
        RECT 727.950 711.600 730.050 712.050 ;
        RECT 697.950 710.400 730.050 711.600 ;
        RECT 697.950 709.950 700.050 710.400 ;
        RECT 727.950 709.950 730.050 710.400 ;
        RECT 736.950 711.600 739.050 712.050 ;
        RECT 769.950 711.600 772.050 712.050 ;
        RECT 736.950 710.400 772.050 711.600 ;
        RECT 736.950 709.950 739.050 710.400 ;
        RECT 769.950 709.950 772.050 710.400 ;
        RECT 775.950 711.600 778.050 712.050 ;
        RECT 781.950 711.600 784.050 712.050 ;
        RECT 775.950 710.400 784.050 711.600 ;
        RECT 775.950 709.950 778.050 710.400 ;
        RECT 781.950 709.950 784.050 710.400 ;
        RECT 790.950 711.600 793.050 712.050 ;
        RECT 802.950 711.600 805.050 712.050 ;
        RECT 790.950 710.400 805.050 711.600 ;
        RECT 790.950 709.950 793.050 710.400 ;
        RECT 802.950 709.950 805.050 710.400 ;
        RECT 865.950 711.600 868.050 712.050 ;
        RECT 907.950 711.600 910.050 712.050 ;
        RECT 865.950 710.400 910.050 711.600 ;
        RECT 865.950 709.950 868.050 710.400 ;
        RECT 907.950 709.950 910.050 710.400 ;
        RECT 583.800 708.600 585.900 709.050 ;
        RECT 557.400 707.400 585.900 708.600 ;
        RECT 418.950 706.950 421.050 707.400 ;
        RECT 454.950 706.950 457.050 707.400 ;
        RECT 583.800 706.950 585.900 707.400 ;
        RECT 586.950 708.600 589.050 709.050 ;
        RECT 652.950 708.600 655.050 709.050 ;
        RECT 586.950 707.400 655.050 708.600 ;
        RECT 586.950 706.950 589.050 707.400 ;
        RECT 652.950 706.950 655.050 707.400 ;
        RECT 670.950 708.600 673.050 709.050 ;
        RECT 718.950 708.600 721.050 709.050 ;
        RECT 670.950 707.400 721.050 708.600 ;
        RECT 670.950 706.950 673.050 707.400 ;
        RECT 718.950 706.950 721.050 707.400 ;
        RECT 739.950 708.600 742.050 709.050 ;
        RECT 826.950 708.600 829.050 709.050 ;
        RECT 739.950 707.400 829.050 708.600 ;
        RECT 739.950 706.950 742.050 707.400 ;
        RECT 826.950 706.950 829.050 707.400 ;
        RECT 847.950 708.600 850.050 709.050 ;
        RECT 907.950 708.600 910.050 708.900 ;
        RECT 847.950 707.400 910.050 708.600 ;
        RECT 847.950 706.950 850.050 707.400 ;
        RECT 907.950 706.800 910.050 707.400 ;
        RECT 934.950 708.600 937.050 709.050 ;
        RECT 961.950 708.600 964.050 709.050 ;
        RECT 976.950 708.600 979.050 709.050 ;
        RECT 934.950 707.400 979.050 708.600 ;
        RECT 934.950 706.950 937.050 707.400 ;
        RECT 961.950 706.950 964.050 707.400 ;
        RECT 976.950 706.950 979.050 707.400 ;
        RECT 166.950 705.600 169.050 706.050 ;
        RECT 211.950 705.600 214.050 706.050 ;
        RECT 166.950 704.400 214.050 705.600 ;
        RECT 166.950 703.950 169.050 704.400 ;
        RECT 211.950 703.950 214.050 704.400 ;
        RECT 349.950 705.600 352.050 706.050 ;
        RECT 367.950 705.600 370.050 706.050 ;
        RECT 391.950 705.600 394.050 706.050 ;
        RECT 517.950 705.600 520.050 706.050 ;
        RECT 349.950 704.400 520.050 705.600 ;
        RECT 349.950 703.950 352.050 704.400 ;
        RECT 367.950 703.950 370.050 704.400 ;
        RECT 391.950 703.950 394.050 704.400 ;
        RECT 517.950 703.950 520.050 704.400 ;
        RECT 532.950 705.600 535.050 706.050 ;
        RECT 547.950 705.600 550.050 706.050 ;
        RECT 655.950 705.600 658.050 705.900 ;
        RECT 664.950 705.600 667.050 706.050 ;
        RECT 799.950 705.600 802.050 706.050 ;
        RECT 532.950 704.400 667.050 705.600 ;
        RECT 532.950 703.950 535.050 704.400 ;
        RECT 547.950 703.950 550.050 704.400 ;
        RECT 655.950 703.800 658.050 704.400 ;
        RECT 664.950 703.950 667.050 704.400 ;
        RECT 770.400 704.400 802.050 705.600 ;
        RECT 4.950 702.600 7.050 703.050 ;
        RECT 28.950 702.600 31.050 703.050 ;
        RECT 46.950 702.600 49.050 703.050 ;
        RECT 4.950 701.400 49.050 702.600 ;
        RECT 4.950 700.950 7.050 701.400 ;
        RECT 28.950 700.950 31.050 701.400 ;
        RECT 46.950 700.950 49.050 701.400 ;
        RECT 415.950 702.600 418.050 703.050 ;
        RECT 448.950 702.600 451.050 703.050 ;
        RECT 415.950 701.400 451.050 702.600 ;
        RECT 415.950 700.950 418.050 701.400 ;
        RECT 448.950 700.950 451.050 701.400 ;
        RECT 457.950 702.600 460.050 703.050 ;
        RECT 511.950 702.600 514.050 703.050 ;
        RECT 457.950 701.400 514.050 702.600 ;
        RECT 457.950 700.950 460.050 701.400 ;
        RECT 511.950 700.950 514.050 701.400 ;
        RECT 550.950 702.600 553.050 703.050 ;
        RECT 607.950 702.600 610.050 703.050 ;
        RECT 660.000 702.600 664.050 703.050 ;
        RECT 550.950 701.400 654.600 702.600 ;
        RECT 550.950 700.950 553.050 701.400 ;
        RECT 607.950 700.950 610.050 701.400 ;
        RECT 307.950 699.600 310.050 700.050 ;
        RECT 316.950 699.600 319.050 700.050 ;
        RECT 325.950 699.600 328.050 700.050 ;
        RECT 484.950 699.600 487.050 700.050 ;
        RECT 307.950 698.400 487.050 699.600 ;
        RECT 307.950 697.950 310.050 698.400 ;
        RECT 316.950 697.950 319.050 698.400 ;
        RECT 325.950 697.950 328.050 698.400 ;
        RECT 484.950 697.950 487.050 698.400 ;
        RECT 586.950 699.600 589.050 700.050 ;
        RECT 649.950 699.600 652.050 700.050 ;
        RECT 586.950 698.400 652.050 699.600 ;
        RECT 653.400 699.600 654.600 701.400 ;
        RECT 659.400 700.950 664.050 702.600 ;
        RECT 667.950 702.600 670.050 703.050 ;
        RECT 736.950 702.600 739.050 703.050 ;
        RECT 667.950 701.400 739.050 702.600 ;
        RECT 667.950 700.950 670.050 701.400 ;
        RECT 736.950 700.950 739.050 701.400 ;
        RECT 742.950 702.600 745.050 703.050 ;
        RECT 770.400 702.600 771.600 704.400 ;
        RECT 799.950 703.950 802.050 704.400 ;
        RECT 844.950 705.600 847.050 706.050 ;
        RECT 910.950 705.600 913.050 706.050 ;
        RECT 844.950 704.400 913.050 705.600 ;
        RECT 844.950 703.950 847.050 704.400 ;
        RECT 910.950 703.950 913.050 704.400 ;
        RECT 916.950 705.600 919.050 706.050 ;
        RECT 949.950 705.600 952.050 706.050 ;
        RECT 916.950 704.400 952.050 705.600 ;
        RECT 916.950 703.950 919.050 704.400 ;
        RECT 949.950 703.950 952.050 704.400 ;
        RECT 742.950 701.400 771.600 702.600 ;
        RECT 793.950 702.600 796.050 703.050 ;
        RECT 814.950 702.600 817.050 703.050 ;
        RECT 793.950 701.400 817.050 702.600 ;
        RECT 742.950 700.950 745.050 701.400 ;
        RECT 793.950 700.950 796.050 701.400 ;
        RECT 814.950 700.950 817.050 701.400 ;
        RECT 847.950 702.600 850.050 703.050 ;
        RECT 901.950 702.600 904.050 703.050 ;
        RECT 847.950 701.400 904.050 702.600 ;
        RECT 847.950 700.950 850.050 701.400 ;
        RECT 901.950 700.950 904.050 701.400 ;
        RECT 907.950 702.600 910.050 703.050 ;
        RECT 955.950 702.600 958.050 703.050 ;
        RECT 907.950 701.400 958.050 702.600 ;
        RECT 907.950 700.950 910.050 701.400 ;
        RECT 955.950 700.950 958.050 701.400 ;
        RECT 659.400 699.600 660.600 700.950 ;
        RECT 653.400 698.400 660.600 699.600 ;
        RECT 661.950 699.600 664.050 699.900 ;
        RECT 760.950 699.600 763.050 700.050 ;
        RECT 661.950 698.400 763.050 699.600 ;
        RECT 586.950 697.950 589.050 698.400 ;
        RECT 649.950 697.950 652.050 698.400 ;
        RECT 661.950 697.800 664.050 698.400 ;
        RECT 760.950 697.950 763.050 698.400 ;
        RECT 769.950 699.600 772.050 700.050 ;
        RECT 787.950 699.600 790.050 700.050 ;
        RECT 769.950 698.400 790.050 699.600 ;
        RECT 769.950 697.950 772.050 698.400 ;
        RECT 787.950 697.950 790.050 698.400 ;
        RECT 805.950 699.600 808.050 700.050 ;
        RECT 877.950 699.600 880.050 700.050 ;
        RECT 805.950 698.400 880.050 699.600 ;
        RECT 805.950 697.950 808.050 698.400 ;
        RECT 877.950 697.950 880.050 698.400 ;
        RECT 895.950 699.600 898.050 700.050 ;
        RECT 934.950 699.600 937.050 700.050 ;
        RECT 895.950 698.400 937.050 699.600 ;
        RECT 895.950 697.950 898.050 698.400 ;
        RECT 934.950 697.950 937.050 698.400 ;
        RECT 424.950 696.600 427.050 697.050 ;
        RECT 505.950 696.600 508.050 697.050 ;
        RECT 424.950 695.400 508.050 696.600 ;
        RECT 424.950 694.950 427.050 695.400 ;
        RECT 505.950 694.950 508.050 695.400 ;
        RECT 541.950 696.600 544.050 697.050 ;
        RECT 580.950 696.600 583.050 697.050 ;
        RECT 541.950 695.400 583.050 696.600 ;
        RECT 541.950 694.950 544.050 695.400 ;
        RECT 580.950 694.950 583.050 695.400 ;
        RECT 637.950 696.600 640.050 697.050 ;
        RECT 676.950 696.600 679.050 697.050 ;
        RECT 637.950 695.400 679.050 696.600 ;
        RECT 637.950 694.950 640.050 695.400 ;
        RECT 676.950 694.950 679.050 695.400 ;
        RECT 757.950 696.600 760.050 697.050 ;
        RECT 781.950 696.600 784.050 697.050 ;
        RECT 757.950 695.400 784.050 696.600 ;
        RECT 757.950 694.950 760.050 695.400 ;
        RECT 781.950 694.950 784.050 695.400 ;
        RECT 805.950 696.600 808.050 696.900 ;
        RECT 814.950 696.600 817.050 697.050 ;
        RECT 805.950 695.400 817.050 696.600 ;
        RECT 805.950 694.800 808.050 695.400 ;
        RECT 814.950 694.950 817.050 695.400 ;
        RECT 823.950 696.600 826.050 697.050 ;
        RECT 847.950 696.600 850.050 697.050 ;
        RECT 823.950 695.400 850.050 696.600 ;
        RECT 823.950 694.950 826.050 695.400 ;
        RECT 847.950 694.950 850.050 695.400 ;
        RECT 856.950 696.600 859.050 697.050 ;
        RECT 871.950 696.600 874.050 697.050 ;
        RECT 856.950 695.400 874.050 696.600 ;
        RECT 856.950 694.950 859.050 695.400 ;
        RECT 871.950 694.950 874.050 695.400 ;
        RECT 883.950 696.600 886.050 697.050 ;
        RECT 946.950 696.600 949.050 697.050 ;
        RECT 883.950 695.400 949.050 696.600 ;
        RECT 883.950 694.950 886.050 695.400 ;
        RECT 946.950 694.950 949.050 695.400 ;
        RECT 964.950 696.600 967.050 697.050 ;
        RECT 1024.950 696.600 1027.050 697.050 ;
        RECT 964.950 695.400 1027.050 696.600 ;
        RECT 964.950 694.950 967.050 695.400 ;
        RECT 1024.950 694.950 1027.050 695.400 ;
        RECT 322.950 693.600 325.050 694.050 ;
        RECT 346.950 693.600 349.050 694.050 ;
        RECT 322.950 692.400 349.050 693.600 ;
        RECT 322.950 691.950 325.050 692.400 ;
        RECT 346.950 691.950 349.050 692.400 ;
        RECT 376.950 693.600 379.050 694.050 ;
        RECT 412.950 693.600 415.050 694.050 ;
        RECT 376.950 692.400 415.050 693.600 ;
        RECT 376.950 691.950 379.050 692.400 ;
        RECT 412.950 691.950 415.050 692.400 ;
        RECT 427.950 693.600 430.050 694.050 ;
        RECT 502.950 693.600 505.050 694.050 ;
        RECT 427.950 692.400 505.050 693.600 ;
        RECT 427.950 691.950 430.050 692.400 ;
        RECT 502.950 691.950 505.050 692.400 ;
        RECT 526.950 693.600 529.050 694.050 ;
        RECT 568.950 693.600 571.050 694.050 ;
        RECT 526.950 692.400 571.050 693.600 ;
        RECT 526.950 691.950 529.050 692.400 ;
        RECT 568.950 691.950 571.050 692.400 ;
        RECT 619.950 693.600 622.050 694.050 ;
        RECT 688.950 693.600 691.050 694.050 ;
        RECT 619.950 692.400 691.050 693.600 ;
        RECT 619.950 691.950 622.050 692.400 ;
        RECT 688.950 691.950 691.050 692.400 ;
        RECT 715.950 693.600 718.050 694.050 ;
        RECT 730.950 693.600 733.050 694.050 ;
        RECT 820.950 693.600 823.050 694.050 ;
        RECT 715.950 692.400 733.050 693.600 ;
        RECT 715.950 691.950 718.050 692.400 ;
        RECT 730.950 691.950 733.050 692.400 ;
        RECT 734.400 692.400 823.050 693.600 ;
        RECT 34.950 687.600 37.050 691.050 ;
        RECT 49.950 690.600 52.050 691.050 ;
        RECT 73.950 690.600 76.050 691.050 ;
        RECT 136.950 690.600 139.050 691.050 ;
        RECT 49.950 689.400 60.600 690.600 ;
        RECT 49.950 688.950 52.050 689.400 ;
        RECT 34.950 687.000 57.600 687.600 ;
        RECT 35.400 686.400 57.600 687.000 ;
        RECT 52.950 681.600 55.050 685.050 ;
        RECT 32.400 681.000 55.050 681.600 ;
        RECT 32.400 680.400 54.600 681.000 ;
        RECT 32.400 678.900 33.600 680.400 ;
        RECT 22.950 678.450 25.050 678.900 ;
        RECT 31.950 678.450 34.050 678.900 ;
        RECT 22.950 677.250 34.050 678.450 ;
        RECT 22.950 676.800 25.050 677.250 ;
        RECT 31.950 676.800 34.050 677.250 ;
        RECT 34.950 675.600 37.050 676.050 ;
        RECT 56.400 675.600 57.600 686.400 ;
        RECT 59.400 684.600 60.600 689.400 ;
        RECT 73.950 689.400 139.050 690.600 ;
        RECT 73.950 688.950 76.050 689.400 ;
        RECT 136.950 688.950 139.050 689.400 ;
        RECT 178.950 690.600 181.050 691.050 ;
        RECT 193.950 690.600 196.050 691.050 ;
        RECT 178.950 689.400 196.050 690.600 ;
        RECT 178.950 688.950 181.050 689.400 ;
        RECT 193.950 688.950 196.050 689.400 ;
        RECT 421.950 690.600 424.050 691.050 ;
        RECT 457.950 690.600 460.050 691.050 ;
        RECT 592.950 690.600 595.050 691.050 ;
        RECT 421.950 689.400 460.050 690.600 ;
        RECT 421.950 688.950 424.050 689.400 ;
        RECT 457.950 688.950 460.050 689.400 ;
        RECT 509.400 689.400 595.050 690.600 ;
        RECT 127.950 687.600 130.050 688.050 ;
        RECT 142.950 687.600 145.050 688.050 ;
        RECT 127.950 686.400 145.050 687.600 ;
        RECT 127.950 685.950 130.050 686.400 ;
        RECT 142.950 685.950 145.050 686.400 ;
        RECT 163.950 687.600 166.050 688.050 ;
        RECT 187.950 687.600 190.050 688.050 ;
        RECT 163.950 686.400 190.050 687.600 ;
        RECT 163.950 685.950 166.050 686.400 ;
        RECT 187.950 685.950 190.050 686.400 ;
        RECT 340.950 687.600 343.050 688.050 ;
        RECT 352.950 687.600 355.050 688.050 ;
        RECT 340.950 686.400 355.050 687.600 ;
        RECT 340.950 685.950 343.050 686.400 ;
        RECT 352.950 685.950 355.050 686.400 ;
        RECT 397.950 687.600 400.050 688.050 ;
        RECT 403.950 687.600 406.050 688.050 ;
        RECT 427.950 687.600 430.050 688.050 ;
        RECT 432.000 687.600 436.050 688.050 ;
        RECT 397.950 686.400 430.050 687.600 ;
        RECT 397.950 685.950 400.050 686.400 ;
        RECT 403.950 685.950 406.050 686.400 ;
        RECT 427.950 685.950 430.050 686.400 ;
        RECT 431.400 685.950 436.050 687.600 ;
        RECT 502.950 687.600 505.050 688.050 ;
        RECT 509.400 687.600 510.600 689.400 ;
        RECT 592.950 688.950 595.050 689.400 ;
        RECT 598.950 690.600 601.050 691.050 ;
        RECT 631.950 690.600 634.050 691.050 ;
        RECT 643.950 690.600 646.050 691.050 ;
        RECT 598.950 689.400 646.050 690.600 ;
        RECT 598.950 688.950 601.050 689.400 ;
        RECT 631.950 688.950 634.050 689.400 ;
        RECT 643.950 688.950 646.050 689.400 ;
        RECT 664.950 690.600 667.050 691.050 ;
        RECT 694.950 690.600 697.050 691.050 ;
        RECT 664.950 689.400 697.050 690.600 ;
        RECT 664.950 688.950 667.050 689.400 ;
        RECT 694.950 688.950 697.050 689.400 ;
        RECT 703.950 690.600 706.050 691.050 ;
        RECT 734.400 690.600 735.600 692.400 ;
        RECT 820.950 691.950 823.050 692.400 ;
        RECT 838.950 693.600 841.050 694.050 ;
        RECT 838.950 692.400 951.600 693.600 ;
        RECT 838.950 691.950 841.050 692.400 ;
        RECT 950.400 691.050 951.600 692.400 ;
        RECT 703.950 689.400 735.600 690.600 ;
        RECT 745.950 690.600 748.050 691.050 ;
        RECT 802.950 690.600 805.050 691.050 ;
        RECT 745.950 689.400 805.050 690.600 ;
        RECT 703.950 688.950 706.050 689.400 ;
        RECT 745.950 688.950 748.050 689.400 ;
        RECT 802.950 688.950 805.050 689.400 ;
        RECT 826.950 690.600 829.050 691.050 ;
        RECT 907.800 690.600 909.900 691.050 ;
        RECT 826.950 689.400 909.900 690.600 ;
        RECT 826.950 688.950 829.050 689.400 ;
        RECT 907.800 688.950 909.900 689.400 ;
        RECT 910.950 690.600 913.050 691.050 ;
        RECT 925.950 690.600 928.050 691.050 ;
        RECT 910.950 689.400 928.050 690.600 ;
        RECT 950.400 689.400 955.050 691.050 ;
        RECT 910.950 688.950 913.050 689.400 ;
        RECT 925.950 688.950 928.050 689.400 ;
        RECT 951.000 688.950 955.050 689.400 ;
        RECT 988.950 690.600 991.050 691.050 ;
        RECT 1000.950 690.600 1003.050 691.050 ;
        RECT 988.950 689.400 1003.050 690.600 ;
        RECT 988.950 688.950 991.050 689.400 ;
        RECT 1000.950 688.950 1003.050 689.400 ;
        RECT 502.950 686.400 510.600 687.600 ;
        RECT 511.950 687.600 514.050 688.050 ;
        RECT 532.950 687.600 535.050 688.050 ;
        RECT 511.950 686.400 535.050 687.600 ;
        RECT 502.950 685.950 505.050 686.400 ;
        RECT 511.950 685.950 514.050 686.400 ;
        RECT 532.950 685.950 535.050 686.400 ;
        RECT 553.950 687.600 556.050 688.050 ;
        RECT 580.950 687.600 583.050 688.050 ;
        RECT 553.950 686.400 583.050 687.600 ;
        RECT 553.950 685.950 556.050 686.400 ;
        RECT 580.950 685.950 583.050 686.400 ;
        RECT 613.950 687.600 616.050 688.050 ;
        RECT 625.950 687.600 628.050 688.050 ;
        RECT 613.950 686.400 628.050 687.600 ;
        RECT 613.950 685.950 616.050 686.400 ;
        RECT 625.950 685.950 628.050 686.400 ;
        RECT 658.950 687.600 661.050 688.050 ;
        RECT 667.950 687.600 670.050 688.050 ;
        RECT 697.950 687.600 700.050 688.050 ;
        RECT 658.950 686.400 700.050 687.600 ;
        RECT 658.950 685.950 661.050 686.400 ;
        RECT 667.950 685.950 670.050 686.400 ;
        RECT 697.950 685.950 700.050 686.400 ;
        RECT 739.950 687.600 742.050 688.050 ;
        RECT 784.950 687.600 787.050 688.050 ;
        RECT 799.950 687.600 802.050 688.050 ;
        RECT 739.950 686.400 787.050 687.600 ;
        RECT 739.950 685.950 742.050 686.400 ;
        RECT 784.950 685.950 787.050 686.400 ;
        RECT 788.400 686.400 802.050 687.600 ;
        RECT 112.950 684.600 115.050 685.200 ;
        RECT 59.400 683.400 115.050 684.600 ;
        RECT 112.950 683.100 115.050 683.400 ;
        RECT 151.950 684.750 154.050 685.200 ;
        RECT 160.950 684.750 163.050 685.200 ;
        RECT 151.950 683.550 163.050 684.750 ;
        RECT 151.950 683.100 154.050 683.550 ;
        RECT 160.950 683.100 163.050 683.550 ;
        RECT 220.950 684.600 223.050 685.050 ;
        RECT 232.950 684.600 235.050 685.200 ;
        RECT 220.950 683.400 235.050 684.600 ;
        RECT 220.950 682.950 223.050 683.400 ;
        RECT 232.950 683.100 235.050 683.400 ;
        RECT 268.950 684.750 271.050 685.200 ;
        RECT 274.950 684.750 277.050 685.200 ;
        RECT 268.950 683.550 277.050 684.750 ;
        RECT 268.950 683.100 271.050 683.550 ;
        RECT 274.950 683.100 277.050 683.550 ;
        RECT 289.950 684.600 292.050 685.200 ;
        RECT 313.950 684.600 316.050 685.200 ;
        RECT 322.950 684.600 325.050 685.050 ;
        RECT 289.950 683.400 325.050 684.600 ;
        RECT 289.950 683.100 292.050 683.400 ;
        RECT 313.950 683.100 316.050 683.400 ;
        RECT 322.950 682.950 325.050 683.400 ;
        RECT 328.950 684.600 331.050 685.050 ;
        RECT 337.950 684.600 340.050 685.200 ;
        RECT 328.950 683.400 340.050 684.600 ;
        RECT 328.950 682.950 331.050 683.400 ;
        RECT 337.950 683.100 340.050 683.400 ;
        RECT 355.950 684.600 358.050 685.050 ;
        RECT 367.950 684.600 370.050 685.200 ;
        RECT 355.950 683.400 370.050 684.600 ;
        RECT 355.950 682.950 358.050 683.400 ;
        RECT 367.950 683.100 370.050 683.400 ;
        RECT 400.950 682.950 403.050 685.050 ;
        RECT 431.400 684.600 432.600 685.950 ;
        RECT 788.400 685.200 789.600 686.400 ;
        RECT 799.950 685.950 802.050 686.400 ;
        RECT 844.950 687.600 847.050 688.050 ;
        RECT 868.950 687.600 871.050 688.050 ;
        RECT 880.950 687.600 883.050 688.050 ;
        RECT 844.950 686.400 867.600 687.600 ;
        RECT 844.950 685.950 847.050 686.400 ;
        RECT 428.400 683.400 432.600 684.600 ;
        RECT 433.950 684.600 436.050 684.900 ;
        RECT 445.950 684.600 448.050 685.200 ;
        RECT 466.950 684.600 469.050 685.200 ;
        RECT 433.950 683.400 469.050 684.600 ;
        RECT 79.950 678.600 82.050 679.050 ;
        RECT 91.950 678.600 94.050 679.050 ;
        RECT 79.950 677.400 94.050 678.600 ;
        RECT 79.950 676.950 82.050 677.400 ;
        RECT 91.950 676.950 94.050 677.400 ;
        RECT 97.950 678.450 100.050 678.900 ;
        RECT 109.950 678.450 112.050 678.900 ;
        RECT 97.950 677.250 112.050 678.450 ;
        RECT 97.950 676.800 100.050 677.250 ;
        RECT 109.950 676.800 112.050 677.250 ;
        RECT 115.950 678.450 118.050 678.900 ;
        RECT 127.950 678.450 130.050 678.900 ;
        RECT 115.950 677.250 130.050 678.450 ;
        RECT 115.950 676.800 118.050 677.250 ;
        RECT 127.950 676.800 130.050 677.250 ;
        RECT 139.950 678.600 142.050 678.900 ;
        RECT 154.950 678.600 157.050 679.050 ;
        RECT 139.950 677.400 157.050 678.600 ;
        RECT 139.950 676.800 142.050 677.400 ;
        RECT 154.950 676.950 157.050 677.400 ;
        RECT 163.950 678.600 166.050 678.900 ;
        RECT 175.950 678.600 178.050 679.050 ;
        RECT 163.950 677.400 178.050 678.600 ;
        RECT 163.950 676.800 166.050 677.400 ;
        RECT 175.950 676.950 178.050 677.400 ;
        RECT 181.950 678.600 184.050 679.050 ;
        RECT 196.950 678.600 199.050 679.050 ;
        RECT 181.950 677.400 199.050 678.600 ;
        RECT 181.950 676.950 184.050 677.400 ;
        RECT 196.950 676.950 199.050 677.400 ;
        RECT 253.950 678.450 256.050 678.900 ;
        RECT 271.800 678.450 273.900 678.900 ;
        RECT 253.950 677.250 273.900 678.450 ;
        RECT 253.950 676.800 256.050 677.250 ;
        RECT 271.800 676.800 273.900 677.250 ;
        RECT 274.950 678.450 277.050 678.900 ;
        RECT 286.950 678.450 289.050 678.900 ;
        RECT 274.950 677.250 289.050 678.450 ;
        RECT 274.950 676.800 277.050 677.250 ;
        RECT 286.950 676.800 289.050 677.250 ;
        RECT 316.950 678.600 319.050 678.900 ;
        RECT 334.950 678.600 337.050 678.900 ;
        RECT 316.950 678.450 337.050 678.600 ;
        RECT 340.950 678.450 343.050 678.900 ;
        RECT 316.950 677.400 343.050 678.450 ;
        RECT 316.950 676.800 319.050 677.400 ;
        RECT 334.950 677.250 343.050 677.400 ;
        RECT 334.950 676.800 337.050 677.250 ;
        RECT 340.950 676.800 343.050 677.250 ;
        RECT 349.950 678.450 352.050 678.900 ;
        RECT 364.950 678.450 367.050 678.900 ;
        RECT 349.950 677.250 367.050 678.450 ;
        RECT 349.950 676.800 352.050 677.250 ;
        RECT 364.950 676.800 367.050 677.250 ;
        RECT 370.950 678.600 373.050 678.900 ;
        RECT 382.950 678.600 385.050 678.900 ;
        RECT 370.950 678.450 385.050 678.600 ;
        RECT 388.950 678.450 391.050 678.900 ;
        RECT 370.950 677.400 391.050 678.450 ;
        RECT 401.400 678.600 402.600 682.950 ;
        RECT 418.950 678.600 421.050 678.900 ;
        RECT 401.400 677.400 421.050 678.600 ;
        RECT 370.950 676.800 373.050 677.400 ;
        RECT 382.950 677.250 391.050 677.400 ;
        RECT 382.950 676.800 385.050 677.250 ;
        RECT 388.950 676.800 391.050 677.250 ;
        RECT 418.950 676.800 421.050 677.400 ;
        RECT 424.950 678.600 427.050 678.900 ;
        RECT 428.400 678.600 429.600 683.400 ;
        RECT 433.950 682.800 436.050 683.400 ;
        RECT 445.950 683.100 448.050 683.400 ;
        RECT 466.950 683.100 469.050 683.400 ;
        RECT 472.950 684.750 475.050 685.200 ;
        RECT 481.950 684.750 484.050 684.900 ;
        RECT 472.950 684.600 484.050 684.750 ;
        RECT 493.950 684.600 496.050 685.200 ;
        RECT 472.950 683.550 496.050 684.600 ;
        RECT 472.950 683.100 475.050 683.550 ;
        RECT 481.950 683.400 496.050 683.550 ;
        RECT 481.950 682.800 484.050 683.400 ;
        RECT 493.950 683.100 496.050 683.400 ;
        RECT 547.950 684.600 550.050 685.200 ;
        RECT 574.950 684.600 577.050 685.200 ;
        RECT 547.950 683.400 564.600 684.600 ;
        RECT 547.950 683.100 550.050 683.400 ;
        RECT 563.400 681.600 564.600 683.400 ;
        RECT 574.950 683.400 579.600 684.600 ;
        RECT 574.950 683.100 577.050 683.400 ;
        RECT 563.400 680.400 570.600 681.600 ;
        RECT 424.950 677.400 429.600 678.600 ;
        RECT 448.950 678.450 451.050 678.900 ;
        RECT 505.950 678.450 508.050 678.900 ;
        RECT 424.950 676.800 427.050 677.400 ;
        RECT 448.950 677.250 508.050 678.450 ;
        RECT 448.950 676.800 451.050 677.250 ;
        RECT 505.950 676.800 508.050 677.250 ;
        RECT 520.950 678.600 523.050 678.900 ;
        RECT 529.950 678.600 532.050 679.050 ;
        RECT 520.950 677.400 532.050 678.600 ;
        RECT 520.950 676.800 523.050 677.400 ;
        RECT 529.950 676.950 532.050 677.400 ;
        RECT 559.950 678.450 562.050 678.900 ;
        RECT 565.950 678.450 568.050 678.900 ;
        RECT 559.950 677.250 568.050 678.450 ;
        RECT 569.400 678.600 570.600 680.400 ;
        RECT 571.950 678.600 574.050 678.900 ;
        RECT 569.400 677.400 574.050 678.600 ;
        RECT 578.400 678.600 579.600 683.400 ;
        RECT 583.950 681.600 586.050 682.050 ;
        RECT 628.950 681.600 631.050 685.050 ;
        RECT 634.950 684.750 637.050 685.200 ;
        RECT 643.950 684.750 646.050 685.200 ;
        RECT 634.950 683.550 646.050 684.750 ;
        RECT 703.950 684.600 706.050 685.200 ;
        RECT 634.950 683.100 637.050 683.550 ;
        RECT 643.950 683.100 646.050 683.550 ;
        RECT 680.400 683.400 706.050 684.600 ;
        RECT 583.950 681.000 631.050 681.600 ;
        RECT 583.950 680.400 630.600 681.000 ;
        RECT 583.950 679.950 586.050 680.400 ;
        RECT 623.400 678.900 624.600 680.400 ;
        RECT 616.950 678.600 619.050 678.900 ;
        RECT 578.400 677.400 619.050 678.600 ;
        RECT 559.950 676.800 562.050 677.250 ;
        RECT 565.950 676.800 568.050 677.250 ;
        RECT 571.950 676.800 574.050 677.400 ;
        RECT 616.950 676.800 619.050 677.400 ;
        RECT 622.950 676.800 625.050 678.900 ;
        RECT 646.950 678.450 649.050 678.900 ;
        RECT 658.950 678.450 661.050 678.900 ;
        RECT 646.950 677.250 661.050 678.450 ;
        RECT 646.950 676.800 649.050 677.250 ;
        RECT 658.950 676.800 661.050 677.250 ;
        RECT 676.950 678.600 679.050 678.900 ;
        RECT 680.400 678.600 681.600 683.400 ;
        RECT 703.950 683.100 706.050 683.400 ;
        RECT 751.950 684.600 754.050 685.200 ;
        RECT 760.950 684.600 763.050 685.050 ;
        RECT 751.950 683.400 763.050 684.600 ;
        RECT 751.950 683.100 754.050 683.400 ;
        RECT 760.950 682.950 763.050 683.400 ;
        RECT 775.950 684.600 778.050 685.200 ;
        RECT 775.950 683.400 783.600 684.600 ;
        RECT 775.950 683.100 778.050 683.400 ;
        RECT 685.950 681.600 688.050 682.050 ;
        RECT 741.000 681.600 745.050 682.050 ;
        RECT 685.950 680.400 702.600 681.600 ;
        RECT 685.950 679.950 688.050 680.400 ;
        RECT 676.950 677.400 681.600 678.600 ;
        RECT 688.950 678.600 691.050 679.050 ;
        RECT 701.400 678.900 702.600 680.400 ;
        RECT 740.400 679.950 745.050 681.600 ;
        RECT 782.400 681.600 783.600 683.400 ;
        RECT 787.950 683.100 790.050 685.200 ;
        RECT 811.950 682.950 814.050 685.050 ;
        RECT 823.800 682.950 825.900 685.050 ;
        RECT 826.950 684.600 829.050 685.200 ;
        RECT 847.950 684.600 850.050 685.200 ;
        RECT 826.950 683.400 850.050 684.600 ;
        RECT 826.950 683.100 829.050 683.400 ;
        RECT 847.950 683.100 850.050 683.400 ;
        RECT 853.950 684.750 856.050 685.200 ;
        RECT 862.950 684.750 865.050 685.200 ;
        RECT 853.950 683.550 865.050 684.750 ;
        RECT 853.950 683.100 856.050 683.550 ;
        RECT 862.950 683.100 865.050 683.550 ;
        RECT 866.400 684.600 867.600 686.400 ;
        RECT 868.950 686.400 883.050 687.600 ;
        RECT 868.950 685.950 871.050 686.400 ;
        RECT 880.950 685.950 883.050 686.400 ;
        RECT 898.950 684.600 901.050 685.200 ;
        RECT 866.400 683.400 901.050 684.600 ;
        RECT 898.950 683.100 901.050 683.400 ;
        RECT 904.950 683.100 907.050 685.200 ;
        RECT 925.950 684.750 928.050 685.200 ;
        RECT 937.950 684.750 940.050 685.200 ;
        RECT 925.950 683.550 940.050 684.750 ;
        RECT 925.950 683.100 928.050 683.550 ;
        RECT 937.950 683.100 940.050 683.550 ;
        RECT 952.950 684.750 955.050 685.200 ;
        RECT 967.950 684.750 970.050 685.200 ;
        RECT 952.950 683.550 970.050 684.750 ;
        RECT 952.950 683.100 955.050 683.550 ;
        RECT 967.950 683.100 970.050 683.550 ;
        RECT 985.950 684.600 988.050 685.050 ;
        RECT 991.950 684.600 994.050 685.200 ;
        RECT 985.950 683.400 994.050 684.600 ;
        RECT 782.400 680.400 786.600 681.600 ;
        RECT 694.950 678.600 697.050 678.900 ;
        RECT 688.950 677.400 697.050 678.600 ;
        RECT 676.950 676.800 679.050 677.400 ;
        RECT 688.950 676.950 691.050 677.400 ;
        RECT 694.950 676.800 697.050 677.400 ;
        RECT 700.950 678.600 703.050 678.900 ;
        RECT 730.950 678.600 733.050 678.900 ;
        RECT 740.400 678.600 741.600 679.950 ;
        RECT 700.950 677.400 741.600 678.600 ;
        RECT 766.950 678.600 769.050 679.050 ;
        RECT 778.950 678.600 781.050 678.900 ;
        RECT 766.950 677.400 781.050 678.600 ;
        RECT 785.400 678.600 786.600 680.400 ;
        RECT 812.400 679.050 813.600 682.950 ;
        RECT 793.950 678.600 796.050 679.050 ;
        RECT 785.400 677.400 796.050 678.600 ;
        RECT 700.950 676.800 703.050 677.400 ;
        RECT 730.950 676.800 733.050 677.400 ;
        RECT 766.950 676.950 769.050 677.400 ;
        RECT 778.950 676.800 781.050 677.400 ;
        RECT 793.950 676.950 796.050 677.400 ;
        RECT 811.950 676.950 814.050 679.050 ;
        RECT 34.950 674.400 57.600 675.600 ;
        RECT 133.950 675.600 136.050 676.050 ;
        RECT 160.950 675.600 163.050 676.050 ;
        RECT 133.950 674.400 163.050 675.600 ;
        RECT 34.950 673.950 37.050 674.400 ;
        RECT 133.950 673.950 136.050 674.400 ;
        RECT 160.950 673.950 163.050 674.400 ;
        RECT 436.950 675.600 439.050 676.050 ;
        RECT 442.950 675.600 445.050 676.050 ;
        RECT 436.950 674.400 445.050 675.600 ;
        RECT 436.950 673.950 439.050 674.400 ;
        RECT 442.950 673.950 445.050 674.400 ;
        RECT 457.950 675.600 460.050 676.050 ;
        RECT 496.950 675.600 499.050 676.050 ;
        RECT 502.950 675.600 505.050 676.050 ;
        RECT 457.950 674.400 505.050 675.600 ;
        RECT 457.950 673.950 460.050 674.400 ;
        RECT 496.950 673.950 499.050 674.400 ;
        RECT 502.950 673.950 505.050 674.400 ;
        RECT 592.950 675.600 595.050 676.050 ;
        RECT 601.950 675.600 604.050 676.050 ;
        RECT 592.950 674.400 604.050 675.600 ;
        RECT 592.950 673.950 595.050 674.400 ;
        RECT 601.950 673.950 604.050 674.400 ;
        RECT 694.950 675.600 697.050 675.750 ;
        RECT 733.950 675.600 736.050 676.050 ;
        RECT 694.950 674.400 736.050 675.600 ;
        RECT 88.950 672.600 91.050 673.050 ;
        RECT 124.950 672.600 127.050 673.050 ;
        RECT 134.400 672.600 135.600 673.950 ;
        RECT 694.950 673.650 697.050 674.400 ;
        RECT 733.950 673.950 736.050 674.400 ;
        RECT 790.950 675.600 793.050 676.050 ;
        RECT 814.950 675.600 817.050 676.050 ;
        RECT 790.950 674.400 817.050 675.600 ;
        RECT 790.950 673.950 793.050 674.400 ;
        RECT 814.950 673.950 817.050 674.400 ;
        RECT 88.950 671.400 135.600 672.600 ;
        RECT 169.950 672.600 172.050 673.050 ;
        RECT 178.950 672.600 181.050 673.050 ;
        RECT 169.950 671.400 181.050 672.600 ;
        RECT 88.950 670.950 91.050 671.400 ;
        RECT 124.950 670.950 127.050 671.400 ;
        RECT 169.950 670.950 172.050 671.400 ;
        RECT 178.950 670.950 181.050 671.400 ;
        RECT 235.950 672.600 238.050 673.050 ;
        RECT 259.950 672.600 262.050 673.050 ;
        RECT 265.950 672.600 268.050 673.050 ;
        RECT 235.950 671.400 268.050 672.600 ;
        RECT 235.950 670.950 238.050 671.400 ;
        RECT 259.950 670.950 262.050 671.400 ;
        RECT 265.950 670.950 268.050 671.400 ;
        RECT 271.950 672.600 274.050 673.050 ;
        RECT 292.950 672.600 295.050 673.050 ;
        RECT 433.950 672.600 436.050 673.050 ;
        RECT 271.950 671.400 436.050 672.600 ;
        RECT 271.950 670.950 274.050 671.400 ;
        RECT 292.950 670.950 295.050 671.400 ;
        RECT 433.950 670.950 436.050 671.400 ;
        RECT 460.950 672.600 463.050 673.050 ;
        RECT 469.950 672.600 472.050 673.050 ;
        RECT 460.950 671.400 472.050 672.600 ;
        RECT 460.950 670.950 463.050 671.400 ;
        RECT 469.950 670.950 472.050 671.400 ;
        RECT 508.950 672.600 511.050 673.050 ;
        RECT 517.950 672.600 520.050 673.050 ;
        RECT 508.950 671.400 520.050 672.600 ;
        RECT 508.950 670.950 511.050 671.400 ;
        RECT 517.950 670.950 520.050 671.400 ;
        RECT 532.950 672.600 535.050 673.050 ;
        RECT 541.950 672.600 544.050 673.050 ;
        RECT 532.950 671.400 544.050 672.600 ;
        RECT 532.950 670.950 535.050 671.400 ;
        RECT 541.950 670.950 544.050 671.400 ;
        RECT 655.950 672.600 658.050 673.050 ;
        RECT 667.950 672.600 670.050 673.050 ;
        RECT 655.950 671.400 670.050 672.600 ;
        RECT 655.950 670.950 658.050 671.400 ;
        RECT 667.950 670.950 670.050 671.400 ;
        RECT 685.950 672.600 688.050 673.050 ;
        RECT 739.950 672.600 742.050 673.050 ;
        RECT 685.950 671.400 742.050 672.600 ;
        RECT 685.950 670.950 688.050 671.400 ;
        RECT 739.950 670.950 742.050 671.400 ;
        RECT 793.950 672.600 796.050 673.050 ;
        RECT 805.950 672.600 808.050 673.050 ;
        RECT 824.400 672.900 825.600 682.950 ;
        RECT 905.400 681.600 906.600 683.100 ;
        RECT 985.950 682.950 988.050 683.400 ;
        RECT 991.950 683.100 994.050 683.400 ;
        RECT 1009.950 684.600 1012.050 685.050 ;
        RECT 1015.950 684.600 1018.050 685.200 ;
        RECT 1009.950 683.400 1018.050 684.600 ;
        RECT 1009.950 682.950 1012.050 683.400 ;
        RECT 1015.950 683.100 1018.050 683.400 ;
        RECT 1021.950 684.750 1024.050 685.200 ;
        RECT 1039.950 684.750 1042.050 685.200 ;
        RECT 1021.950 683.550 1042.050 684.750 ;
        RECT 1021.950 683.100 1024.050 683.550 ;
        RECT 1039.950 683.100 1042.050 683.550 ;
        RECT 916.950 681.600 919.050 682.050 ;
        RECT 905.400 680.400 919.050 681.600 ;
        RECT 916.950 679.950 919.050 680.400 ;
        RECT 986.400 679.050 987.600 682.950 ;
        RECT 829.950 678.450 832.050 678.900 ;
        RECT 838.950 678.450 841.050 678.900 ;
        RECT 829.950 677.250 841.050 678.450 ;
        RECT 829.950 676.800 832.050 677.250 ;
        RECT 838.950 676.800 841.050 677.250 ;
        RECT 862.950 678.600 865.050 679.050 ;
        RECT 871.950 678.600 874.050 678.900 ;
        RECT 862.950 677.400 874.050 678.600 ;
        RECT 862.950 676.950 865.050 677.400 ;
        RECT 871.950 676.800 874.050 677.400 ;
        RECT 883.950 678.600 886.050 679.050 ;
        RECT 907.950 678.600 910.050 678.900 ;
        RECT 883.950 677.400 910.050 678.600 ;
        RECT 883.950 676.950 886.050 677.400 ;
        RECT 907.950 676.800 910.050 677.400 ;
        RECT 925.950 678.600 928.050 679.050 ;
        RECT 943.950 678.600 946.050 678.900 ;
        RECT 925.950 677.400 946.050 678.600 ;
        RECT 925.950 676.950 928.050 677.400 ;
        RECT 943.950 676.800 946.050 677.400 ;
        RECT 955.950 678.450 958.050 678.900 ;
        RECT 964.950 678.450 967.050 678.900 ;
        RECT 955.950 677.250 967.050 678.450 ;
        RECT 955.950 676.800 958.050 677.250 ;
        RECT 964.950 676.800 967.050 677.250 ;
        RECT 985.950 676.950 988.050 679.050 ;
        RECT 1003.950 678.600 1006.050 679.050 ;
        RECT 1012.950 678.600 1015.050 678.900 ;
        RECT 1003.950 677.400 1015.050 678.600 ;
        RECT 1003.950 676.950 1006.050 677.400 ;
        RECT 1012.950 676.800 1015.050 677.400 ;
        RECT 1016.400 676.050 1017.600 683.100 ;
        RECT 826.950 675.600 829.050 676.050 ;
        RECT 850.950 675.600 853.050 676.050 ;
        RECT 826.950 674.400 853.050 675.600 ;
        RECT 826.950 673.950 829.050 674.400 ;
        RECT 850.950 673.950 853.050 674.400 ;
        RECT 889.950 675.600 892.050 676.050 ;
        RECT 901.800 675.600 903.900 676.050 ;
        RECT 889.950 674.400 903.900 675.600 ;
        RECT 889.950 673.950 892.050 674.400 ;
        RECT 901.800 673.950 903.900 674.400 ;
        RECT 904.950 675.600 907.050 676.050 ;
        RECT 913.950 675.600 916.050 676.050 ;
        RECT 904.950 674.400 916.050 675.600 ;
        RECT 904.950 673.950 907.050 674.400 ;
        RECT 913.950 673.950 916.050 674.400 ;
        RECT 1015.950 673.950 1018.050 676.050 ;
        RECT 793.950 671.400 808.050 672.600 ;
        RECT 793.950 670.950 796.050 671.400 ;
        RECT 805.950 670.950 808.050 671.400 ;
        RECT 823.950 670.800 826.050 672.900 ;
        RECT 919.950 672.600 922.050 673.050 ;
        RECT 928.950 672.600 931.050 673.050 ;
        RECT 919.950 671.400 931.050 672.600 ;
        RECT 919.950 670.950 922.050 671.400 ;
        RECT 928.950 670.950 931.050 671.400 ;
        RECT 946.950 672.600 949.050 673.050 ;
        RECT 952.950 672.600 955.050 672.900 ;
        RECT 946.950 671.400 955.050 672.600 ;
        RECT 946.950 670.950 949.050 671.400 ;
        RECT 952.950 670.800 955.050 671.400 ;
        RECT 964.950 672.600 967.050 673.050 ;
        RECT 982.950 672.600 985.050 673.050 ;
        RECT 964.950 671.400 985.050 672.600 ;
        RECT 964.950 670.950 967.050 671.400 ;
        RECT 982.950 670.950 985.050 671.400 ;
        RECT 580.950 669.600 583.050 670.050 ;
        RECT 628.950 669.600 631.050 670.050 ;
        RECT 580.950 668.400 631.050 669.600 ;
        RECT 580.950 667.950 583.050 668.400 ;
        RECT 628.950 667.950 631.050 668.400 ;
        RECT 670.950 669.600 673.050 670.050 ;
        RECT 679.950 669.600 682.050 670.050 ;
        RECT 670.950 668.400 682.050 669.600 ;
        RECT 670.950 667.950 673.050 668.400 ;
        RECT 679.950 667.950 682.050 668.400 ;
        RECT 709.950 669.600 712.050 670.050 ;
        RECT 739.800 669.600 741.900 669.900 ;
        RECT 709.950 668.400 741.900 669.600 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 739.800 667.800 741.900 668.400 ;
        RECT 742.950 669.600 745.050 670.050 ;
        RECT 754.950 669.600 757.050 670.050 ;
        RECT 742.950 668.400 757.050 669.600 ;
        RECT 742.950 667.950 745.050 668.400 ;
        RECT 754.950 667.950 757.050 668.400 ;
        RECT 820.950 669.600 823.050 670.050 ;
        RECT 868.800 669.600 870.900 669.900 ;
        RECT 820.950 668.400 870.900 669.600 ;
        RECT 820.950 667.950 823.050 668.400 ;
        RECT 868.800 667.800 870.900 668.400 ;
        RECT 871.950 669.600 874.050 670.050 ;
        RECT 931.950 669.600 934.050 670.050 ;
        RECT 871.950 668.400 934.050 669.600 ;
        RECT 871.950 667.950 874.050 668.400 ;
        RECT 931.950 667.950 934.050 668.400 ;
        RECT 940.950 669.600 943.050 670.050 ;
        RECT 970.950 669.600 973.050 670.050 ;
        RECT 940.950 668.400 973.050 669.600 ;
        RECT 940.950 667.950 943.050 668.400 ;
        RECT 970.950 667.950 973.050 668.400 ;
        RECT 1003.950 669.600 1006.050 670.050 ;
        RECT 1018.950 669.600 1021.050 670.050 ;
        RECT 1003.950 668.400 1021.050 669.600 ;
        RECT 1003.950 667.950 1006.050 668.400 ;
        RECT 1018.950 667.950 1021.050 668.400 ;
        RECT 148.950 666.600 151.050 667.050 ;
        RECT 172.950 666.600 175.050 667.050 ;
        RECT 148.950 665.400 175.050 666.600 ;
        RECT 148.950 664.950 151.050 665.400 ;
        RECT 172.950 664.950 175.050 665.400 ;
        RECT 364.950 666.600 367.050 667.050 ;
        RECT 379.950 666.600 382.050 667.050 ;
        RECT 445.950 666.600 448.050 667.050 ;
        RECT 364.950 665.400 448.050 666.600 ;
        RECT 364.950 664.950 367.050 665.400 ;
        RECT 379.950 664.950 382.050 665.400 ;
        RECT 445.950 664.950 448.050 665.400 ;
        RECT 568.950 666.600 571.050 667.050 ;
        RECT 604.950 666.600 607.050 667.050 ;
        RECT 568.950 665.400 607.050 666.600 ;
        RECT 568.950 664.950 571.050 665.400 ;
        RECT 604.950 664.950 607.050 665.400 ;
        RECT 622.950 666.600 625.050 667.050 ;
        RECT 643.950 666.600 646.050 667.050 ;
        RECT 622.950 665.400 646.050 666.600 ;
        RECT 622.950 664.950 625.050 665.400 ;
        RECT 643.950 664.950 646.050 665.400 ;
        RECT 682.950 666.600 685.050 667.050 ;
        RECT 721.800 666.600 723.900 667.050 ;
        RECT 682.950 665.400 723.900 666.600 ;
        RECT 682.950 664.950 685.050 665.400 ;
        RECT 721.800 664.950 723.900 665.400 ;
        RECT 724.950 666.600 727.050 667.050 ;
        RECT 733.950 666.600 736.050 667.050 ;
        RECT 724.950 665.400 736.050 666.600 ;
        RECT 724.950 664.950 727.050 665.400 ;
        RECT 733.950 664.950 736.050 665.400 ;
        RECT 814.950 666.600 817.050 667.050 ;
        RECT 862.950 666.600 865.050 667.050 ;
        RECT 814.950 665.400 865.050 666.600 ;
        RECT 814.950 664.950 817.050 665.400 ;
        RECT 862.950 664.950 865.050 665.400 ;
        RECT 916.950 666.600 919.050 667.050 ;
        RECT 934.950 666.600 937.050 667.050 ;
        RECT 973.950 666.600 976.050 667.050 ;
        RECT 994.950 666.600 997.050 667.050 ;
        RECT 916.950 665.400 997.050 666.600 ;
        RECT 916.950 664.950 919.050 665.400 ;
        RECT 934.950 664.950 937.050 665.400 ;
        RECT 973.950 664.950 976.050 665.400 ;
        RECT 994.950 664.950 997.050 665.400 ;
        RECT 334.950 663.600 337.050 664.050 ;
        RECT 460.950 663.600 463.050 664.050 ;
        RECT 334.950 662.400 463.050 663.600 ;
        RECT 334.950 661.950 337.050 662.400 ;
        RECT 460.950 661.950 463.050 662.400 ;
        RECT 493.950 663.600 496.050 664.050 ;
        RECT 514.950 663.600 517.050 664.050 ;
        RECT 544.950 663.600 547.050 664.050 ;
        RECT 493.950 662.400 547.050 663.600 ;
        RECT 493.950 661.950 496.050 662.400 ;
        RECT 514.950 661.950 517.050 662.400 ;
        RECT 544.950 661.950 547.050 662.400 ;
        RECT 553.950 663.600 556.050 664.050 ;
        RECT 601.950 663.600 604.050 664.050 ;
        RECT 553.950 662.400 604.050 663.600 ;
        RECT 553.950 661.950 556.050 662.400 ;
        RECT 601.950 661.950 604.050 662.400 ;
        RECT 631.950 663.600 634.050 664.050 ;
        RECT 679.950 663.600 682.050 664.050 ;
        RECT 742.950 663.600 745.050 664.050 ;
        RECT 631.950 662.400 682.050 663.600 ;
        RECT 631.950 661.950 634.050 662.400 ;
        RECT 679.950 661.950 682.050 662.400 ;
        RECT 722.400 662.400 745.050 663.600 ;
        RECT 34.950 660.600 37.050 661.050 ;
        RECT 46.950 660.600 49.050 661.050 ;
        RECT 34.950 659.400 49.050 660.600 ;
        RECT 34.950 658.950 37.050 659.400 ;
        RECT 46.950 658.950 49.050 659.400 ;
        RECT 310.950 660.600 313.050 661.050 ;
        RECT 319.950 660.600 322.050 661.050 ;
        RECT 310.950 659.400 322.050 660.600 ;
        RECT 310.950 658.950 313.050 659.400 ;
        RECT 319.950 658.950 322.050 659.400 ;
        RECT 379.950 660.600 382.050 661.050 ;
        RECT 466.950 660.600 469.050 661.050 ;
        RECT 478.950 660.600 481.050 661.050 ;
        RECT 496.950 660.600 499.050 661.050 ;
        RECT 589.950 660.600 592.050 661.050 ;
        RECT 379.950 659.400 592.050 660.600 ;
        RECT 379.950 658.950 382.050 659.400 ;
        RECT 466.950 658.950 469.050 659.400 ;
        RECT 478.950 658.950 481.050 659.400 ;
        RECT 496.950 658.950 499.050 659.400 ;
        RECT 589.950 658.950 592.050 659.400 ;
        RECT 616.950 660.600 619.050 661.050 ;
        RECT 676.950 660.600 679.050 661.050 ;
        RECT 616.950 659.400 679.050 660.600 ;
        RECT 616.950 658.950 619.050 659.400 ;
        RECT 676.950 658.950 679.050 659.400 ;
        RECT 682.950 660.600 685.050 661.050 ;
        RECT 722.400 660.600 723.600 662.400 ;
        RECT 742.950 661.950 745.050 662.400 ;
        RECT 748.950 663.600 751.050 664.050 ;
        RECT 760.950 663.600 763.050 664.050 ;
        RECT 748.950 662.400 763.050 663.600 ;
        RECT 748.950 661.950 751.050 662.400 ;
        RECT 760.950 661.950 763.050 662.400 ;
        RECT 796.950 663.600 799.050 664.050 ;
        RECT 883.950 663.600 886.050 664.050 ;
        RECT 796.950 662.400 886.050 663.600 ;
        RECT 796.950 661.950 799.050 662.400 ;
        RECT 883.950 661.950 886.050 662.400 ;
        RECT 895.950 663.600 898.050 664.050 ;
        RECT 982.950 663.600 985.050 664.050 ;
        RECT 895.950 662.400 985.050 663.600 ;
        RECT 895.950 661.950 898.050 662.400 ;
        RECT 982.950 661.950 985.050 662.400 ;
        RECT 682.950 659.400 723.600 660.600 ;
        RECT 724.950 660.600 727.050 661.050 ;
        RECT 733.950 660.600 736.050 661.050 ;
        RECT 724.950 659.400 736.050 660.600 ;
        RECT 682.950 658.950 685.050 659.400 ;
        RECT 724.950 658.950 727.050 659.400 ;
        RECT 733.950 658.950 736.050 659.400 ;
        RECT 739.950 660.600 742.050 661.050 ;
        RECT 775.950 660.600 778.050 661.050 ;
        RECT 790.950 660.600 793.050 661.050 ;
        RECT 739.950 659.400 793.050 660.600 ;
        RECT 739.950 658.950 742.050 659.400 ;
        RECT 775.950 658.950 778.050 659.400 ;
        RECT 790.950 658.950 793.050 659.400 ;
        RECT 826.950 660.600 829.050 661.050 ;
        RECT 835.950 660.600 838.050 661.050 ;
        RECT 826.950 659.400 838.050 660.600 ;
        RECT 826.950 658.950 829.050 659.400 ;
        RECT 835.950 658.950 838.050 659.400 ;
        RECT 853.950 660.600 856.050 661.050 ;
        RECT 877.950 660.600 880.050 661.050 ;
        RECT 853.950 659.400 880.050 660.600 ;
        RECT 853.950 658.950 856.050 659.400 ;
        RECT 877.950 658.950 880.050 659.400 ;
        RECT 916.950 660.600 919.050 661.050 ;
        RECT 934.950 660.600 937.050 661.050 ;
        RECT 940.950 660.600 943.050 661.050 ;
        RECT 916.950 659.400 943.050 660.600 ;
        RECT 916.950 658.950 919.050 659.400 ;
        RECT 934.950 658.950 937.050 659.400 ;
        RECT 940.950 658.950 943.050 659.400 ;
        RECT 946.950 660.600 949.050 661.050 ;
        RECT 976.950 660.600 979.050 661.050 ;
        RECT 946.950 659.400 979.050 660.600 ;
        RECT 946.950 658.950 949.050 659.400 ;
        RECT 976.950 658.950 979.050 659.400 ;
        RECT 994.950 660.600 997.050 661.050 ;
        RECT 1033.950 660.600 1036.050 661.050 ;
        RECT 994.950 659.400 1036.050 660.600 ;
        RECT 994.950 658.950 997.050 659.400 ;
        RECT 1033.950 658.950 1036.050 659.400 ;
        RECT 178.950 657.600 181.050 658.050 ;
        RECT 190.950 657.600 193.050 658.050 ;
        RECT 178.950 656.400 193.050 657.600 ;
        RECT 178.950 655.950 181.050 656.400 ;
        RECT 190.950 655.950 193.050 656.400 ;
        RECT 223.950 657.600 226.050 658.050 ;
        RECT 238.950 657.600 241.050 658.050 ;
        RECT 223.950 656.400 241.050 657.600 ;
        RECT 223.950 655.950 226.050 656.400 ;
        RECT 238.950 655.950 241.050 656.400 ;
        RECT 292.950 657.600 295.050 658.050 ;
        RECT 328.950 657.600 331.050 658.050 ;
        RECT 292.950 656.400 331.050 657.600 ;
        RECT 292.950 655.950 295.050 656.400 ;
        RECT 328.950 655.950 331.050 656.400 ;
        RECT 409.950 657.600 412.050 658.050 ;
        RECT 418.950 657.600 421.050 658.050 ;
        RECT 409.950 656.400 421.050 657.600 ;
        RECT 409.950 655.950 412.050 656.400 ;
        RECT 418.950 655.950 421.050 656.400 ;
        RECT 439.950 657.600 442.050 658.050 ;
        RECT 454.950 657.600 457.050 658.050 ;
        RECT 613.950 657.600 616.050 658.050 ;
        RECT 721.950 657.600 724.050 658.050 ;
        RECT 736.950 657.600 739.050 658.050 ;
        RECT 439.950 656.400 462.600 657.600 ;
        RECT 439.950 655.950 442.050 656.400 ;
        RECT 454.950 655.950 457.050 656.400 ;
        RECT 244.950 654.600 247.050 655.050 ;
        RECT 400.950 654.600 403.050 655.050 ;
        RECT 406.950 654.600 409.050 655.050 ;
        RECT 244.950 653.400 348.600 654.600 ;
        RECT 244.950 652.950 247.050 653.400 ;
        RECT 16.950 650.100 19.050 652.200 ;
        RECT 22.950 651.750 25.050 652.200 ;
        RECT 28.950 651.750 31.050 652.200 ;
        RECT 22.950 651.600 31.050 651.750 ;
        RECT 40.950 651.600 43.050 652.200 ;
        RECT 73.950 651.600 76.050 652.050 ;
        RECT 22.950 650.550 76.050 651.600 ;
        RECT 22.950 650.100 25.050 650.550 ;
        RECT 28.950 650.400 76.050 650.550 ;
        RECT 28.950 650.100 31.050 650.400 ;
        RECT 40.950 650.100 43.050 650.400 ;
        RECT 17.400 648.600 18.600 650.100 ;
        RECT 73.950 649.950 76.050 650.400 ;
        RECT 85.950 651.600 88.050 652.050 ;
        RECT 94.950 651.600 97.050 652.050 ;
        RECT 85.950 650.400 97.050 651.600 ;
        RECT 85.950 649.950 88.050 650.400 ;
        RECT 94.950 649.950 97.050 650.400 ;
        RECT 172.950 651.750 175.050 652.200 ;
        RECT 184.950 651.750 187.050 652.200 ;
        RECT 172.950 650.550 187.050 651.750 ;
        RECT 172.950 650.100 175.050 650.550 ;
        RECT 184.950 650.100 187.050 650.550 ;
        RECT 202.950 651.750 205.050 652.200 ;
        RECT 211.950 651.750 214.050 652.200 ;
        RECT 202.950 650.550 214.050 651.750 ;
        RECT 202.950 650.100 205.050 650.550 ;
        RECT 211.950 650.100 214.050 650.550 ;
        RECT 220.950 651.600 223.050 652.050 ;
        RECT 220.950 650.400 228.600 651.600 ;
        RECT 220.950 649.950 223.050 650.400 ;
        RECT 148.950 648.600 151.050 649.200 ;
        RECT 17.400 647.400 39.600 648.600 ;
        RECT 10.950 645.600 13.050 646.050 ;
        RECT 38.400 645.900 39.600 647.400 ;
        RECT 80.400 647.400 151.050 648.600 ;
        RECT 80.400 646.050 81.600 647.400 ;
        RECT 148.950 647.100 151.050 647.400 ;
        RECT 157.950 648.750 160.050 649.200 ;
        RECT 214.950 648.750 217.050 649.200 ;
        RECT 157.950 647.550 217.050 648.750 ;
        RECT 157.950 647.100 160.050 647.550 ;
        RECT 214.950 647.100 217.050 647.550 ;
        RECT 19.950 645.600 22.050 645.900 ;
        RECT 10.950 644.400 22.050 645.600 ;
        RECT 10.950 643.950 13.050 644.400 ;
        RECT 19.950 643.800 22.050 644.400 ;
        RECT 37.950 645.450 40.050 645.900 ;
        RECT 43.950 645.450 46.050 645.900 ;
        RECT 37.950 644.250 46.050 645.450 ;
        RECT 37.950 643.800 40.050 644.250 ;
        RECT 43.950 643.800 46.050 644.250 ;
        RECT 70.950 645.600 73.050 645.900 ;
        RECT 79.950 645.600 82.050 646.050 ;
        RECT 70.950 644.400 82.050 645.600 ;
        RECT 70.950 643.800 73.050 644.400 ;
        RECT 79.950 643.950 82.050 644.400 ;
        RECT 121.950 645.600 124.050 646.050 ;
        RECT 227.400 645.900 228.600 650.400 ;
        RECT 229.950 650.100 232.050 652.200 ;
        RECT 250.950 651.600 253.050 652.200 ;
        RECT 256.950 651.600 259.050 652.200 ;
        RECT 268.950 651.600 271.050 652.050 ;
        RECT 277.950 651.600 280.050 652.200 ;
        RECT 304.950 651.600 307.050 652.200 ;
        RECT 334.950 651.600 337.050 652.200 ;
        RECT 250.950 650.400 255.600 651.600 ;
        RECT 250.950 650.100 253.050 650.400 ;
        RECT 181.950 645.600 184.050 645.900 ;
        RECT 121.950 644.400 184.050 645.600 ;
        RECT 121.950 643.950 124.050 644.400 ;
        RECT 181.950 643.800 184.050 644.400 ;
        RECT 226.950 643.800 229.050 645.900 ;
        RECT 230.400 645.600 231.600 650.100 ;
        RECT 254.400 648.600 255.600 650.400 ;
        RECT 256.950 650.400 271.050 651.600 ;
        RECT 256.950 650.100 259.050 650.400 ;
        RECT 268.950 649.950 271.050 650.400 ;
        RECT 272.400 650.400 307.050 651.600 ;
        RECT 272.400 648.600 273.600 650.400 ;
        RECT 277.950 650.100 280.050 650.400 ;
        RECT 304.950 650.100 307.050 650.400 ;
        RECT 314.400 650.400 337.050 651.600 ;
        RECT 254.400 647.400 273.600 648.600 ;
        RECT 235.950 645.600 238.050 646.050 ;
        RECT 314.400 645.900 315.600 650.400 ;
        RECT 334.950 650.100 337.050 650.400 ;
        RECT 340.950 651.600 343.050 652.200 ;
        RECT 347.400 651.600 348.600 653.400 ;
        RECT 400.950 653.400 409.050 654.600 ;
        RECT 461.400 654.600 462.600 656.400 ;
        RECT 613.950 656.400 630.600 657.600 ;
        RECT 613.950 655.950 616.050 656.400 ;
        RECT 469.950 654.600 472.050 655.050 ;
        RECT 505.950 654.600 508.050 655.050 ;
        RECT 461.400 653.400 508.050 654.600 ;
        RECT 400.950 652.950 403.050 653.400 ;
        RECT 406.950 652.950 409.050 653.400 ;
        RECT 469.950 652.950 472.050 653.400 ;
        RECT 505.950 652.950 508.050 653.400 ;
        RECT 535.950 654.600 538.050 655.050 ;
        RECT 547.950 654.600 550.050 655.050 ;
        RECT 629.400 654.600 630.600 656.400 ;
        RECT 721.950 656.400 739.050 657.600 ;
        RECT 721.950 655.950 724.050 656.400 ;
        RECT 736.950 655.950 739.050 656.400 ;
        RECT 751.950 657.600 754.050 658.050 ;
        RECT 763.950 657.600 766.050 658.050 ;
        RECT 751.950 656.400 766.050 657.600 ;
        RECT 751.950 655.950 754.050 656.400 ;
        RECT 763.950 655.950 766.050 656.400 ;
        RECT 910.950 657.600 913.050 658.050 ;
        RECT 943.950 657.600 946.050 658.050 ;
        RECT 910.950 656.400 946.050 657.600 ;
        RECT 910.950 655.950 913.050 656.400 ;
        RECT 943.950 655.950 946.050 656.400 ;
        RECT 679.950 654.600 682.050 655.050 ;
        RECT 535.950 653.400 550.050 654.600 ;
        RECT 535.950 652.950 538.050 653.400 ;
        RECT 547.950 652.950 550.050 653.400 ;
        RECT 596.400 653.400 627.600 654.600 ;
        RECT 629.400 653.400 682.050 654.600 ;
        RECT 358.950 651.600 361.050 652.200 ;
        RECT 376.800 651.600 378.900 652.050 ;
        RECT 340.950 650.400 345.600 651.600 ;
        RECT 347.400 650.400 378.900 651.600 ;
        RECT 340.950 650.100 343.050 650.400 ;
        RECT 344.400 646.050 345.600 650.400 ;
        RECT 358.950 650.100 361.050 650.400 ;
        RECT 376.800 649.950 378.900 650.400 ;
        RECT 379.950 651.600 384.000 652.050 ;
        RECT 385.950 651.600 388.050 652.200 ;
        RECT 397.950 651.600 400.050 652.050 ;
        RECT 379.950 649.950 384.600 651.600 ;
        RECT 385.950 650.400 400.050 651.600 ;
        RECT 385.950 650.100 388.050 650.400 ;
        RECT 397.950 649.950 400.050 650.400 ;
        RECT 403.950 651.600 408.000 652.050 ;
        RECT 409.950 651.600 412.050 652.200 ;
        RECT 430.950 651.600 433.050 652.050 ;
        RECT 403.950 649.950 408.600 651.600 ;
        RECT 409.950 650.400 433.050 651.600 ;
        RECT 409.950 650.100 412.050 650.400 ;
        RECT 430.950 649.950 433.050 650.400 ;
        RECT 436.950 651.600 439.050 652.200 ;
        RECT 457.950 651.600 460.050 652.200 ;
        RECT 436.950 650.400 460.050 651.600 ;
        RECT 436.950 650.100 439.050 650.400 ;
        RECT 457.950 650.100 460.050 650.400 ;
        RECT 511.950 651.600 514.050 652.200 ;
        RECT 529.950 651.600 532.050 652.200 ;
        RECT 511.950 650.400 532.050 651.600 ;
        RECT 511.950 650.100 514.050 650.400 ;
        RECT 230.400 644.400 238.050 645.600 ;
        RECT 235.950 643.950 238.050 644.400 ;
        RECT 259.950 645.450 262.050 645.900 ;
        RECT 265.950 645.450 268.050 645.900 ;
        RECT 259.950 644.250 268.050 645.450 ;
        RECT 259.950 643.800 262.050 644.250 ;
        RECT 265.950 643.800 268.050 644.250 ;
        RECT 286.950 645.450 289.050 645.900 ;
        RECT 292.950 645.450 295.050 645.900 ;
        RECT 286.950 644.250 295.050 645.450 ;
        RECT 286.950 643.800 289.050 644.250 ;
        RECT 292.950 643.800 295.050 644.250 ;
        RECT 313.950 643.800 316.050 645.900 ;
        RECT 325.950 645.450 328.050 645.900 ;
        RECT 331.950 645.450 334.050 645.900 ;
        RECT 325.950 644.250 334.050 645.450 ;
        RECT 325.950 643.800 328.050 644.250 ;
        RECT 331.950 643.800 334.050 644.250 ;
        RECT 343.950 643.950 346.050 646.050 ;
        RECT 383.400 645.900 384.600 649.950 ;
        RECT 407.400 645.900 408.600 649.950 ;
        RECT 515.400 646.050 516.600 650.400 ;
        RECT 529.950 650.100 532.050 650.400 ;
        RECT 538.950 649.950 541.050 652.050 ;
        RECT 550.800 649.950 552.900 652.050 ;
        RECT 553.950 650.100 556.050 652.200 ;
        RECT 565.950 651.600 568.050 652.050 ;
        RECT 577.950 651.600 580.050 652.200 ;
        RECT 596.400 652.050 597.600 653.400 ;
        RECT 565.950 650.400 580.050 651.600 ;
        RECT 539.400 646.050 540.600 649.950 ;
        RECT 551.400 646.050 552.600 649.950 ;
        RECT 382.950 643.800 385.050 645.900 ;
        RECT 388.950 645.600 391.050 645.900 ;
        RECT 406.950 645.600 409.050 645.900 ;
        RECT 388.950 644.400 409.050 645.600 ;
        RECT 388.950 643.800 391.050 644.400 ;
        RECT 406.950 643.800 409.050 644.400 ;
        RECT 460.950 645.450 463.050 645.900 ;
        RECT 466.950 645.450 469.050 645.900 ;
        RECT 460.950 644.250 469.050 645.450 ;
        RECT 460.950 643.800 463.050 644.250 ;
        RECT 466.950 643.800 469.050 644.250 ;
        RECT 472.950 645.600 475.050 646.050 ;
        RECT 478.950 645.600 481.050 645.900 ;
        RECT 472.950 644.400 481.050 645.600 ;
        RECT 472.950 643.950 475.050 644.400 ;
        RECT 478.950 643.800 481.050 644.400 ;
        RECT 484.950 645.600 487.050 645.900 ;
        RECT 496.950 645.600 499.050 646.050 ;
        RECT 484.950 644.400 499.050 645.600 ;
        RECT 484.950 643.800 487.050 644.400 ;
        RECT 496.950 643.950 499.050 644.400 ;
        RECT 514.950 643.950 517.050 646.050 ;
        RECT 523.950 645.600 526.050 646.050 ;
        RECT 532.950 645.600 535.050 645.900 ;
        RECT 523.950 644.400 535.050 645.600 ;
        RECT 523.950 643.950 526.050 644.400 ;
        RECT 532.950 643.800 535.050 644.400 ;
        RECT 538.950 643.950 541.050 646.050 ;
        RECT 550.950 643.950 553.050 646.050 ;
        RECT 554.400 645.600 555.600 650.100 ;
        RECT 565.950 649.950 568.050 650.400 ;
        RECT 577.950 650.100 580.050 650.400 ;
        RECT 595.950 648.600 598.050 652.050 ;
        RECT 607.950 651.600 610.050 652.050 ;
        RECT 607.950 650.400 621.600 651.600 ;
        RECT 607.950 649.950 610.050 650.400 ;
        RECT 587.400 648.000 598.050 648.600 ;
        RECT 587.400 647.400 597.600 648.000 ;
        RECT 574.950 645.600 577.050 645.900 ;
        RECT 554.400 644.400 577.050 645.600 ;
        RECT 574.950 643.800 577.050 644.400 ;
        RECT 580.950 645.600 583.050 645.900 ;
        RECT 587.400 645.600 588.600 647.400 ;
        RECT 620.400 646.050 621.600 650.400 ;
        RECT 580.950 644.400 588.600 645.600 ;
        RECT 589.950 645.450 592.050 645.900 ;
        RECT 598.950 645.450 601.050 645.900 ;
        RECT 580.950 643.800 583.050 644.400 ;
        RECT 589.950 644.250 601.050 645.450 ;
        RECT 589.950 643.800 592.050 644.250 ;
        RECT 598.950 643.800 601.050 644.250 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 626.400 645.900 627.600 653.400 ;
        RECT 679.950 652.950 682.050 653.400 ;
        RECT 727.950 654.600 730.050 655.050 ;
        RECT 736.950 654.600 739.050 654.900 ;
        RECT 727.950 653.400 739.050 654.600 ;
        RECT 727.950 652.950 730.050 653.400 ;
        RECT 736.950 652.800 739.050 653.400 ;
        RECT 745.950 654.600 748.050 655.050 ;
        RECT 754.950 654.600 757.050 655.050 ;
        RECT 745.950 653.400 757.050 654.600 ;
        RECT 745.950 652.950 748.050 653.400 ;
        RECT 754.950 652.950 757.050 653.400 ;
        RECT 778.950 654.600 781.050 655.050 ;
        RECT 840.000 654.600 844.050 655.050 ;
        RECT 778.950 653.400 798.600 654.600 ;
        RECT 778.950 652.950 781.050 653.400 ;
        RECT 634.950 651.600 637.050 652.050 ;
        RECT 640.950 651.600 643.050 652.050 ;
        RECT 634.950 650.400 643.050 651.600 ;
        RECT 634.950 649.950 637.050 650.400 ;
        RECT 640.950 649.950 643.050 650.400 ;
        RECT 652.950 651.750 655.050 652.200 ;
        RECT 664.950 651.750 667.050 652.200 ;
        RECT 652.950 650.550 667.050 651.750 ;
        RECT 652.950 650.100 655.050 650.550 ;
        RECT 664.950 650.100 667.050 650.550 ;
        RECT 682.950 651.750 685.050 652.200 ;
        RECT 688.950 651.750 691.050 652.200 ;
        RECT 682.950 650.550 691.050 651.750 ;
        RECT 703.950 651.600 706.050 652.200 ;
        RECT 682.950 650.100 685.050 650.550 ;
        RECT 688.950 650.100 691.050 650.550 ;
        RECT 698.400 650.400 706.050 651.600 ;
        RECT 698.400 646.050 699.600 650.400 ;
        RECT 703.950 650.100 706.050 650.400 ;
        RECT 721.950 651.600 726.000 652.050 ;
        RECT 721.950 649.950 726.600 651.600 ;
        RECT 625.950 643.800 628.050 645.900 ;
        RECT 643.950 645.450 646.050 646.050 ;
        RECT 649.950 645.450 652.050 645.900 ;
        RECT 643.950 644.250 652.050 645.450 ;
        RECT 643.950 643.950 646.050 644.250 ;
        RECT 649.950 643.800 652.050 644.250 ;
        RECT 664.950 645.600 667.050 646.050 ;
        RECT 679.950 645.600 682.050 645.900 ;
        RECT 664.950 644.400 682.050 645.600 ;
        RECT 664.950 643.950 667.050 644.400 ;
        RECT 679.950 643.800 682.050 644.400 ;
        RECT 697.950 643.950 700.050 646.050 ;
        RECT 725.400 645.900 726.600 649.950 ;
        RECT 742.950 648.600 745.050 652.050 ;
        RECT 754.950 651.600 757.050 652.200 ;
        RECT 793.950 651.600 796.050 652.200 ;
        RECT 754.950 650.400 796.050 651.600 ;
        RECT 754.950 650.100 757.050 650.400 ;
        RECT 793.950 650.100 796.050 650.400 ;
        RECT 742.950 648.000 753.600 648.600 ;
        RECT 743.400 647.400 754.050 648.000 ;
        RECT 724.950 643.800 727.050 645.900 ;
        RECT 751.950 643.950 754.050 647.400 ;
        RECT 797.400 645.900 798.600 653.400 ;
        RECT 839.400 652.950 844.050 654.600 ;
        RECT 856.950 654.600 859.050 654.900 ;
        RECT 865.950 654.600 868.050 655.050 ;
        RECT 856.950 653.400 868.050 654.600 ;
        RECT 814.950 650.100 817.050 652.200 ;
        RECT 829.950 651.600 832.050 652.050 ;
        RECT 835.950 651.600 838.050 652.050 ;
        RECT 829.950 650.400 838.050 651.600 ;
        RECT 769.950 645.450 772.050 645.900 ;
        RECT 784.950 645.450 787.050 645.900 ;
        RECT 769.950 644.250 787.050 645.450 ;
        RECT 769.950 643.800 772.050 644.250 ;
        RECT 784.950 643.800 787.050 644.250 ;
        RECT 796.950 643.800 799.050 645.900 ;
        RECT 815.400 645.600 816.600 650.100 ;
        RECT 829.950 649.950 832.050 650.400 ;
        RECT 835.950 649.950 838.050 650.400 ;
        RECT 815.400 645.000 822.600 645.600 ;
        RECT 815.400 644.400 823.050 645.000 ;
        RECT 205.950 642.600 208.050 643.050 ;
        RECT 223.950 642.600 226.050 642.750 ;
        RECT 205.950 641.400 226.050 642.600 ;
        RECT 205.950 640.950 208.050 641.400 ;
        RECT 223.950 640.650 226.050 641.400 ;
        RECT 253.950 642.600 256.050 643.050 ;
        RECT 280.950 642.600 283.050 643.050 ;
        RECT 253.950 641.400 283.050 642.600 ;
        RECT 253.950 640.950 256.050 641.400 ;
        RECT 280.950 640.950 283.050 641.400 ;
        RECT 307.950 642.600 310.050 643.050 ;
        RECT 337.950 642.600 340.050 643.050 ;
        RECT 307.950 641.400 340.050 642.600 ;
        RECT 307.950 640.950 310.050 641.400 ;
        RECT 337.950 640.950 340.050 641.400 ;
        RECT 454.950 642.600 457.050 643.050 ;
        RECT 469.950 642.600 472.050 643.050 ;
        RECT 454.950 641.400 472.050 642.600 ;
        RECT 454.950 640.950 457.050 641.400 ;
        RECT 469.950 640.950 472.050 641.400 ;
        RECT 643.950 642.600 646.050 642.900 ;
        RECT 655.950 642.600 658.050 643.050 ;
        RECT 643.950 641.400 658.050 642.600 ;
        RECT 643.950 640.800 646.050 641.400 ;
        RECT 655.950 640.950 658.050 641.400 ;
        RECT 793.950 642.600 796.050 643.050 ;
        RECT 808.950 642.600 811.050 643.050 ;
        RECT 793.950 641.400 811.050 642.600 ;
        RECT 793.950 640.950 796.050 641.400 ;
        RECT 808.950 640.950 811.050 641.400 ;
        RECT 820.950 640.950 823.050 644.400 ;
        RECT 34.950 639.600 37.050 640.050 ;
        RECT 49.950 639.600 52.050 640.050 ;
        RECT 34.950 638.400 52.050 639.600 ;
        RECT 34.950 637.950 37.050 638.400 ;
        RECT 49.950 637.950 52.050 638.400 ;
        RECT 64.950 639.600 67.050 640.050 ;
        RECT 85.950 639.600 88.050 640.050 ;
        RECT 97.950 639.600 100.050 640.050 ;
        RECT 64.950 638.400 100.050 639.600 ;
        RECT 64.950 637.950 67.050 638.400 ;
        RECT 85.950 637.950 88.050 638.400 ;
        RECT 97.950 637.950 100.050 638.400 ;
        RECT 403.950 639.600 406.050 640.050 ;
        RECT 412.950 639.600 415.050 640.050 ;
        RECT 442.950 639.600 445.050 640.050 ;
        RECT 493.950 639.600 496.050 640.050 ;
        RECT 403.950 638.400 496.050 639.600 ;
        RECT 403.950 637.950 406.050 638.400 ;
        RECT 412.950 637.950 415.050 638.400 ;
        RECT 442.950 637.950 445.050 638.400 ;
        RECT 493.950 637.950 496.050 638.400 ;
        RECT 508.950 639.600 511.050 640.050 ;
        RECT 520.800 639.600 522.900 640.050 ;
        RECT 508.950 638.400 522.900 639.600 ;
        RECT 508.950 637.950 511.050 638.400 ;
        RECT 520.800 637.950 522.900 638.400 ;
        RECT 523.950 639.600 526.050 640.050 ;
        RECT 646.950 639.600 649.050 640.050 ;
        RECT 523.950 638.400 649.050 639.600 ;
        RECT 523.950 637.950 526.050 638.400 ;
        RECT 646.950 637.950 649.050 638.400 ;
        RECT 688.950 639.600 691.050 640.050 ;
        RECT 709.950 639.600 712.050 640.050 ;
        RECT 688.950 638.400 712.050 639.600 ;
        RECT 688.950 637.950 691.050 638.400 ;
        RECT 709.950 637.950 712.050 638.400 ;
        RECT 760.950 639.600 763.050 640.050 ;
        RECT 778.950 639.600 781.050 640.050 ;
        RECT 760.950 638.400 781.050 639.600 ;
        RECT 760.950 637.950 763.050 638.400 ;
        RECT 778.950 637.950 781.050 638.400 ;
        RECT 796.950 639.600 799.050 640.050 ;
        RECT 817.950 639.600 820.050 640.050 ;
        RECT 796.950 638.400 820.050 639.600 ;
        RECT 839.400 639.600 840.600 652.950 ;
        RECT 856.950 652.800 859.050 653.400 ;
        RECT 865.950 652.950 868.050 653.400 ;
        RECT 886.950 654.600 889.050 654.900 ;
        RECT 892.950 654.600 895.050 655.050 ;
        RECT 886.950 653.400 895.050 654.600 ;
        RECT 886.950 652.800 889.050 653.400 ;
        RECT 892.950 652.950 895.050 653.400 ;
        RECT 883.950 651.600 886.050 652.050 ;
        RECT 895.950 651.600 898.050 652.200 ;
        RECT 883.950 650.400 898.050 651.600 ;
        RECT 883.950 649.950 886.050 650.400 ;
        RECT 895.950 650.100 898.050 650.400 ;
        RECT 907.950 651.600 910.050 652.050 ;
        RECT 913.950 651.600 916.050 652.050 ;
        RECT 907.950 650.400 916.050 651.600 ;
        RECT 907.950 649.950 910.050 650.400 ;
        RECT 913.950 649.950 916.050 650.400 ;
        RECT 931.950 651.600 936.000 652.050 ;
        RECT 949.950 651.600 952.050 652.050 ;
        RECT 970.950 651.600 973.050 652.200 ;
        RECT 931.950 649.950 936.600 651.600 ;
        RECT 949.950 650.400 973.050 651.600 ;
        RECT 949.950 649.950 952.050 650.400 ;
        RECT 970.950 650.100 973.050 650.400 ;
        RECT 994.950 650.100 997.050 652.200 ;
        RECT 880.950 648.600 883.050 649.050 ;
        RECT 842.400 647.400 883.050 648.600 ;
        RECT 935.400 648.600 936.600 649.950 ;
        RECT 935.400 647.400 957.600 648.600 ;
        RECT 842.400 645.900 843.600 647.400 ;
        RECT 880.950 646.950 883.050 647.400 ;
        RECT 841.950 643.800 844.050 645.900 ;
        RECT 913.950 645.600 916.050 646.050 ;
        RECT 925.950 645.600 928.050 646.050 ;
        RECT 913.950 644.400 928.050 645.600 ;
        RECT 913.950 643.950 916.050 644.400 ;
        RECT 925.950 643.950 928.050 644.400 ;
        RECT 946.950 645.600 949.050 645.900 ;
        RECT 952.950 645.600 955.050 646.050 ;
        RECT 946.950 644.400 955.050 645.600 ;
        RECT 946.950 643.800 949.050 644.400 ;
        RECT 952.950 643.950 955.050 644.400 ;
        RECT 886.950 642.600 889.050 643.050 ;
        RECT 898.950 642.600 901.050 643.050 ;
        RECT 886.950 641.400 901.050 642.600 ;
        RECT 886.950 640.950 889.050 641.400 ;
        RECT 898.950 640.950 901.050 641.400 ;
        RECT 931.950 642.600 934.050 642.900 ;
        RECT 946.950 642.600 949.050 643.050 ;
        RECT 931.950 641.400 949.050 642.600 ;
        RECT 956.400 642.600 957.600 647.400 ;
        RECT 971.400 646.050 972.600 650.100 ;
        RECT 971.400 644.400 976.050 646.050 ;
        RECT 972.000 643.950 976.050 644.400 ;
        RECT 964.950 642.600 967.050 643.050 ;
        RECT 956.400 641.400 967.050 642.600 ;
        RECT 931.950 640.800 934.050 641.400 ;
        RECT 946.950 640.950 949.050 641.400 ;
        RECT 964.950 640.950 967.050 641.400 ;
        RECT 988.950 642.600 991.050 643.050 ;
        RECT 995.400 642.600 996.600 650.100 ;
        RECT 988.950 641.400 996.600 642.600 ;
        RECT 988.950 640.950 991.050 641.400 ;
        RECT 844.950 639.600 847.050 640.050 ;
        RECT 839.400 638.400 847.050 639.600 ;
        RECT 796.950 637.950 799.050 638.400 ;
        RECT 817.950 637.950 820.050 638.400 ;
        RECT 844.950 637.950 847.050 638.400 ;
        RECT 889.950 639.600 892.050 640.050 ;
        RECT 895.950 639.600 898.050 640.050 ;
        RECT 889.950 638.400 898.050 639.600 ;
        RECT 889.950 637.950 892.050 638.400 ;
        RECT 895.950 637.950 898.050 638.400 ;
        RECT 211.950 636.600 214.050 637.050 ;
        RECT 235.950 636.600 238.050 637.050 ;
        RECT 310.950 636.600 313.050 637.050 ;
        RECT 343.950 636.600 346.050 637.050 ;
        RECT 211.950 635.400 346.050 636.600 ;
        RECT 211.950 634.950 214.050 635.400 ;
        RECT 235.950 634.950 238.050 635.400 ;
        RECT 310.950 634.950 313.050 635.400 ;
        RECT 343.950 634.950 346.050 635.400 ;
        RECT 448.950 636.600 451.050 637.050 ;
        RECT 457.950 636.600 460.050 637.050 ;
        RECT 448.950 635.400 460.050 636.600 ;
        RECT 448.950 634.950 451.050 635.400 ;
        RECT 457.950 634.950 460.050 635.400 ;
        RECT 481.950 636.600 484.050 637.050 ;
        RECT 502.950 636.600 505.050 637.050 ;
        RECT 481.950 635.400 505.050 636.600 ;
        RECT 481.950 634.950 484.050 635.400 ;
        RECT 502.950 634.950 505.050 635.400 ;
        RECT 547.950 636.600 550.050 637.050 ;
        RECT 556.950 636.600 559.050 637.050 ;
        RECT 616.950 636.600 619.050 637.050 ;
        RECT 547.950 635.400 619.050 636.600 ;
        RECT 547.950 634.950 550.050 635.400 ;
        RECT 556.950 634.950 559.050 635.400 ;
        RECT 616.950 634.950 619.050 635.400 ;
        RECT 631.950 636.600 634.050 637.050 ;
        RECT 706.950 636.600 709.050 637.050 ;
        RECT 631.950 635.400 709.050 636.600 ;
        RECT 631.950 634.950 634.050 635.400 ;
        RECT 706.950 634.950 709.050 635.400 ;
        RECT 712.950 636.600 715.050 636.900 ;
        RECT 766.950 636.600 769.050 637.050 ;
        RECT 712.950 635.400 769.050 636.600 ;
        RECT 712.950 634.800 715.050 635.400 ;
        RECT 766.950 634.950 769.050 635.400 ;
        RECT 784.950 636.600 787.050 637.050 ;
        RECT 862.950 636.600 865.050 637.050 ;
        RECT 784.950 635.400 865.050 636.600 ;
        RECT 784.950 634.950 787.050 635.400 ;
        RECT 862.950 634.950 865.050 635.400 ;
        RECT 889.950 636.600 892.050 636.900 ;
        RECT 901.950 636.600 904.050 640.050 ;
        RECT 940.950 639.600 943.050 639.900 ;
        RECT 955.950 639.600 958.050 640.050 ;
        RECT 940.950 638.400 958.050 639.600 ;
        RECT 940.950 637.800 943.050 638.400 ;
        RECT 955.950 637.950 958.050 638.400 ;
        RECT 967.950 639.600 970.050 640.050 ;
        RECT 973.950 639.600 976.050 640.050 ;
        RECT 967.950 638.400 976.050 639.600 ;
        RECT 967.950 637.950 970.050 638.400 ;
        RECT 973.950 637.950 976.050 638.400 ;
        RECT 889.950 636.000 904.050 636.600 ;
        RECT 904.950 636.600 907.050 637.050 ;
        RECT 922.950 636.600 925.050 637.050 ;
        RECT 889.950 635.400 903.600 636.000 ;
        RECT 904.950 635.400 925.050 636.600 ;
        RECT 889.950 634.800 892.050 635.400 ;
        RECT 904.950 634.950 907.050 635.400 ;
        RECT 922.950 634.950 925.050 635.400 ;
        RECT 991.950 636.600 994.050 637.050 ;
        RECT 1012.950 636.600 1015.050 637.050 ;
        RECT 991.950 635.400 1015.050 636.600 ;
        RECT 991.950 634.950 994.050 635.400 ;
        RECT 1012.950 634.950 1015.050 635.400 ;
        RECT 160.950 633.600 163.050 634.050 ;
        RECT 181.950 633.600 184.050 634.050 ;
        RECT 160.950 632.400 184.050 633.600 ;
        RECT 160.950 631.950 163.050 632.400 ;
        RECT 181.950 631.950 184.050 632.400 ;
        RECT 232.950 633.600 235.050 634.050 ;
        RECT 325.950 633.600 328.050 634.050 ;
        RECT 232.950 632.400 328.050 633.600 ;
        RECT 232.950 631.950 235.050 632.400 ;
        RECT 325.950 631.950 328.050 632.400 ;
        RECT 589.950 633.600 592.050 634.050 ;
        RECT 610.950 633.600 613.050 634.050 ;
        RECT 589.950 632.400 613.050 633.600 ;
        RECT 589.950 631.950 592.050 632.400 ;
        RECT 610.950 631.950 613.050 632.400 ;
        RECT 715.950 633.600 718.050 634.050 ;
        RECT 769.950 633.600 772.050 634.050 ;
        RECT 715.950 632.400 772.050 633.600 ;
        RECT 715.950 631.950 718.050 632.400 ;
        RECT 769.950 631.950 772.050 632.400 ;
        RECT 796.950 633.600 799.050 634.050 ;
        RECT 890.400 633.600 891.600 634.800 ;
        RECT 796.950 632.400 891.600 633.600 ;
        RECT 964.950 633.600 967.050 634.050 ;
        RECT 973.950 633.600 976.050 634.050 ;
        RECT 964.950 632.400 976.050 633.600 ;
        RECT 796.950 631.950 799.050 632.400 ;
        RECT 964.950 631.950 967.050 632.400 ;
        RECT 973.950 631.950 976.050 632.400 ;
        RECT 79.950 630.600 82.050 631.050 ;
        RECT 127.950 630.600 130.050 631.050 ;
        RECT 79.950 629.400 130.050 630.600 ;
        RECT 79.950 628.950 82.050 629.400 ;
        RECT 127.950 628.950 130.050 629.400 ;
        RECT 214.950 630.600 217.050 631.050 ;
        RECT 253.950 630.600 256.050 631.050 ;
        RECT 214.950 629.400 256.050 630.600 ;
        RECT 214.950 628.950 217.050 629.400 ;
        RECT 253.950 628.950 256.050 629.400 ;
        RECT 466.950 630.600 469.050 631.050 ;
        RECT 514.950 630.600 517.050 631.050 ;
        RECT 466.950 629.400 517.050 630.600 ;
        RECT 466.950 628.950 469.050 629.400 ;
        RECT 514.950 628.950 517.050 629.400 ;
        RECT 520.950 630.600 523.050 631.050 ;
        RECT 565.950 630.600 568.050 631.050 ;
        RECT 520.950 629.400 568.050 630.600 ;
        RECT 520.950 628.950 523.050 629.400 ;
        RECT 565.950 628.950 568.050 629.400 ;
        RECT 571.950 630.600 574.050 631.050 ;
        RECT 697.950 630.600 700.050 631.050 ;
        RECT 772.950 630.600 775.050 631.050 ;
        RECT 571.950 629.400 700.050 630.600 ;
        RECT 571.950 628.950 574.050 629.400 ;
        RECT 697.950 628.950 700.050 629.400 ;
        RECT 701.400 629.400 775.050 630.600 ;
        RECT 130.950 627.600 133.050 628.050 ;
        RECT 331.950 627.600 334.050 628.050 ;
        RECT 373.950 627.600 376.050 628.050 ;
        RECT 130.950 626.400 159.600 627.600 ;
        RECT 130.950 625.950 133.050 626.400 ;
        RECT 158.400 624.600 159.600 626.400 ;
        RECT 331.950 626.400 376.050 627.600 ;
        RECT 331.950 625.950 334.050 626.400 ;
        RECT 373.950 625.950 376.050 626.400 ;
        RECT 511.950 627.600 514.050 628.050 ;
        RECT 517.950 627.600 520.050 628.050 ;
        RECT 511.950 626.400 520.050 627.600 ;
        RECT 511.950 625.950 514.050 626.400 ;
        RECT 517.950 625.950 520.050 626.400 ;
        RECT 592.950 627.600 595.050 628.050 ;
        RECT 610.950 627.600 613.050 628.050 ;
        RECT 592.950 626.400 613.050 627.600 ;
        RECT 592.950 625.950 595.050 626.400 ;
        RECT 610.950 625.950 613.050 626.400 ;
        RECT 679.950 627.600 682.050 628.050 ;
        RECT 701.400 627.600 702.600 629.400 ;
        RECT 772.950 628.950 775.050 629.400 ;
        RECT 778.950 630.600 781.050 631.050 ;
        RECT 850.950 630.600 853.050 631.050 ;
        RECT 778.950 629.400 853.050 630.600 ;
        RECT 778.950 628.950 781.050 629.400 ;
        RECT 850.950 628.950 853.050 629.400 ;
        RECT 910.950 630.600 913.050 631.050 ;
        RECT 916.950 630.600 919.050 631.050 ;
        RECT 910.950 629.400 919.050 630.600 ;
        RECT 910.950 628.950 913.050 629.400 ;
        RECT 916.950 628.950 919.050 629.400 ;
        RECT 934.950 630.600 937.050 631.050 ;
        RECT 955.950 630.600 958.050 631.050 ;
        RECT 934.950 629.400 958.050 630.600 ;
        RECT 934.950 628.950 937.050 629.400 ;
        RECT 955.950 628.950 958.050 629.400 ;
        RECT 961.950 630.600 964.050 631.050 ;
        RECT 1012.950 630.600 1015.050 631.050 ;
        RECT 961.950 629.400 1015.050 630.600 ;
        RECT 961.950 628.950 964.050 629.400 ;
        RECT 1012.950 628.950 1015.050 629.400 ;
        RECT 718.950 627.600 721.050 628.050 ;
        RECT 679.950 626.400 702.600 627.600 ;
        RECT 704.400 626.400 721.050 627.600 ;
        RECT 679.950 625.950 682.050 626.400 ;
        RECT 172.950 624.600 175.050 625.050 ;
        RECT 158.400 623.400 175.050 624.600 ;
        RECT 172.950 622.950 175.050 623.400 ;
        RECT 325.950 624.600 328.050 625.050 ;
        RECT 394.950 624.600 397.050 625.050 ;
        RECT 613.950 624.600 616.050 625.050 ;
        RECT 325.950 623.400 397.050 624.600 ;
        RECT 325.950 622.950 328.050 623.400 ;
        RECT 394.950 622.950 397.050 623.400 ;
        RECT 485.400 623.400 616.050 624.600 ;
        RECT 124.950 621.600 127.050 622.050 ;
        RECT 151.950 621.600 154.050 622.050 ;
        RECT 124.950 620.400 154.050 621.600 ;
        RECT 124.950 619.950 127.050 620.400 ;
        RECT 151.950 619.950 154.050 620.400 ;
        RECT 376.950 621.600 379.050 622.050 ;
        RECT 439.950 621.600 442.050 622.050 ;
        RECT 376.950 620.400 442.050 621.600 ;
        RECT 376.950 619.950 379.050 620.400 ;
        RECT 439.950 619.950 442.050 620.400 ;
        RECT 478.950 621.600 481.050 622.050 ;
        RECT 485.400 621.600 486.600 623.400 ;
        RECT 613.950 622.950 616.050 623.400 ;
        RECT 628.950 624.600 631.050 625.050 ;
        RECT 658.950 624.600 661.050 625.050 ;
        RECT 676.950 624.600 679.050 625.050 ;
        RECT 704.400 624.600 705.600 626.400 ;
        RECT 718.950 625.950 721.050 626.400 ;
        RECT 727.950 627.600 730.050 628.050 ;
        RECT 802.950 627.600 805.050 628.050 ;
        RECT 727.950 626.400 805.050 627.600 ;
        RECT 727.950 625.950 730.050 626.400 ;
        RECT 802.950 625.950 805.050 626.400 ;
        RECT 844.950 627.600 847.050 628.050 ;
        RECT 874.950 627.600 877.050 628.050 ;
        RECT 844.950 626.400 877.050 627.600 ;
        RECT 844.950 625.950 847.050 626.400 ;
        RECT 874.950 625.950 877.050 626.400 ;
        RECT 892.950 627.600 895.050 628.050 ;
        RECT 928.950 627.600 931.050 628.050 ;
        RECT 949.950 627.600 952.050 628.050 ;
        RECT 892.950 626.400 952.050 627.600 ;
        RECT 892.950 625.950 895.050 626.400 ;
        RECT 928.950 625.950 931.050 626.400 ;
        RECT 949.950 625.950 952.050 626.400 ;
        RECT 628.950 623.400 645.600 624.600 ;
        RECT 628.950 622.950 631.050 623.400 ;
        RECT 478.950 620.400 486.600 621.600 ;
        RECT 544.950 621.600 547.050 622.050 ;
        RECT 640.950 621.600 643.050 622.050 ;
        RECT 544.950 620.400 643.050 621.600 ;
        RECT 644.400 621.600 645.600 623.400 ;
        RECT 658.950 623.400 705.600 624.600 ;
        RECT 709.950 624.600 712.050 625.050 ;
        RECT 847.950 624.600 850.050 625.050 ;
        RECT 853.950 624.600 856.050 625.050 ;
        RECT 883.950 624.600 886.050 625.050 ;
        RECT 919.950 624.600 922.050 625.050 ;
        RECT 709.950 623.400 922.050 624.600 ;
        RECT 658.950 622.950 661.050 623.400 ;
        RECT 676.950 622.950 679.050 623.400 ;
        RECT 709.950 622.950 712.050 623.400 ;
        RECT 847.950 622.950 850.050 623.400 ;
        RECT 853.950 622.950 856.050 623.400 ;
        RECT 883.950 622.950 886.050 623.400 ;
        RECT 919.950 622.950 922.050 623.400 ;
        RECT 721.950 621.600 724.050 622.050 ;
        RECT 644.400 620.400 724.050 621.600 ;
        RECT 478.950 619.950 481.050 620.400 ;
        RECT 544.950 619.950 547.050 620.400 ;
        RECT 640.950 619.950 643.050 620.400 ;
        RECT 721.950 619.950 724.050 620.400 ;
        RECT 748.950 621.600 751.050 622.050 ;
        RECT 757.950 621.600 760.050 622.050 ;
        RECT 748.950 620.400 760.050 621.600 ;
        RECT 748.950 619.950 751.050 620.400 ;
        RECT 757.950 619.950 760.050 620.400 ;
        RECT 763.950 621.600 766.050 622.050 ;
        RECT 790.950 621.600 793.050 622.050 ;
        RECT 763.950 620.400 793.050 621.600 ;
        RECT 763.950 619.950 766.050 620.400 ;
        RECT 790.950 619.950 793.050 620.400 ;
        RECT 802.950 621.600 805.050 622.050 ;
        RECT 844.950 621.600 847.050 622.050 ;
        RECT 910.950 621.600 913.050 622.050 ;
        RECT 973.950 621.600 976.050 622.050 ;
        RECT 1018.950 621.600 1021.050 622.050 ;
        RECT 802.950 620.400 847.050 621.600 ;
        RECT 802.950 619.950 805.050 620.400 ;
        RECT 844.950 619.950 847.050 620.400 ;
        RECT 887.400 620.400 945.600 621.600 ;
        RECT 118.950 618.600 121.050 619.050 ;
        RECT 136.950 618.600 139.050 619.050 ;
        RECT 142.950 618.600 145.050 619.050 ;
        RECT 118.950 617.400 145.050 618.600 ;
        RECT 118.950 616.950 121.050 617.400 ;
        RECT 136.950 616.950 139.050 617.400 ;
        RECT 142.950 616.950 145.050 617.400 ;
        RECT 238.950 618.600 241.050 619.050 ;
        RECT 250.950 618.600 253.050 619.050 ;
        RECT 262.950 618.600 265.050 619.050 ;
        RECT 238.950 617.400 265.050 618.600 ;
        RECT 238.950 616.950 241.050 617.400 ;
        RECT 250.950 616.950 253.050 617.400 ;
        RECT 262.950 616.950 265.050 617.400 ;
        RECT 460.950 618.600 463.050 619.050 ;
        RECT 529.950 618.600 532.050 619.050 ;
        RECT 460.950 617.400 532.050 618.600 ;
        RECT 460.950 616.950 463.050 617.400 ;
        RECT 529.950 616.950 532.050 617.400 ;
        RECT 586.950 618.600 589.050 619.050 ;
        RECT 613.950 618.600 616.050 619.050 ;
        RECT 586.950 617.400 616.050 618.600 ;
        RECT 586.950 616.950 589.050 617.400 ;
        RECT 613.950 616.950 616.050 617.400 ;
        RECT 646.950 618.600 649.050 619.050 ;
        RECT 712.950 618.600 715.050 619.050 ;
        RECT 646.950 617.400 715.050 618.600 ;
        RECT 646.950 616.950 649.050 617.400 ;
        RECT 712.950 616.950 715.050 617.400 ;
        RECT 766.950 618.600 769.050 619.050 ;
        RECT 775.950 618.600 778.050 619.050 ;
        RECT 766.950 617.400 778.050 618.600 ;
        RECT 766.950 616.950 769.050 617.400 ;
        RECT 775.950 616.950 778.050 617.400 ;
        RECT 802.950 618.600 805.050 618.900 ;
        RECT 856.950 618.600 859.050 619.050 ;
        RECT 802.950 617.400 859.050 618.600 ;
        RECT 802.950 616.800 805.050 617.400 ;
        RECT 856.950 616.950 859.050 617.400 ;
        RECT 862.950 618.600 865.050 619.050 ;
        RECT 887.400 618.600 888.600 620.400 ;
        RECT 910.950 619.950 913.050 620.400 ;
        RECT 862.950 617.400 888.600 618.600 ;
        RECT 901.950 618.600 904.050 619.050 ;
        RECT 931.950 618.600 934.050 619.050 ;
        RECT 901.950 617.400 934.050 618.600 ;
        RECT 944.400 618.600 945.600 620.400 ;
        RECT 973.950 620.400 1021.050 621.600 ;
        RECT 973.950 619.950 976.050 620.400 ;
        RECT 1018.950 619.950 1021.050 620.400 ;
        RECT 1036.950 621.600 1039.050 622.050 ;
        RECT 1042.950 621.600 1045.050 622.050 ;
        RECT 1036.950 620.400 1045.050 621.600 ;
        RECT 1036.950 619.950 1039.050 620.400 ;
        RECT 1042.950 619.950 1045.050 620.400 ;
        RECT 970.950 618.600 973.050 619.050 ;
        RECT 944.400 617.400 973.050 618.600 ;
        RECT 862.950 616.950 865.050 617.400 ;
        RECT 901.950 616.950 904.050 617.400 ;
        RECT 931.950 616.950 934.050 617.400 ;
        RECT 970.950 616.950 973.050 617.400 ;
        RECT 25.950 615.600 28.050 616.050 ;
        RECT 31.950 615.600 34.050 616.050 ;
        RECT 202.950 615.600 205.050 616.050 ;
        RECT 25.950 614.400 205.050 615.600 ;
        RECT 25.950 613.950 28.050 614.400 ;
        RECT 31.950 613.950 34.050 614.400 ;
        RECT 202.950 613.950 205.050 614.400 ;
        RECT 346.950 615.600 349.050 616.050 ;
        RECT 379.950 615.600 382.050 616.050 ;
        RECT 394.950 615.600 397.050 616.050 ;
        RECT 346.950 614.400 397.050 615.600 ;
        RECT 346.950 613.950 349.050 614.400 ;
        RECT 379.950 613.950 382.050 614.400 ;
        RECT 394.950 613.950 397.050 614.400 ;
        RECT 400.950 615.600 403.050 616.050 ;
        RECT 406.950 615.600 409.050 616.050 ;
        RECT 415.950 615.600 418.050 616.050 ;
        RECT 400.950 614.400 418.050 615.600 ;
        RECT 400.950 613.950 403.050 614.400 ;
        RECT 406.950 613.950 409.050 614.400 ;
        RECT 415.950 613.950 418.050 614.400 ;
        RECT 553.950 615.600 556.050 616.050 ;
        RECT 568.950 615.600 571.050 616.050 ;
        RECT 553.950 614.400 571.050 615.600 ;
        RECT 553.950 613.950 556.050 614.400 ;
        RECT 568.950 613.950 571.050 614.400 ;
        RECT 619.950 615.600 622.050 616.050 ;
        RECT 631.950 615.600 634.050 616.050 ;
        RECT 619.950 614.400 634.050 615.600 ;
        RECT 619.950 613.950 622.050 614.400 ;
        RECT 631.950 613.950 634.050 614.400 ;
        RECT 664.950 615.600 667.050 616.050 ;
        RECT 703.950 615.600 706.050 616.050 ;
        RECT 736.950 615.600 739.050 616.050 ;
        RECT 805.950 615.600 808.050 616.050 ;
        RECT 664.950 614.400 699.600 615.600 ;
        RECT 664.950 613.950 667.050 614.400 ;
        RECT 698.400 613.050 699.600 614.400 ;
        RECT 703.950 614.400 808.050 615.600 ;
        RECT 703.950 613.950 706.050 614.400 ;
        RECT 736.950 613.950 739.050 614.400 ;
        RECT 805.950 613.950 808.050 614.400 ;
        RECT 973.950 615.600 976.050 616.050 ;
        RECT 979.950 615.600 982.050 616.050 ;
        RECT 973.950 614.400 982.050 615.600 ;
        RECT 973.950 613.950 976.050 614.400 ;
        RECT 979.950 613.950 982.050 614.400 ;
        RECT 121.950 612.600 124.050 613.050 ;
        RECT 142.950 612.600 145.050 613.050 ;
        RECT 166.950 612.600 169.050 613.050 ;
        RECT 178.950 612.600 181.050 613.050 ;
        RECT 241.950 612.600 244.050 613.050 ;
        RECT 121.950 611.400 141.600 612.600 ;
        RECT 121.950 610.950 124.050 611.400 ;
        RECT 64.950 609.600 67.050 610.050 ;
        RECT 109.950 609.600 112.050 610.050 ;
        RECT 64.950 608.400 112.050 609.600 ;
        RECT 140.400 609.600 141.600 611.400 ;
        RECT 142.950 611.400 181.050 612.600 ;
        RECT 142.950 610.950 145.050 611.400 ;
        RECT 166.950 610.950 169.050 611.400 ;
        RECT 178.950 610.950 181.050 611.400 ;
        RECT 233.400 611.400 244.050 612.600 ;
        RECT 160.950 609.600 163.050 610.050 ;
        RECT 140.400 608.400 163.050 609.600 ;
        RECT 64.950 607.950 67.050 608.400 ;
        RECT 109.950 607.950 112.050 608.400 ;
        RECT 160.950 607.950 163.050 608.400 ;
        RECT 193.950 609.600 196.050 610.050 ;
        RECT 214.950 609.600 217.050 610.050 ;
        RECT 193.950 608.400 217.050 609.600 ;
        RECT 193.950 607.950 196.050 608.400 ;
        RECT 214.950 607.950 217.050 608.400 ;
        RECT 37.800 606.000 39.900 607.050 ;
        RECT 40.950 606.600 43.050 607.050 ;
        RECT 157.950 606.750 160.050 607.200 ;
        RECT 163.950 606.750 166.050 607.200 ;
        RECT 37.800 604.950 40.050 606.000 ;
        RECT 40.950 605.400 63.600 606.600 ;
        RECT 40.950 604.950 43.050 605.400 ;
        RECT 37.950 603.600 40.050 604.950 ;
        RECT 58.950 603.600 61.050 604.050 ;
        RECT 37.950 603.000 61.050 603.600 ;
        RECT 38.250 602.400 61.050 603.000 ;
        RECT 58.950 601.950 61.050 602.400 ;
        RECT 34.950 600.600 37.050 601.050 ;
        RECT 43.950 600.600 46.050 600.900 ;
        RECT 34.950 599.400 46.050 600.600 ;
        RECT 34.950 598.950 37.050 599.400 ;
        RECT 43.950 598.800 46.050 599.400 ;
        RECT 62.400 597.600 63.600 605.400 ;
        RECT 157.950 605.550 166.050 606.750 ;
        RECT 157.950 605.100 160.050 605.550 ;
        RECT 163.950 605.100 166.050 605.550 ;
        RECT 220.950 606.750 223.050 607.200 ;
        RECT 226.950 606.750 229.050 607.200 ;
        RECT 233.400 607.050 234.600 611.400 ;
        RECT 241.950 610.950 244.050 611.400 ;
        RECT 283.950 612.600 286.050 613.050 ;
        RECT 298.950 612.600 301.050 613.050 ;
        RECT 283.950 611.400 301.050 612.600 ;
        RECT 283.950 610.950 286.050 611.400 ;
        RECT 298.950 610.950 301.050 611.400 ;
        RECT 382.950 612.600 385.050 613.050 ;
        RECT 397.950 612.600 400.050 613.050 ;
        RECT 382.950 611.400 400.050 612.600 ;
        RECT 382.950 610.950 385.050 611.400 ;
        RECT 397.950 610.950 400.050 611.400 ;
        RECT 445.950 612.600 448.050 613.050 ;
        RECT 493.950 612.600 496.050 613.050 ;
        RECT 445.950 611.400 496.050 612.600 ;
        RECT 445.950 610.950 448.050 611.400 ;
        RECT 493.950 610.950 496.050 611.400 ;
        RECT 244.950 607.950 247.050 610.050 ;
        RECT 376.950 609.600 379.050 610.050 ;
        RECT 400.950 609.600 403.050 610.050 ;
        RECT 376.950 608.400 403.050 609.600 ;
        RECT 376.950 607.950 379.050 608.400 ;
        RECT 400.950 607.950 403.050 608.400 ;
        RECT 409.950 609.600 412.050 610.050 ;
        RECT 418.950 609.600 421.050 610.050 ;
        RECT 409.950 608.400 421.050 609.600 ;
        RECT 409.950 607.950 412.050 608.400 ;
        RECT 418.950 607.950 421.050 608.400 ;
        RECT 436.950 609.600 439.050 610.050 ;
        RECT 469.950 609.600 472.050 610.050 ;
        RECT 436.950 608.400 472.050 609.600 ;
        RECT 436.950 607.950 439.050 608.400 ;
        RECT 469.950 607.950 472.050 608.400 ;
        RECT 499.950 609.600 502.050 610.050 ;
        RECT 505.800 609.600 507.900 610.050 ;
        RECT 499.950 608.400 507.900 609.600 ;
        RECT 499.950 607.950 502.050 608.400 ;
        RECT 505.800 607.950 507.900 608.400 ;
        RECT 508.950 609.600 511.050 610.050 ;
        RECT 538.950 609.600 541.050 610.050 ;
        RECT 508.950 608.400 541.050 609.600 ;
        RECT 541.950 609.600 544.050 613.050 ;
        RECT 565.950 612.600 568.050 613.050 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 565.950 611.400 598.050 612.600 ;
        RECT 565.950 610.950 568.050 611.400 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 697.950 612.600 700.050 613.050 ;
        RECT 751.950 612.600 754.050 613.050 ;
        RECT 769.950 612.600 772.050 613.050 ;
        RECT 697.950 611.400 735.600 612.600 ;
        RECT 697.950 610.950 700.050 611.400 ;
        RECT 580.950 609.600 583.050 610.050 ;
        RECT 619.950 609.600 622.050 610.050 ;
        RECT 541.950 609.000 622.050 609.600 ;
        RECT 542.400 608.400 622.050 609.000 ;
        RECT 508.950 607.950 511.050 608.400 ;
        RECT 538.950 607.950 541.050 608.400 ;
        RECT 580.950 607.950 583.050 608.400 ;
        RECT 619.950 607.950 622.050 608.400 ;
        RECT 640.950 609.600 643.050 610.050 ;
        RECT 652.950 609.600 655.050 610.050 ;
        RECT 640.950 608.400 655.050 609.600 ;
        RECT 640.950 607.950 643.050 608.400 ;
        RECT 652.950 607.950 655.050 608.400 ;
        RECT 667.950 609.600 670.050 610.050 ;
        RECT 685.950 609.600 688.050 610.050 ;
        RECT 724.950 609.600 727.050 610.050 ;
        RECT 667.950 608.400 727.050 609.600 ;
        RECT 734.400 609.600 735.600 611.400 ;
        RECT 751.950 611.400 772.050 612.600 ;
        RECT 751.950 610.950 754.050 611.400 ;
        RECT 769.950 610.950 772.050 611.400 ;
        RECT 787.950 612.600 790.050 613.050 ;
        RECT 826.950 612.600 829.050 613.050 ;
        RECT 787.950 611.400 829.050 612.600 ;
        RECT 787.950 610.950 790.050 611.400 ;
        RECT 826.950 610.950 829.050 611.400 ;
        RECT 835.950 612.600 838.050 613.050 ;
        RECT 841.950 612.600 844.050 613.050 ;
        RECT 835.950 611.400 844.050 612.600 ;
        RECT 835.950 610.950 838.050 611.400 ;
        RECT 841.950 610.950 844.050 611.400 ;
        RECT 859.950 612.600 862.050 613.050 ;
        RECT 868.950 612.600 871.050 613.050 ;
        RECT 859.950 611.400 871.050 612.600 ;
        RECT 859.950 610.950 862.050 611.400 ;
        RECT 868.950 610.950 871.050 611.400 ;
        RECT 946.950 612.600 949.050 613.050 ;
        RECT 958.950 612.600 961.050 613.050 ;
        RECT 946.950 611.400 961.050 612.600 ;
        RECT 946.950 610.950 949.050 611.400 ;
        RECT 958.950 610.950 961.050 611.400 ;
        RECT 964.950 612.600 967.050 613.050 ;
        RECT 982.950 612.600 985.050 613.050 ;
        RECT 964.950 611.400 985.050 612.600 ;
        RECT 964.950 610.950 967.050 611.400 ;
        RECT 982.950 610.950 985.050 611.400 ;
        RECT 1024.950 612.600 1027.050 613.050 ;
        RECT 1036.950 612.600 1039.050 613.050 ;
        RECT 1024.950 611.400 1039.050 612.600 ;
        RECT 1024.950 610.950 1027.050 611.400 ;
        RECT 1036.950 610.950 1039.050 611.400 ;
        RECT 781.950 609.600 784.050 610.050 ;
        RECT 734.400 608.400 784.050 609.600 ;
        RECT 667.950 607.950 670.050 608.400 ;
        RECT 685.950 607.950 688.050 608.400 ;
        RECT 724.950 607.950 727.050 608.400 ;
        RECT 781.950 607.950 784.050 608.400 ;
        RECT 790.950 609.600 793.050 610.050 ;
        RECT 832.950 609.600 835.050 610.050 ;
        RECT 790.950 608.400 835.050 609.600 ;
        RECT 790.950 607.950 793.050 608.400 ;
        RECT 832.950 607.950 835.050 608.400 ;
        RECT 850.950 609.600 853.050 610.050 ;
        RECT 913.950 609.600 916.050 610.050 ;
        RECT 850.950 608.400 882.600 609.600 ;
        RECT 850.950 607.950 853.050 608.400 ;
        RECT 220.950 605.550 229.050 606.750 ;
        RECT 220.950 605.100 223.050 605.550 ;
        RECT 226.950 605.100 229.050 605.550 ;
        RECT 232.950 604.950 235.050 607.050 ;
        RECT 79.950 603.750 82.050 604.200 ;
        RECT 100.950 603.750 103.050 604.200 ;
        RECT 79.950 602.550 103.050 603.750 ;
        RECT 79.950 602.100 82.050 602.550 ;
        RECT 100.950 602.100 103.050 602.550 ;
        RECT 106.950 603.450 109.050 603.900 ;
        RECT 127.950 603.450 130.050 603.900 ;
        RECT 106.950 602.250 130.050 603.450 ;
        RECT 106.950 601.800 109.050 602.250 ;
        RECT 127.950 601.800 130.050 602.250 ;
        RECT 139.950 600.600 142.050 600.900 ;
        RECT 154.950 600.600 157.050 601.050 ;
        RECT 139.950 599.400 157.050 600.600 ;
        RECT 139.950 598.800 142.050 599.400 ;
        RECT 154.950 598.950 157.050 599.400 ;
        RECT 202.950 600.600 205.050 601.050 ;
        RECT 245.400 600.900 246.600 607.950 ;
        RECT 268.950 606.600 271.050 607.050 ;
        RECT 280.950 606.750 283.050 607.200 ;
        RECT 289.950 606.750 292.050 607.200 ;
        RECT 280.950 606.600 292.050 606.750 ;
        RECT 268.950 605.550 292.050 606.600 ;
        RECT 268.950 605.400 283.050 605.550 ;
        RECT 268.950 604.950 271.050 605.400 ;
        RECT 280.950 605.100 283.050 605.400 ;
        RECT 289.950 605.100 292.050 605.550 ;
        RECT 295.950 606.600 298.050 607.200 ;
        RECT 304.950 606.600 307.050 607.050 ;
        RECT 295.950 605.400 307.050 606.600 ;
        RECT 295.950 605.100 298.050 605.400 ;
        RECT 304.950 604.950 307.050 605.400 ;
        RECT 361.950 606.750 364.050 607.200 ;
        RECT 367.950 606.750 370.050 607.200 ;
        RECT 361.950 605.550 370.050 606.750 ;
        RECT 361.950 605.100 364.050 605.550 ;
        RECT 367.950 605.100 370.050 605.550 ;
        RECT 448.950 606.750 451.050 607.200 ;
        RECT 454.950 606.750 457.050 607.200 ;
        RECT 448.950 605.550 457.050 606.750 ;
        RECT 562.950 606.600 565.050 607.050 ;
        RECT 448.950 605.100 451.050 605.550 ;
        RECT 454.950 605.100 457.050 605.550 ;
        RECT 518.400 605.400 565.050 606.600 ;
        RECT 211.950 600.600 214.050 600.900 ;
        RECT 202.950 599.400 214.050 600.600 ;
        RECT 202.950 598.950 205.050 599.400 ;
        RECT 211.950 598.800 214.050 599.400 ;
        RECT 232.950 600.450 235.050 600.900 ;
        RECT 238.950 600.450 241.050 600.900 ;
        RECT 232.950 599.250 241.050 600.450 ;
        RECT 232.950 598.800 235.050 599.250 ;
        RECT 238.950 598.800 241.050 599.250 ;
        RECT 244.950 598.800 247.050 600.900 ;
        RECT 256.950 600.450 259.050 600.900 ;
        RECT 265.950 600.450 268.050 600.900 ;
        RECT 256.950 599.250 268.050 600.450 ;
        RECT 256.950 598.800 259.050 599.250 ;
        RECT 265.950 598.800 268.050 599.250 ;
        RECT 310.950 600.450 313.050 600.900 ;
        RECT 322.950 600.450 325.050 600.900 ;
        RECT 310.950 599.250 325.050 600.450 ;
        RECT 310.950 598.800 313.050 599.250 ;
        RECT 322.950 598.800 325.050 599.250 ;
        RECT 349.950 600.450 352.050 600.900 ;
        RECT 358.950 600.450 361.050 600.900 ;
        RECT 349.950 599.250 361.050 600.450 ;
        RECT 349.950 598.800 352.050 599.250 ;
        RECT 358.950 598.800 361.050 599.250 ;
        RECT 373.950 600.450 376.050 600.900 ;
        RECT 379.950 600.450 382.050 600.900 ;
        RECT 373.950 599.250 382.050 600.450 ;
        RECT 373.950 598.800 376.050 599.250 ;
        RECT 379.950 598.800 382.050 599.250 ;
        RECT 421.950 600.450 424.050 600.900 ;
        RECT 433.950 600.450 436.050 600.900 ;
        RECT 421.950 599.250 436.050 600.450 ;
        RECT 421.950 598.800 424.050 599.250 ;
        RECT 433.950 598.800 436.050 599.250 ;
        RECT 439.950 600.450 442.050 600.900 ;
        RECT 445.950 600.450 448.050 600.900 ;
        RECT 439.950 599.250 448.050 600.450 ;
        RECT 439.950 598.800 442.050 599.250 ;
        RECT 445.950 598.800 448.050 599.250 ;
        RECT 460.950 600.600 463.050 601.050 ;
        RECT 518.400 600.900 519.600 605.400 ;
        RECT 562.950 604.950 565.050 605.400 ;
        RECT 601.950 606.600 604.050 607.200 ;
        RECT 664.950 606.600 667.050 607.200 ;
        RECT 601.950 605.400 667.050 606.600 ;
        RECT 601.950 605.100 604.050 605.400 ;
        RECT 664.950 605.100 667.050 605.400 ;
        RECT 670.950 606.600 673.050 607.200 ;
        RECT 730.950 606.600 733.050 607.200 ;
        RECT 742.950 606.600 745.050 607.050 ;
        RECT 670.950 605.400 681.600 606.600 ;
        RECT 670.950 605.100 673.050 605.400 ;
        RECT 607.950 603.600 610.050 604.050 ;
        RECT 655.950 603.600 658.050 604.050 ;
        RECT 607.950 602.400 658.050 603.600 ;
        RECT 607.950 601.950 610.050 602.400 ;
        RECT 655.950 601.950 658.050 602.400 ;
        RECT 680.400 601.050 681.600 605.400 ;
        RECT 730.950 605.400 745.050 606.600 ;
        RECT 730.950 605.100 733.050 605.400 ;
        RECT 742.950 604.950 745.050 605.400 ;
        RECT 748.950 606.600 751.050 607.050 ;
        RECT 766.950 606.600 769.050 607.050 ;
        RECT 748.950 605.400 769.050 606.600 ;
        RECT 748.950 604.950 751.050 605.400 ;
        RECT 766.950 604.950 769.050 605.400 ;
        RECT 799.950 606.750 802.050 607.200 ;
        RECT 814.950 606.750 817.050 607.200 ;
        RECT 799.950 605.550 817.050 606.750 ;
        RECT 799.950 605.100 802.050 605.550 ;
        RECT 814.950 605.100 817.050 605.550 ;
        RECT 823.950 606.600 826.050 607.050 ;
        RECT 829.950 606.600 832.050 607.050 ;
        RECT 823.950 605.400 832.050 606.600 ;
        RECT 833.400 606.600 834.600 607.950 ;
        RECT 835.950 606.600 838.050 607.200 ;
        RECT 833.400 605.400 838.050 606.600 ;
        RECT 823.950 604.950 826.050 605.400 ;
        RECT 829.950 604.950 832.050 605.400 ;
        RECT 835.950 605.100 838.050 605.400 ;
        RECT 856.950 605.100 859.050 607.200 ;
        RECT 862.950 605.100 865.050 607.200 ;
        RECT 881.400 606.600 882.600 608.400 ;
        RECT 908.400 608.400 916.050 609.600 ;
        RECT 892.950 606.600 895.050 607.050 ;
        RECT 881.400 605.400 895.050 606.600 ;
        RECT 820.950 603.600 823.050 604.050 ;
        RECT 788.400 602.400 823.050 603.600 ;
        RECT 469.950 600.600 472.050 600.900 ;
        RECT 460.950 599.400 472.050 600.600 ;
        RECT 460.950 598.950 463.050 599.400 ;
        RECT 469.950 598.800 472.050 599.400 ;
        RECT 484.950 600.450 487.050 600.900 ;
        RECT 496.950 600.450 499.050 600.900 ;
        RECT 484.950 599.250 499.050 600.450 ;
        RECT 484.950 598.800 487.050 599.250 ;
        RECT 496.950 598.800 499.050 599.250 ;
        RECT 517.950 598.800 520.050 600.900 ;
        RECT 523.950 600.450 526.050 600.900 ;
        RECT 529.950 600.450 532.050 600.900 ;
        RECT 523.950 599.250 532.050 600.450 ;
        RECT 523.950 598.800 526.050 599.250 ;
        RECT 529.950 598.800 532.050 599.250 ;
        RECT 613.950 600.600 616.050 601.050 ;
        RECT 622.950 600.600 625.050 600.900 ;
        RECT 613.950 599.400 625.050 600.600 ;
        RECT 613.950 598.950 616.050 599.400 ;
        RECT 622.950 598.800 625.050 599.400 ;
        RECT 640.950 600.450 643.050 600.900 ;
        RECT 652.950 600.450 655.050 601.050 ;
        RECT 640.950 599.250 655.050 600.450 ;
        RECT 640.950 598.800 643.050 599.250 ;
        RECT 652.950 598.950 655.050 599.250 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 788.400 600.900 789.600 602.400 ;
        RECT 820.950 601.950 823.050 602.400 ;
        RECT 826.950 603.600 831.000 604.050 ;
        RECT 826.950 601.950 831.600 603.600 ;
        RECT 688.950 600.450 691.050 600.900 ;
        RECT 694.950 600.450 697.050 600.900 ;
        RECT 688.950 599.250 697.050 600.450 ;
        RECT 688.950 598.800 691.050 599.250 ;
        RECT 694.950 598.800 697.050 599.250 ;
        RECT 721.950 600.450 724.050 600.900 ;
        RECT 727.950 600.450 730.050 600.900 ;
        RECT 721.950 599.250 730.050 600.450 ;
        RECT 721.950 598.800 724.050 599.250 ;
        RECT 727.950 598.800 730.050 599.250 ;
        RECT 751.950 600.450 754.050 600.900 ;
        RECT 760.950 600.450 763.050 600.900 ;
        RECT 751.950 599.250 763.050 600.450 ;
        RECT 751.950 598.800 754.050 599.250 ;
        RECT 760.950 598.800 763.050 599.250 ;
        RECT 787.950 598.800 790.050 600.900 ;
        RECT 799.950 600.600 802.050 601.050 ;
        RECT 817.950 600.600 820.050 601.050 ;
        RECT 799.950 599.400 820.050 600.600 ;
        RECT 830.400 600.600 831.600 601.950 ;
        RECT 853.950 600.600 856.050 601.050 ;
        RECT 830.400 599.400 856.050 600.600 ;
        RECT 857.400 600.600 858.600 605.100 ;
        RECT 863.400 603.600 864.600 605.100 ;
        RECT 892.950 604.950 895.050 605.400 ;
        RECT 863.400 602.400 867.600 603.600 ;
        RECT 866.400 600.600 867.600 602.400 ;
        RECT 880.950 600.600 883.050 600.900 ;
        RECT 857.400 600.000 864.600 600.600 ;
        RECT 857.400 599.400 865.050 600.000 ;
        RECT 866.400 599.400 883.050 600.600 ;
        RECT 799.950 598.950 802.050 599.400 ;
        RECT 817.950 598.950 820.050 599.400 ;
        RECT 853.950 598.950 856.050 599.400 ;
        RECT 64.950 597.600 67.050 598.050 ;
        RECT 115.950 597.600 118.050 598.050 ;
        RECT 62.400 596.400 118.050 597.600 ;
        RECT 64.950 595.950 67.050 596.400 ;
        RECT 115.950 595.950 118.050 596.400 ;
        RECT 190.950 597.600 193.050 598.050 ;
        RECT 199.950 597.600 202.050 598.050 ;
        RECT 190.950 596.400 202.050 597.600 ;
        RECT 190.950 595.950 193.050 596.400 ;
        RECT 199.950 595.950 202.050 596.400 ;
        RECT 292.950 597.600 295.050 598.050 ;
        RECT 316.950 597.600 319.050 598.050 ;
        RECT 292.950 596.400 319.050 597.600 ;
        RECT 359.400 597.600 360.600 598.800 ;
        RECT 598.950 597.600 601.050 598.050 ;
        RECT 359.400 596.400 601.050 597.600 ;
        RECT 292.950 595.950 295.050 596.400 ;
        RECT 316.950 595.950 319.050 596.400 ;
        RECT 598.950 595.950 601.050 596.400 ;
        RECT 673.950 597.600 676.050 598.050 ;
        RECT 706.950 597.600 709.050 598.050 ;
        RECT 718.950 597.600 721.050 598.050 ;
        RECT 733.950 597.600 736.050 598.050 ;
        RECT 673.950 596.400 684.600 597.600 ;
        RECT 673.950 595.950 676.050 596.400 ;
        RECT 28.950 594.600 31.050 595.050 ;
        RECT 52.950 594.600 55.050 595.050 ;
        RECT 28.950 593.400 55.050 594.600 ;
        RECT 28.950 592.950 31.050 593.400 ;
        RECT 52.950 592.950 55.050 593.400 ;
        RECT 181.950 594.600 184.050 595.050 ;
        RECT 220.950 594.600 223.050 595.050 ;
        RECT 181.950 593.400 223.050 594.600 ;
        RECT 181.950 592.950 184.050 593.400 ;
        RECT 220.950 592.950 223.050 593.400 ;
        RECT 469.950 594.600 472.050 595.050 ;
        RECT 493.950 594.600 496.050 595.050 ;
        RECT 568.950 594.600 571.050 595.050 ;
        RECT 469.950 593.400 571.050 594.600 ;
        RECT 469.950 592.950 472.050 593.400 ;
        RECT 493.950 592.950 496.050 593.400 ;
        RECT 568.950 592.950 571.050 593.400 ;
        RECT 667.950 594.600 670.050 595.050 ;
        RECT 676.950 594.600 679.050 595.050 ;
        RECT 667.950 593.400 679.050 594.600 ;
        RECT 683.400 594.600 684.600 596.400 ;
        RECT 706.950 596.400 736.050 597.600 ;
        RECT 706.950 595.950 709.050 596.400 ;
        RECT 718.950 595.950 721.050 596.400 ;
        RECT 733.950 595.950 736.050 596.400 ;
        RECT 835.950 597.600 838.050 598.050 ;
        RECT 841.950 597.600 844.050 598.050 ;
        RECT 835.950 596.400 844.050 597.600 ;
        RECT 835.950 595.950 838.050 596.400 ;
        RECT 841.950 595.950 844.050 596.400 ;
        RECT 862.950 595.950 865.050 599.400 ;
        RECT 880.950 598.800 883.050 599.400 ;
        RECT 886.950 600.600 889.050 600.900 ;
        RECT 901.950 600.600 904.050 601.050 ;
        RECT 908.400 600.900 909.600 608.400 ;
        RECT 913.950 607.950 916.050 608.400 ;
        RECT 973.950 609.600 976.050 610.050 ;
        RECT 1000.950 609.600 1003.050 610.050 ;
        RECT 1018.950 609.600 1021.050 610.050 ;
        RECT 973.950 608.400 981.600 609.600 ;
        RECT 973.950 607.950 976.050 608.400 ;
        RECT 916.950 606.600 919.050 607.200 ;
        RECT 925.950 606.600 928.050 607.050 ;
        RECT 934.950 606.600 937.050 607.200 ;
        RECT 955.950 606.600 958.050 607.050 ;
        RECT 916.950 605.400 928.050 606.600 ;
        RECT 916.950 605.100 919.050 605.400 ;
        RECT 886.950 599.400 904.050 600.600 ;
        RECT 886.950 598.800 889.050 599.400 ;
        RECT 901.950 598.950 904.050 599.400 ;
        RECT 907.950 598.800 910.050 600.900 ;
        RECT 917.400 600.600 918.600 605.100 ;
        RECT 925.950 604.950 928.050 605.400 ;
        RECT 932.400 605.400 937.050 606.600 ;
        RECT 925.950 603.600 928.050 603.900 ;
        RECT 932.400 603.600 933.600 605.400 ;
        RECT 934.950 605.100 937.050 605.400 ;
        RECT 947.400 605.400 958.050 606.600 ;
        RECT 925.950 602.400 933.600 603.600 ;
        RECT 925.950 601.800 928.050 602.400 ;
        RECT 947.400 601.050 948.600 605.400 ;
        RECT 955.950 604.950 958.050 605.400 ;
        RECT 964.950 604.950 967.050 607.050 ;
        RECT 965.400 601.050 966.600 604.950 ;
        RECT 931.950 600.600 934.050 601.050 ;
        RECT 917.400 599.400 934.050 600.600 ;
        RECT 931.950 598.950 934.050 599.400 ;
        RECT 943.950 599.400 948.600 601.050 ;
        RECT 952.950 600.600 955.050 601.050 ;
        RECT 958.950 600.600 961.050 600.900 ;
        RECT 952.950 599.400 961.050 600.600 ;
        RECT 943.950 598.950 948.000 599.400 ;
        RECT 952.950 598.950 955.050 599.400 ;
        RECT 958.950 598.800 961.050 599.400 ;
        RECT 964.950 598.950 967.050 601.050 ;
        RECT 980.400 600.900 981.600 608.400 ;
        RECT 1000.950 608.400 1021.050 609.600 ;
        RECT 1000.950 607.950 1003.050 608.400 ;
        RECT 1018.950 607.950 1021.050 608.400 ;
        RECT 982.950 606.600 985.050 607.200 ;
        RECT 988.950 606.600 991.050 607.050 ;
        RECT 982.950 605.400 991.050 606.600 ;
        RECT 982.950 605.100 985.050 605.400 ;
        RECT 988.950 604.950 991.050 605.400 ;
        RECT 1033.950 604.950 1036.050 607.050 ;
        RECT 1034.400 601.050 1035.600 604.950 ;
        RECT 979.950 598.800 982.050 600.900 ;
        RECT 997.950 600.450 1000.050 600.900 ;
        RECT 1003.950 600.450 1006.050 600.900 ;
        RECT 997.950 599.250 1006.050 600.450 ;
        RECT 997.950 598.800 1000.050 599.250 ;
        RECT 1003.950 598.800 1006.050 599.250 ;
        RECT 1018.950 600.600 1021.050 601.050 ;
        RECT 1024.950 600.600 1027.050 601.050 ;
        RECT 1018.950 599.400 1027.050 600.600 ;
        RECT 1018.950 598.950 1021.050 599.400 ;
        RECT 1024.950 598.950 1027.050 599.400 ;
        RECT 1033.950 598.950 1036.050 601.050 ;
        RECT 889.950 597.600 892.050 598.050 ;
        RECT 895.950 597.600 898.050 598.050 ;
        RECT 889.950 596.400 898.050 597.600 ;
        RECT 889.950 595.950 892.050 596.400 ;
        RECT 895.950 595.950 898.050 596.400 ;
        RECT 919.950 597.600 922.050 598.050 ;
        RECT 925.950 597.600 928.050 598.050 ;
        RECT 919.950 596.400 928.050 597.600 ;
        RECT 919.950 595.950 922.050 596.400 ;
        RECT 925.950 595.950 928.050 596.400 ;
        RECT 733.950 594.600 736.050 594.900 ;
        RECT 683.400 593.400 736.050 594.600 ;
        RECT 667.950 592.950 670.050 593.400 ;
        RECT 676.950 592.950 679.050 593.400 ;
        RECT 733.950 592.800 736.050 593.400 ;
        RECT 844.950 594.600 847.050 595.050 ;
        RECT 859.950 594.600 862.050 595.050 ;
        RECT 844.950 593.400 862.050 594.600 ;
        RECT 844.950 592.950 847.050 593.400 ;
        RECT 859.950 592.950 862.050 593.400 ;
        RECT 865.950 594.600 868.050 595.050 ;
        RECT 892.950 594.600 895.050 595.050 ;
        RECT 865.950 593.400 895.050 594.600 ;
        RECT 865.950 592.950 868.050 593.400 ;
        RECT 892.950 592.950 895.050 593.400 ;
        RECT 916.950 594.600 919.050 595.050 ;
        RECT 937.950 594.600 940.050 595.050 ;
        RECT 916.950 593.400 940.050 594.600 ;
        RECT 916.950 592.950 919.050 593.400 ;
        RECT 937.950 592.950 940.050 593.400 ;
        RECT 970.950 594.600 973.050 595.050 ;
        RECT 985.950 594.600 988.050 595.050 ;
        RECT 970.950 593.400 988.050 594.600 ;
        RECT 970.950 592.950 973.050 593.400 ;
        RECT 985.950 592.950 988.050 593.400 ;
        RECT 112.950 591.600 115.050 592.050 ;
        RECT 118.950 591.600 121.050 592.050 ;
        RECT 71.400 591.000 121.050 591.600 ;
        RECT 70.950 590.400 121.050 591.000 ;
        RECT 70.950 586.950 73.050 590.400 ;
        RECT 112.950 589.950 115.050 590.400 ;
        RECT 118.950 589.950 121.050 590.400 ;
        RECT 160.950 591.600 163.050 592.050 ;
        RECT 172.950 591.600 175.050 592.050 ;
        RECT 160.950 590.400 175.050 591.600 ;
        RECT 160.950 589.950 163.050 590.400 ;
        RECT 172.950 589.950 175.050 590.400 ;
        RECT 232.950 591.600 235.050 592.050 ;
        RECT 343.950 591.600 346.050 592.050 ;
        RECT 232.950 590.400 346.050 591.600 ;
        RECT 232.950 589.950 235.050 590.400 ;
        RECT 343.950 589.950 346.050 590.400 ;
        RECT 418.950 591.600 421.050 592.050 ;
        RECT 436.950 591.600 439.050 592.050 ;
        RECT 418.950 590.400 439.050 591.600 ;
        RECT 418.950 589.950 421.050 590.400 ;
        RECT 436.950 589.950 439.050 590.400 ;
        RECT 448.950 591.600 451.050 592.050 ;
        RECT 553.950 591.600 556.050 592.050 ;
        RECT 448.950 590.400 556.050 591.600 ;
        RECT 448.950 589.950 451.050 590.400 ;
        RECT 553.950 589.950 556.050 590.400 ;
        RECT 592.950 591.600 595.050 592.050 ;
        RECT 673.950 591.600 676.050 592.050 ;
        RECT 592.950 590.400 676.050 591.600 ;
        RECT 592.950 589.950 595.050 590.400 ;
        RECT 673.950 589.950 676.050 590.400 ;
        RECT 679.950 591.600 682.050 592.050 ;
        RECT 718.800 591.600 720.900 592.050 ;
        RECT 679.950 590.400 720.900 591.600 ;
        RECT 679.950 589.950 682.050 590.400 ;
        RECT 718.800 589.950 720.900 590.400 ;
        RECT 721.950 591.600 724.050 592.050 ;
        RECT 772.950 591.600 775.050 591.900 ;
        RECT 796.950 591.600 799.050 592.050 ;
        RECT 721.950 590.400 735.600 591.600 ;
        RECT 721.950 589.950 724.050 590.400 ;
        RECT 79.950 588.600 82.050 589.050 ;
        RECT 100.950 588.600 103.050 589.050 ;
        RECT 79.950 587.400 103.050 588.600 ;
        RECT 79.950 586.950 82.050 587.400 ;
        RECT 100.950 586.950 103.050 587.400 ;
        RECT 127.950 588.600 130.050 589.050 ;
        RECT 205.950 588.600 208.050 589.050 ;
        RECT 127.950 587.400 208.050 588.600 ;
        RECT 127.950 586.950 130.050 587.400 ;
        RECT 205.950 586.950 208.050 587.400 ;
        RECT 505.950 588.600 508.050 589.050 ;
        RECT 601.950 588.600 604.050 589.050 ;
        RECT 637.950 588.600 640.050 589.050 ;
        RECT 505.950 587.400 582.600 588.600 ;
        RECT 505.950 586.950 508.050 587.400 ;
        RECT 166.950 585.600 169.050 586.050 ;
        RECT 178.950 585.600 181.050 586.050 ;
        RECT 166.950 584.400 181.050 585.600 ;
        RECT 166.950 583.950 169.050 584.400 ;
        RECT 178.950 583.950 181.050 584.400 ;
        RECT 271.950 585.600 274.050 586.050 ;
        RECT 361.950 585.600 364.050 586.050 ;
        RECT 271.950 584.400 364.050 585.600 ;
        RECT 271.950 583.950 274.050 584.400 ;
        RECT 361.950 583.950 364.050 584.400 ;
        RECT 427.950 585.600 430.050 586.050 ;
        RECT 574.950 585.600 577.050 586.050 ;
        RECT 427.950 584.400 577.050 585.600 ;
        RECT 581.400 585.600 582.600 587.400 ;
        RECT 601.950 587.400 640.050 588.600 ;
        RECT 601.950 586.950 604.050 587.400 ;
        RECT 637.950 586.950 640.050 587.400 ;
        RECT 655.950 588.600 658.050 589.050 ;
        RECT 712.950 588.600 715.050 589.050 ;
        RECT 655.950 587.400 715.050 588.600 ;
        RECT 734.400 588.600 735.600 590.400 ;
        RECT 772.950 590.400 799.050 591.600 ;
        RECT 772.950 589.800 775.050 590.400 ;
        RECT 796.950 589.950 799.050 590.400 ;
        RECT 940.950 591.600 943.050 592.050 ;
        RECT 958.950 591.600 961.050 592.050 ;
        RECT 940.950 590.400 961.050 591.600 ;
        RECT 940.950 589.950 943.050 590.400 ;
        RECT 958.950 589.950 961.050 590.400 ;
        RECT 976.950 591.600 979.050 592.050 ;
        RECT 982.950 591.600 985.050 592.050 ;
        RECT 976.950 590.400 985.050 591.600 ;
        RECT 976.950 589.950 979.050 590.400 ;
        RECT 982.950 589.950 985.050 590.400 ;
        RECT 997.950 591.600 1000.050 592.050 ;
        RECT 1033.950 591.600 1036.050 592.050 ;
        RECT 997.950 590.400 1036.050 591.600 ;
        RECT 997.950 589.950 1000.050 590.400 ;
        RECT 1033.950 589.950 1036.050 590.400 ;
        RECT 748.950 588.600 751.050 589.050 ;
        RECT 734.400 587.400 751.050 588.600 ;
        RECT 655.950 586.950 658.050 587.400 ;
        RECT 712.950 586.950 715.050 587.400 ;
        RECT 748.950 586.950 751.050 587.400 ;
        RECT 769.950 588.600 772.050 589.050 ;
        RECT 787.950 588.600 790.050 589.050 ;
        RECT 769.950 587.400 790.050 588.600 ;
        RECT 769.950 586.950 772.050 587.400 ;
        RECT 787.950 586.950 790.050 587.400 ;
        RECT 829.950 588.600 832.050 589.050 ;
        RECT 850.950 588.600 853.050 589.050 ;
        RECT 829.950 587.400 853.050 588.600 ;
        RECT 829.950 586.950 832.050 587.400 ;
        RECT 850.950 586.950 853.050 587.400 ;
        RECT 898.950 588.600 901.050 589.050 ;
        RECT 919.950 588.600 922.050 589.050 ;
        RECT 898.950 587.400 922.050 588.600 ;
        RECT 898.950 586.950 901.050 587.400 ;
        RECT 919.950 586.950 922.050 587.400 ;
        RECT 925.950 588.600 928.050 589.050 ;
        RECT 937.950 588.600 940.050 589.050 ;
        RECT 925.950 587.400 940.050 588.600 ;
        RECT 925.950 586.950 928.050 587.400 ;
        RECT 937.950 586.950 940.050 587.400 ;
        RECT 673.950 585.600 676.050 586.050 ;
        RECT 775.950 585.600 778.050 586.050 ;
        RECT 799.950 585.600 802.050 586.050 ;
        RECT 826.950 585.600 829.050 586.050 ;
        RECT 581.400 584.400 829.050 585.600 ;
        RECT 427.950 583.950 430.050 584.400 ;
        RECT 574.950 583.950 577.050 584.400 ;
        RECT 673.950 583.950 676.050 584.400 ;
        RECT 775.950 583.950 778.050 584.400 ;
        RECT 799.950 583.950 802.050 584.400 ;
        RECT 826.950 583.950 829.050 584.400 ;
        RECT 832.950 585.600 835.050 586.050 ;
        RECT 856.950 585.600 859.050 586.050 ;
        RECT 832.950 584.400 859.050 585.600 ;
        RECT 832.950 583.950 835.050 584.400 ;
        RECT 856.950 583.950 859.050 584.400 ;
        RECT 871.950 585.600 874.050 586.050 ;
        RECT 895.950 585.600 898.050 586.050 ;
        RECT 871.950 584.400 898.050 585.600 ;
        RECT 871.950 583.950 874.050 584.400 ;
        RECT 895.950 583.950 898.050 584.400 ;
        RECT 955.950 585.600 958.050 586.050 ;
        RECT 976.950 585.600 979.050 586.050 ;
        RECT 955.950 584.400 979.050 585.600 ;
        RECT 955.950 583.950 958.050 584.400 ;
        RECT 976.950 583.950 979.050 584.400 ;
        RECT 1012.950 585.600 1015.050 586.050 ;
        RECT 1042.950 585.600 1045.050 586.050 ;
        RECT 1012.950 584.400 1045.050 585.600 ;
        RECT 1012.950 583.950 1015.050 584.400 ;
        RECT 1042.950 583.950 1045.050 584.400 ;
        RECT 58.950 582.600 61.050 583.050 ;
        RECT 91.950 582.600 94.050 583.050 ;
        RECT 58.950 581.400 94.050 582.600 ;
        RECT 58.950 580.950 61.050 581.400 ;
        RECT 91.950 580.950 94.050 581.400 ;
        RECT 145.950 582.600 148.050 583.050 ;
        RECT 157.950 582.600 160.050 583.050 ;
        RECT 223.950 582.600 226.050 583.050 ;
        RECT 145.950 581.400 162.600 582.600 ;
        RECT 145.950 580.950 148.050 581.400 ;
        RECT 157.950 580.950 160.050 581.400 ;
        RECT 161.400 579.600 162.600 581.400 ;
        RECT 182.400 581.400 226.050 582.600 ;
        RECT 182.400 579.600 183.600 581.400 ;
        RECT 223.950 580.950 226.050 581.400 ;
        RECT 244.950 582.600 247.050 583.050 ;
        RECT 331.950 582.600 334.050 583.050 ;
        RECT 244.950 581.400 334.050 582.600 ;
        RECT 244.950 580.950 247.050 581.400 ;
        RECT 331.950 580.950 334.050 581.400 ;
        RECT 397.950 582.600 400.050 583.050 ;
        RECT 454.950 582.600 457.050 583.050 ;
        RECT 514.950 582.600 517.050 583.050 ;
        RECT 397.950 581.400 517.050 582.600 ;
        RECT 397.950 580.950 400.050 581.400 ;
        RECT 454.950 580.950 457.050 581.400 ;
        RECT 514.950 580.950 517.050 581.400 ;
        RECT 577.950 582.600 580.050 583.050 ;
        RECT 586.950 582.600 589.050 583.050 ;
        RECT 607.950 582.600 610.050 583.050 ;
        RECT 634.950 582.600 637.050 583.050 ;
        RECT 688.950 582.600 691.050 583.050 ;
        RECT 727.950 582.600 730.050 583.050 ;
        RECT 760.950 582.600 763.050 583.050 ;
        RECT 577.950 581.400 660.600 582.600 ;
        RECT 577.950 580.950 580.050 581.400 ;
        RECT 586.950 580.950 589.050 581.400 ;
        RECT 607.950 580.950 610.050 581.400 ;
        RECT 634.950 580.950 637.050 581.400 ;
        RECT 161.400 578.400 183.600 579.600 ;
        RECT 367.950 579.600 370.050 580.050 ;
        RECT 400.950 579.600 403.050 580.050 ;
        RECT 367.950 578.400 403.050 579.600 ;
        RECT 367.950 577.950 370.050 578.400 ;
        RECT 400.950 577.950 403.050 578.400 ;
        RECT 421.950 579.600 424.050 580.050 ;
        RECT 532.950 579.600 535.050 580.050 ;
        RECT 544.950 579.600 547.050 580.050 ;
        RECT 421.950 578.400 441.600 579.600 ;
        RECT 421.950 577.950 424.050 578.400 ;
        RECT 49.950 576.600 52.050 577.050 ;
        RECT 58.950 576.600 61.050 577.050 ;
        RECT 49.950 575.400 61.050 576.600 ;
        RECT 49.950 574.950 52.050 575.400 ;
        RECT 58.950 574.950 61.050 575.400 ;
        RECT 136.950 576.600 139.050 577.050 ;
        RECT 148.950 576.600 151.050 577.050 ;
        RECT 136.950 575.400 151.050 576.600 ;
        RECT 136.950 574.950 139.050 575.400 ;
        RECT 148.950 574.950 151.050 575.400 ;
        RECT 271.950 576.600 274.050 577.050 ;
        RECT 277.950 576.600 280.050 577.050 ;
        RECT 271.950 575.400 280.050 576.600 ;
        RECT 440.400 576.600 441.600 578.400 ;
        RECT 532.950 578.400 547.050 579.600 ;
        RECT 659.400 579.600 660.600 581.400 ;
        RECT 688.950 581.400 723.600 582.600 ;
        RECT 688.950 580.950 691.050 581.400 ;
        RECT 667.950 579.600 670.050 580.050 ;
        RECT 659.400 578.400 670.050 579.600 ;
        RECT 722.400 579.600 723.600 581.400 ;
        RECT 727.950 581.400 763.050 582.600 ;
        RECT 727.950 580.950 730.050 581.400 ;
        RECT 760.950 580.950 763.050 581.400 ;
        RECT 841.950 582.600 844.050 583.050 ;
        RECT 868.950 582.600 871.050 583.050 ;
        RECT 916.950 582.600 919.050 583.050 ;
        RECT 841.950 581.400 871.050 582.600 ;
        RECT 841.950 580.950 844.050 581.400 ;
        RECT 868.950 580.950 871.050 581.400 ;
        RECT 896.400 581.400 919.050 582.600 ;
        RECT 754.950 579.600 757.050 580.050 ;
        RECT 722.400 578.400 757.050 579.600 ;
        RECT 532.950 577.950 535.050 578.400 ;
        RECT 544.950 577.950 547.050 578.400 ;
        RECT 667.950 577.950 670.050 578.400 ;
        RECT 754.950 577.950 757.050 578.400 ;
        RECT 811.950 579.600 814.050 580.050 ;
        RECT 820.950 579.600 823.050 580.050 ;
        RECT 811.950 578.400 823.050 579.600 ;
        RECT 811.950 577.950 814.050 578.400 ;
        RECT 820.950 577.950 823.050 578.400 ;
        RECT 865.950 579.600 868.050 580.050 ;
        RECT 896.400 579.600 897.600 581.400 ;
        RECT 916.950 580.950 919.050 581.400 ;
        RECT 925.950 582.600 928.050 583.050 ;
        RECT 934.950 582.600 937.050 583.050 ;
        RECT 925.950 581.400 937.050 582.600 ;
        RECT 925.950 580.950 928.050 581.400 ;
        RECT 934.950 580.950 937.050 581.400 ;
        RECT 940.950 582.600 943.050 583.050 ;
        RECT 952.950 582.600 955.050 583.050 ;
        RECT 940.950 581.400 955.050 582.600 ;
        RECT 940.950 580.950 943.050 581.400 ;
        RECT 952.950 580.950 955.050 581.400 ;
        RECT 994.950 582.600 997.050 583.050 ;
        RECT 1000.950 582.600 1003.050 583.050 ;
        RECT 994.950 581.400 1003.050 582.600 ;
        RECT 994.950 580.950 997.050 581.400 ;
        RECT 1000.950 580.950 1003.050 581.400 ;
        RECT 1009.950 582.600 1012.050 583.050 ;
        RECT 1039.950 582.600 1042.050 583.050 ;
        RECT 1009.950 581.400 1042.050 582.600 ;
        RECT 1009.950 580.950 1012.050 581.400 ;
        RECT 1039.950 580.950 1042.050 581.400 ;
        RECT 865.950 578.400 897.600 579.600 ;
        RECT 898.950 579.600 901.050 580.050 ;
        RECT 907.950 579.600 910.050 580.050 ;
        RECT 898.950 578.400 910.050 579.600 ;
        RECT 865.950 577.950 868.050 578.400 ;
        RECT 898.950 577.950 901.050 578.400 ;
        RECT 907.950 577.950 910.050 578.400 ;
        RECT 964.950 579.600 967.050 580.050 ;
        RECT 979.950 579.600 982.050 580.050 ;
        RECT 964.950 578.400 982.050 579.600 ;
        RECT 964.950 577.950 967.050 578.400 ;
        RECT 979.950 577.950 982.050 578.400 ;
        RECT 985.950 579.600 988.050 580.050 ;
        RECT 994.950 579.600 997.050 579.900 ;
        RECT 1036.950 579.600 1039.050 580.050 ;
        RECT 985.950 578.400 997.050 579.600 ;
        RECT 985.950 577.950 988.050 578.400 ;
        RECT 994.950 577.800 997.050 578.400 ;
        RECT 1031.400 578.400 1039.050 579.600 ;
        RECT 454.950 576.600 457.050 577.050 ;
        RECT 440.400 575.400 457.050 576.600 ;
        RECT 271.950 574.950 274.050 575.400 ;
        RECT 277.950 574.950 280.050 575.400 ;
        RECT 454.950 574.950 457.050 575.400 ;
        RECT 487.950 576.600 490.050 577.050 ;
        RECT 502.950 576.600 505.050 577.050 ;
        RECT 487.950 575.400 505.050 576.600 ;
        RECT 487.950 574.950 490.050 575.400 ;
        RECT 502.950 574.950 505.050 575.400 ;
        RECT 511.950 576.600 514.050 577.050 ;
        RECT 523.950 576.600 526.050 577.050 ;
        RECT 511.950 575.400 526.050 576.600 ;
        RECT 511.950 574.950 514.050 575.400 ;
        RECT 523.950 574.950 526.050 575.400 ;
        RECT 610.950 576.600 613.050 577.050 ;
        RECT 679.950 576.600 682.050 577.050 ;
        RECT 610.950 575.400 682.050 576.600 ;
        RECT 610.950 574.950 613.050 575.400 ;
        RECT 679.950 574.950 682.050 575.400 ;
        RECT 694.950 576.600 697.050 577.050 ;
        RECT 712.950 576.600 715.050 577.050 ;
        RECT 694.950 575.400 715.050 576.600 ;
        RECT 694.950 574.950 697.050 575.400 ;
        RECT 712.950 574.950 715.050 575.400 ;
        RECT 718.950 576.600 721.050 577.050 ;
        RECT 772.950 576.600 775.050 577.050 ;
        RECT 816.000 576.600 820.050 577.050 ;
        RECT 718.950 575.400 775.050 576.600 ;
        RECT 718.950 574.950 721.050 575.400 ;
        RECT 772.950 574.950 775.050 575.400 ;
        RECT 815.400 574.950 820.050 576.600 ;
        RECT 871.950 576.600 874.050 577.050 ;
        RECT 886.950 576.600 889.050 577.050 ;
        RECT 871.950 575.400 889.050 576.600 ;
        RECT 871.950 574.950 874.050 575.400 ;
        RECT 886.950 574.950 889.050 575.400 ;
        RECT 913.950 576.600 916.050 577.050 ;
        RECT 931.950 576.600 934.050 577.050 ;
        RECT 913.950 575.400 934.050 576.600 ;
        RECT 913.950 574.950 916.050 575.400 ;
        RECT 19.950 573.600 22.050 574.200 ;
        RECT 37.950 573.750 40.050 574.200 ;
        RECT 46.950 573.750 49.050 574.200 ;
        RECT 37.950 573.600 49.050 573.750 ;
        RECT 19.950 572.550 49.050 573.600 ;
        RECT 19.950 572.400 40.050 572.550 ;
        RECT 19.950 572.100 22.050 572.400 ;
        RECT 37.950 572.100 40.050 572.400 ;
        RECT 46.950 572.100 49.050 572.550 ;
        RECT 97.950 573.750 100.050 574.200 ;
        RECT 106.950 573.750 109.050 574.200 ;
        RECT 97.950 572.550 109.050 573.750 ;
        RECT 97.950 572.100 100.050 572.550 ;
        RECT 106.950 572.100 109.050 572.550 ;
        RECT 118.950 572.100 121.050 574.200 ;
        RECT 160.950 573.600 163.050 574.200 ;
        RECT 208.950 573.600 211.050 574.050 ;
        RECT 235.950 573.600 238.050 574.200 ;
        RECT 160.950 572.400 180.600 573.600 ;
        RECT 160.950 572.100 163.050 572.400 ;
        RECT 119.400 568.050 120.600 572.100 ;
        RECT 179.400 570.900 180.600 572.400 ;
        RECT 208.950 572.400 238.050 573.600 ;
        RECT 208.950 571.950 211.050 572.400 ;
        RECT 235.950 572.100 238.050 572.400 ;
        RECT 280.950 573.750 283.050 574.200 ;
        RECT 292.950 573.750 295.050 574.200 ;
        RECT 280.950 572.550 295.050 573.750 ;
        RECT 280.950 572.100 283.050 572.550 ;
        RECT 292.950 572.100 295.050 572.550 ;
        RECT 340.950 573.600 343.050 574.200 ;
        RECT 352.800 573.600 354.900 574.050 ;
        RECT 340.950 572.400 354.900 573.600 ;
        RECT 340.950 572.100 343.050 572.400 ;
        RECT 352.800 571.950 354.900 572.400 ;
        RECT 355.950 573.750 358.050 574.200 ;
        RECT 373.950 573.750 376.050 574.200 ;
        RECT 355.950 572.550 376.050 573.750 ;
        RECT 355.950 572.100 358.050 572.550 ;
        RECT 373.950 572.100 376.050 572.550 ;
        RECT 391.950 573.600 394.050 573.900 ;
        RECT 406.950 573.600 409.050 574.050 ;
        RECT 430.950 573.600 433.050 574.200 ;
        RECT 391.950 572.400 409.050 573.600 ;
        RECT 391.950 571.800 394.050 572.400 ;
        RECT 406.950 571.950 409.050 572.400 ;
        RECT 410.400 572.400 433.050 573.600 ;
        RECT 178.950 568.800 181.050 570.900 ;
        RECT 199.950 570.600 202.050 571.050 ;
        RECT 325.950 570.600 328.050 571.050 ;
        RECT 410.400 570.600 411.600 572.400 ;
        RECT 430.950 572.100 433.050 572.400 ;
        RECT 436.950 573.750 439.050 574.200 ;
        RECT 442.950 573.750 445.050 574.200 ;
        RECT 436.950 572.550 445.050 573.750 ;
        RECT 436.950 572.100 439.050 572.550 ;
        RECT 442.950 572.100 445.050 572.550 ;
        RECT 460.950 573.600 463.050 574.200 ;
        RECT 484.950 573.600 487.050 574.200 ;
        RECT 460.950 572.400 487.050 573.600 ;
        RECT 460.950 572.100 463.050 572.400 ;
        RECT 484.950 572.100 487.050 572.400 ;
        RECT 508.950 573.600 511.050 574.050 ;
        RECT 520.950 573.600 523.050 574.050 ;
        RECT 508.950 572.400 523.050 573.600 ;
        RECT 508.950 571.950 511.050 572.400 ;
        RECT 520.950 571.950 523.050 572.400 ;
        RECT 538.950 573.600 541.050 574.200 ;
        RECT 550.950 573.600 553.050 574.050 ;
        RECT 559.950 573.600 562.050 574.200 ;
        RECT 538.950 572.400 562.050 573.600 ;
        RECT 538.950 572.100 541.050 572.400 ;
        RECT 550.950 571.950 553.050 572.400 ;
        RECT 559.950 572.100 562.050 572.400 ;
        RECT 565.950 572.100 568.050 574.200 ;
        RECT 613.950 573.600 616.050 574.200 ;
        RECT 643.950 573.750 646.050 574.200 ;
        RECT 655.950 573.750 658.050 574.200 ;
        RECT 613.950 572.400 642.600 573.600 ;
        RECT 613.950 572.100 616.050 572.400 ;
        RECT 199.950 569.400 225.600 570.600 ;
        RECT 199.950 568.950 202.050 569.400 ;
        RECT 22.950 567.450 25.050 567.900 ;
        RECT 28.950 567.600 31.050 567.900 ;
        RECT 43.950 567.600 46.050 567.900 ;
        RECT 28.950 567.450 46.050 567.600 ;
        RECT 22.950 566.400 46.050 567.450 ;
        RECT 22.950 566.250 31.050 566.400 ;
        RECT 22.950 565.800 25.050 566.250 ;
        RECT 28.950 565.800 31.050 566.250 ;
        RECT 43.950 565.800 46.050 566.400 ;
        RECT 49.950 567.600 52.050 567.900 ;
        RECT 49.950 566.400 90.600 567.600 ;
        RECT 49.950 565.800 52.050 566.400 ;
        RECT 37.950 564.600 40.050 565.050 ;
        RECT 49.950 564.600 52.050 564.750 ;
        RECT 37.950 563.400 52.050 564.600 ;
        RECT 89.400 564.600 90.600 566.400 ;
        RECT 115.950 566.400 120.600 568.050 ;
        RECT 127.950 567.600 130.050 568.050 ;
        RECT 145.950 567.600 148.050 567.900 ;
        RECT 127.950 566.400 148.050 567.600 ;
        RECT 224.400 567.600 225.600 569.400 ;
        RECT 325.950 569.400 411.600 570.600 ;
        RECT 475.950 570.600 478.050 571.050 ;
        RECT 499.950 570.600 502.050 571.050 ;
        RECT 475.950 569.400 502.050 570.600 ;
        RECT 325.950 568.950 328.050 569.400 ;
        RECT 475.950 568.950 478.050 569.400 ;
        RECT 499.950 568.950 502.050 569.400 ;
        RECT 526.950 570.600 529.050 571.050 ;
        RECT 566.400 570.600 567.600 572.100 ;
        RECT 526.950 569.400 567.600 570.600 ;
        RECT 526.950 568.950 529.050 569.400 ;
        RECT 232.950 567.600 235.050 568.050 ;
        RECT 224.400 566.400 235.050 567.600 ;
        RECT 115.950 565.950 120.000 566.400 ;
        RECT 127.950 565.950 130.050 566.400 ;
        RECT 145.950 565.800 148.050 566.400 ;
        RECT 232.950 565.950 235.050 566.400 ;
        RECT 250.950 567.450 253.050 567.900 ;
        RECT 262.950 567.450 265.050 567.900 ;
        RECT 250.950 566.250 265.050 567.450 ;
        RECT 250.950 565.800 253.050 566.250 ;
        RECT 262.950 565.800 265.050 566.250 ;
        RECT 268.950 567.600 271.050 567.900 ;
        RECT 289.950 567.600 292.050 567.900 ;
        RECT 307.950 567.600 310.050 568.050 ;
        RECT 268.950 566.400 310.050 567.600 ;
        RECT 268.950 565.800 271.050 566.400 ;
        RECT 289.950 565.800 292.050 566.400 ;
        RECT 307.950 565.950 310.050 566.400 ;
        RECT 331.950 567.450 334.050 567.900 ;
        RECT 343.950 567.450 346.050 567.900 ;
        RECT 331.950 566.250 346.050 567.450 ;
        RECT 331.950 565.800 334.050 566.250 ;
        RECT 343.950 565.800 346.050 566.250 ;
        RECT 352.950 567.450 355.050 567.900 ;
        RECT 370.950 567.450 373.050 567.900 ;
        RECT 352.950 566.250 373.050 567.450 ;
        RECT 352.950 565.800 355.050 566.250 ;
        RECT 370.950 565.800 373.050 566.250 ;
        RECT 433.950 567.600 436.050 567.900 ;
        RECT 433.950 566.400 438.600 567.600 ;
        RECT 433.950 565.800 436.050 566.400 ;
        RECT 94.950 564.600 97.050 565.050 ;
        RECT 89.400 563.400 97.050 564.600 ;
        RECT 37.950 562.950 40.050 563.400 ;
        RECT 49.950 562.650 52.050 563.400 ;
        RECT 94.950 562.950 97.050 563.400 ;
        RECT 109.950 564.450 112.050 564.900 ;
        RECT 154.950 564.450 157.050 564.900 ;
        RECT 109.950 563.250 157.050 564.450 ;
        RECT 437.400 564.600 438.600 566.400 ;
        RECT 463.950 567.450 466.050 567.900 ;
        RECT 469.950 567.450 472.050 567.900 ;
        RECT 463.950 566.250 472.050 567.450 ;
        RECT 463.950 565.800 466.050 566.250 ;
        RECT 469.950 565.800 472.050 566.250 ;
        RECT 511.950 567.600 514.050 567.900 ;
        RECT 523.950 567.600 526.050 568.050 ;
        RECT 511.950 566.400 526.050 567.600 ;
        RECT 511.950 565.800 514.050 566.400 ;
        RECT 523.950 565.950 526.050 566.400 ;
        RECT 544.950 567.600 547.050 568.050 ;
        RECT 641.400 567.900 642.600 572.400 ;
        RECT 643.950 572.550 658.050 573.750 ;
        RECT 643.950 572.100 646.050 572.550 ;
        RECT 655.950 572.100 658.050 572.550 ;
        RECT 691.950 573.600 696.000 574.050 ;
        RECT 697.950 573.600 700.050 574.200 ;
        RECT 709.950 573.600 712.050 574.050 ;
        RECT 691.950 571.950 696.600 573.600 ;
        RECT 697.950 572.400 712.050 573.600 ;
        RECT 697.950 572.100 700.050 572.400 ;
        RECT 709.950 571.950 712.050 572.400 ;
        RECT 724.950 573.750 727.050 574.200 ;
        RECT 736.950 573.750 739.050 574.200 ;
        RECT 724.950 572.550 739.050 573.750 ;
        RECT 724.950 572.100 727.050 572.550 ;
        RECT 736.950 572.100 739.050 572.550 ;
        RECT 775.950 573.600 778.050 574.200 ;
        RECT 784.950 573.600 787.050 574.050 ;
        RECT 815.400 573.600 816.600 574.950 ;
        RECT 775.950 572.400 787.050 573.600 ;
        RECT 775.950 572.100 778.050 572.400 ;
        RECT 784.950 571.950 787.050 572.400 ;
        RECT 791.400 572.400 816.600 573.600 ;
        RECT 868.950 573.600 871.050 574.050 ;
        RECT 874.950 573.600 877.050 574.050 ;
        RECT 892.950 573.600 895.050 574.050 ;
        RECT 907.950 573.600 910.050 574.200 ;
        RECT 868.950 572.400 877.050 573.600 ;
        RECT 556.950 567.600 559.050 567.900 ;
        RECT 544.950 566.400 559.050 567.600 ;
        RECT 544.950 565.950 547.050 566.400 ;
        RECT 556.950 565.800 559.050 566.400 ;
        RECT 568.950 567.600 571.050 567.900 ;
        RECT 616.950 567.600 619.050 567.900 ;
        RECT 568.950 566.400 619.050 567.600 ;
        RECT 568.950 565.800 571.050 566.400 ;
        RECT 616.950 565.800 619.050 566.400 ;
        RECT 640.950 565.800 643.050 567.900 ;
        RECT 655.950 567.600 658.050 568.050 ;
        RECT 695.400 567.900 696.600 571.950 ;
        RECT 791.400 570.600 792.600 572.400 ;
        RECT 868.950 571.950 871.050 572.400 ;
        RECT 874.950 571.950 877.050 572.400 ;
        RECT 884.400 572.400 910.050 573.600 ;
        RECT 865.950 570.600 868.050 571.050 ;
        RECT 782.400 570.000 792.600 570.600 ;
        RECT 781.950 569.400 792.600 570.000 ;
        RECT 854.400 569.400 868.050 570.600 ;
        RECT 670.950 567.600 673.050 567.900 ;
        RECT 655.950 566.400 673.050 567.600 ;
        RECT 655.950 565.950 658.050 566.400 ;
        RECT 670.950 565.800 673.050 566.400 ;
        RECT 676.950 567.450 679.050 567.900 ;
        RECT 682.950 567.450 685.050 567.900 ;
        RECT 676.950 566.250 685.050 567.450 ;
        RECT 676.950 565.800 679.050 566.250 ;
        RECT 682.950 565.800 685.050 566.250 ;
        RECT 694.950 565.800 697.050 567.900 ;
        RECT 700.950 567.600 703.050 567.900 ;
        RECT 721.950 567.600 724.050 567.900 ;
        RECT 700.950 566.400 724.050 567.600 ;
        RECT 700.950 565.800 703.050 566.400 ;
        RECT 721.950 565.800 724.050 566.400 ;
        RECT 730.950 567.600 733.050 567.900 ;
        RECT 739.950 567.600 742.050 567.900 ;
        RECT 730.950 567.450 742.050 567.600 ;
        RECT 748.950 567.450 751.050 567.900 ;
        RECT 730.950 566.400 751.050 567.450 ;
        RECT 730.950 565.800 733.050 566.400 ;
        RECT 739.950 566.250 751.050 566.400 ;
        RECT 739.950 565.800 742.050 566.250 ;
        RECT 748.950 565.800 751.050 566.250 ;
        RECT 763.950 567.450 766.050 567.900 ;
        RECT 772.950 567.450 775.050 567.900 ;
        RECT 763.950 566.250 775.050 567.450 ;
        RECT 763.950 565.800 766.050 566.250 ;
        RECT 772.950 565.800 775.050 566.250 ;
        RECT 781.950 565.950 784.050 569.400 ;
        RECT 811.950 567.450 814.050 567.900 ;
        RECT 817.950 567.450 820.050 567.900 ;
        RECT 811.950 566.250 820.050 567.450 ;
        RECT 811.950 565.800 814.050 566.250 ;
        RECT 817.950 565.800 820.050 566.250 ;
        RECT 478.950 564.600 481.050 565.050 ;
        RECT 508.950 564.600 511.050 565.050 ;
        RECT 535.950 564.600 538.050 565.050 ;
        RECT 437.400 564.000 462.600 564.600 ;
        RECT 437.400 563.400 463.050 564.000 ;
        RECT 109.950 562.800 112.050 563.250 ;
        RECT 154.950 562.800 157.050 563.250 ;
        RECT 106.950 561.600 109.050 562.050 ;
        RECT 127.950 561.600 130.050 562.050 ;
        RECT 106.950 560.400 130.050 561.600 ;
        RECT 106.950 559.950 109.050 560.400 ;
        RECT 127.950 559.950 130.050 560.400 ;
        RECT 220.950 561.600 223.050 562.050 ;
        RECT 304.950 561.600 307.050 561.900 ;
        RECT 220.950 560.400 307.050 561.600 ;
        RECT 220.950 559.950 223.050 560.400 ;
        RECT 304.950 559.800 307.050 560.400 ;
        RECT 331.950 561.600 334.050 562.050 ;
        RECT 364.950 561.600 367.050 562.050 ;
        RECT 331.950 560.400 367.050 561.600 ;
        RECT 331.950 559.950 334.050 560.400 ;
        RECT 364.950 559.950 367.050 560.400 ;
        RECT 460.950 559.950 463.050 563.400 ;
        RECT 478.950 563.400 511.050 564.600 ;
        RECT 478.950 562.950 481.050 563.400 ;
        RECT 508.950 562.950 511.050 563.400 ;
        RECT 512.400 563.400 538.050 564.600 ;
        RECT 499.950 561.600 502.050 562.050 ;
        RECT 512.400 561.600 513.600 563.400 ;
        RECT 535.950 562.950 538.050 563.400 ;
        RECT 652.950 564.600 655.050 565.050 ;
        RECT 667.950 564.600 670.050 565.050 ;
        RECT 652.950 563.400 670.050 564.600 ;
        RECT 652.950 562.950 655.050 563.400 ;
        RECT 667.950 562.950 670.050 563.400 ;
        RECT 712.950 564.600 715.050 565.050 ;
        RECT 724.950 564.600 727.050 565.050 ;
        RECT 712.950 563.400 727.050 564.600 ;
        RECT 712.950 562.950 715.050 563.400 ;
        RECT 724.950 562.950 727.050 563.400 ;
        RECT 775.950 564.600 778.050 565.050 ;
        RECT 808.950 564.600 811.050 565.050 ;
        RECT 854.400 564.600 855.600 569.400 ;
        RECT 865.950 568.950 868.050 569.400 ;
        RECT 884.400 567.900 885.600 572.400 ;
        RECT 892.950 571.950 895.050 572.400 ;
        RECT 907.950 572.100 910.050 572.400 ;
        RECT 925.950 571.800 928.050 575.400 ;
        RECT 931.950 574.950 934.050 575.400 ;
        RECT 952.950 576.600 955.050 577.050 ;
        RECT 964.950 576.600 967.050 576.900 ;
        RECT 952.950 575.400 967.050 576.600 ;
        RECT 952.950 574.950 955.050 575.400 ;
        RECT 964.950 574.800 967.050 575.400 ;
        RECT 970.950 576.600 973.050 577.050 ;
        RECT 970.950 575.400 993.600 576.600 ;
        RECT 970.950 574.950 973.050 575.400 ;
        RECT 943.950 570.600 946.050 574.050 ;
        RECT 955.950 573.600 958.050 574.050 ;
        RECT 988.950 573.600 991.050 574.200 ;
        RECT 955.950 572.400 963.600 573.600 ;
        RECT 955.950 571.950 958.050 572.400 ;
        RECT 943.950 570.000 957.600 570.600 ;
        RECT 944.400 569.400 958.050 570.000 ;
        RECT 883.950 565.800 886.050 567.900 ;
        RECT 919.950 567.600 922.050 568.050 ;
        RECT 937.950 567.600 940.050 567.900 ;
        RECT 919.950 566.400 940.050 567.600 ;
        RECT 919.950 565.950 922.050 566.400 ;
        RECT 937.950 565.800 940.050 566.400 ;
        RECT 955.950 565.950 958.050 569.400 ;
        RECT 962.400 567.900 963.600 572.400 ;
        RECT 968.400 572.400 991.050 573.600 ;
        RECT 992.400 573.600 993.600 575.400 ;
        RECT 1015.950 573.600 1018.050 574.200 ;
        RECT 1031.400 574.050 1032.600 578.400 ;
        RECT 1036.950 577.950 1039.050 578.400 ;
        RECT 992.400 572.400 1018.050 573.600 ;
        RECT 968.400 567.900 969.600 572.400 ;
        RECT 988.950 572.100 991.050 572.400 ;
        RECT 1015.950 572.100 1018.050 572.400 ;
        RECT 1027.950 572.400 1032.600 574.050 ;
        RECT 1016.400 570.600 1017.600 572.100 ;
        RECT 1027.950 571.950 1032.000 572.400 ;
        RECT 1036.800 572.100 1038.900 574.200 ;
        RECT 1016.400 570.000 1020.600 570.600 ;
        RECT 1016.400 569.400 1021.050 570.000 ;
        RECT 961.950 565.800 964.050 567.900 ;
        RECT 967.950 565.800 970.050 567.900 ;
        RECT 973.950 567.450 976.050 567.900 ;
        RECT 985.950 567.450 988.050 567.900 ;
        RECT 973.950 566.250 988.050 567.450 ;
        RECT 973.950 565.800 976.050 566.250 ;
        RECT 985.950 565.800 988.050 566.250 ;
        RECT 991.950 567.600 994.050 567.900 ;
        RECT 1003.950 567.600 1006.050 568.050 ;
        RECT 1012.950 567.600 1015.050 567.900 ;
        RECT 991.950 566.400 1015.050 567.600 ;
        RECT 991.950 565.800 994.050 566.400 ;
        RECT 1003.950 565.950 1006.050 566.400 ;
        RECT 1012.950 565.800 1015.050 566.400 ;
        RECT 1018.950 565.950 1021.050 569.400 ;
        RECT 1030.950 567.600 1033.050 568.050 ;
        RECT 1037.400 567.600 1038.600 572.100 ;
        RECT 1039.950 571.950 1042.050 574.050 ;
        RECT 1040.400 568.050 1041.600 571.950 ;
        RECT 1030.950 566.400 1038.600 567.600 ;
        RECT 1030.950 565.950 1033.050 566.400 ;
        RECT 1039.950 565.950 1042.050 568.050 ;
        RECT 775.950 563.400 855.600 564.600 ;
        RECT 859.950 564.600 862.050 565.050 ;
        RECT 871.950 564.600 874.050 565.050 ;
        RECT 859.950 563.400 874.050 564.600 ;
        RECT 775.950 562.950 778.050 563.400 ;
        RECT 808.950 562.950 811.050 563.400 ;
        RECT 859.950 562.950 862.050 563.400 ;
        RECT 871.950 562.950 874.050 563.400 ;
        RECT 913.950 564.600 916.050 565.050 ;
        RECT 931.950 564.600 934.050 565.050 ;
        RECT 913.950 563.400 934.050 564.600 ;
        RECT 913.950 562.950 916.050 563.400 ;
        RECT 931.950 562.950 934.050 563.400 ;
        RECT 967.950 564.600 970.050 564.750 ;
        RECT 979.950 564.600 982.050 565.050 ;
        RECT 967.950 563.400 982.050 564.600 ;
        RECT 967.950 562.650 970.050 563.400 ;
        RECT 979.950 562.950 982.050 563.400 ;
        RECT 499.950 560.400 513.600 561.600 ;
        RECT 514.950 561.600 517.050 562.050 ;
        RECT 577.950 561.600 580.050 562.050 ;
        RECT 514.950 560.400 580.050 561.600 ;
        RECT 499.950 559.950 502.050 560.400 ;
        RECT 514.950 559.950 517.050 560.400 ;
        RECT 577.950 559.950 580.050 560.400 ;
        RECT 649.950 561.600 652.050 562.050 ;
        RECT 676.950 561.600 679.050 562.050 ;
        RECT 649.950 560.400 679.050 561.600 ;
        RECT 649.950 559.950 652.050 560.400 ;
        RECT 676.950 559.950 679.050 560.400 ;
        RECT 688.950 561.600 691.050 562.050 ;
        RECT 694.950 561.600 697.050 562.050 ;
        RECT 688.950 560.400 697.050 561.600 ;
        RECT 688.950 559.950 691.050 560.400 ;
        RECT 694.950 559.950 697.050 560.400 ;
        RECT 736.950 561.600 739.050 562.050 ;
        RECT 754.950 561.600 757.050 562.050 ;
        RECT 781.950 561.600 784.050 562.050 ;
        RECT 736.950 560.400 784.050 561.600 ;
        RECT 736.950 559.950 739.050 560.400 ;
        RECT 754.950 559.950 757.050 560.400 ;
        RECT 781.950 559.950 784.050 560.400 ;
        RECT 865.950 561.600 868.050 562.050 ;
        RECT 898.950 561.600 901.050 562.050 ;
        RECT 952.950 561.600 955.050 562.050 ;
        RECT 964.950 561.600 967.050 562.050 ;
        RECT 865.950 560.400 901.050 561.600 ;
        RECT 865.950 559.950 868.050 560.400 ;
        RECT 898.950 559.950 901.050 560.400 ;
        RECT 935.400 560.400 945.600 561.600 ;
        RECT 935.400 559.050 936.600 560.400 ;
        RECT 136.950 558.600 139.050 559.050 ;
        RECT 217.950 558.600 220.050 559.050 ;
        RECT 136.950 557.400 220.050 558.600 ;
        RECT 136.950 556.950 139.050 557.400 ;
        RECT 217.950 556.950 220.050 557.400 ;
        RECT 226.950 558.600 229.050 559.050 ;
        RECT 289.950 558.600 292.050 559.050 ;
        RECT 226.950 557.400 292.050 558.600 ;
        RECT 226.950 556.950 229.050 557.400 ;
        RECT 289.950 556.950 292.050 557.400 ;
        RECT 337.950 558.600 340.050 559.050 ;
        RECT 343.950 558.600 346.050 559.050 ;
        RECT 337.950 557.400 346.050 558.600 ;
        RECT 337.950 556.950 340.050 557.400 ;
        RECT 343.950 556.950 346.050 557.400 ;
        RECT 361.950 558.600 364.050 559.050 ;
        RECT 436.950 558.600 439.050 559.050 ;
        RECT 361.950 557.400 439.050 558.600 ;
        RECT 361.950 556.950 364.050 557.400 ;
        RECT 436.950 556.950 439.050 557.400 ;
        RECT 442.950 558.600 445.050 559.050 ;
        RECT 457.950 558.600 460.050 559.050 ;
        RECT 442.950 557.400 460.050 558.600 ;
        RECT 442.950 556.950 445.050 557.400 ;
        RECT 457.950 556.950 460.050 557.400 ;
        RECT 484.950 558.600 487.050 559.050 ;
        RECT 616.950 558.600 619.050 559.050 ;
        RECT 484.950 557.400 619.050 558.600 ;
        RECT 484.950 556.950 487.050 557.400 ;
        RECT 616.950 556.950 619.050 557.400 ;
        RECT 646.950 558.600 649.050 559.050 ;
        RECT 709.950 558.600 712.050 559.050 ;
        RECT 646.950 557.400 712.050 558.600 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 709.950 556.950 712.050 557.400 ;
        RECT 742.950 558.600 745.050 559.050 ;
        RECT 778.800 558.600 780.900 559.050 ;
        RECT 742.950 557.400 780.900 558.600 ;
        RECT 742.950 556.950 745.050 557.400 ;
        RECT 778.800 556.950 780.900 557.400 ;
        RECT 781.950 558.600 784.050 558.900 ;
        RECT 832.800 558.600 834.900 559.050 ;
        RECT 781.950 557.400 834.900 558.600 ;
        RECT 781.950 556.800 784.050 557.400 ;
        RECT 832.800 556.950 834.900 557.400 ;
        RECT 835.950 558.600 838.050 559.050 ;
        RECT 850.950 558.600 853.050 559.050 ;
        RECT 835.950 557.400 853.050 558.600 ;
        RECT 835.950 556.950 838.050 557.400 ;
        RECT 850.950 556.950 853.050 557.400 ;
        RECT 862.950 558.600 865.050 559.050 ;
        RECT 892.950 558.600 895.050 559.050 ;
        RECT 862.950 557.400 895.050 558.600 ;
        RECT 862.950 556.950 865.050 557.400 ;
        RECT 892.950 556.950 895.050 557.400 ;
        RECT 898.950 558.600 901.050 558.900 ;
        RECT 916.950 558.600 919.050 559.050 ;
        RECT 898.950 557.400 919.050 558.600 ;
        RECT 898.950 556.800 901.050 557.400 ;
        RECT 916.950 556.950 919.050 557.400 ;
        RECT 931.950 557.400 936.600 559.050 ;
        RECT 944.400 558.600 945.600 560.400 ;
        RECT 952.950 560.400 967.050 561.600 ;
        RECT 952.950 559.950 955.050 560.400 ;
        RECT 964.950 559.950 967.050 560.400 ;
        RECT 961.950 558.600 964.050 559.050 ;
        RECT 944.400 557.400 964.050 558.600 ;
        RECT 931.950 556.950 936.000 557.400 ;
        RECT 961.950 556.950 964.050 557.400 ;
        RECT 976.950 558.600 979.050 559.050 ;
        RECT 1012.950 558.600 1015.050 559.050 ;
        RECT 976.950 557.400 1015.050 558.600 ;
        RECT 976.950 556.950 979.050 557.400 ;
        RECT 1012.950 556.950 1015.050 557.400 ;
        RECT 115.950 555.600 118.050 556.050 ;
        RECT 220.950 555.600 223.050 556.050 ;
        RECT 115.950 554.400 223.050 555.600 ;
        RECT 115.950 553.950 118.050 554.400 ;
        RECT 220.950 553.950 223.050 554.400 ;
        RECT 352.950 555.600 355.050 556.050 ;
        RECT 403.950 555.600 406.050 556.050 ;
        RECT 352.950 554.400 406.050 555.600 ;
        RECT 352.950 553.950 355.050 554.400 ;
        RECT 403.950 553.950 406.050 554.400 ;
        RECT 460.950 555.600 463.050 556.050 ;
        RECT 481.950 555.600 484.050 556.050 ;
        RECT 460.950 554.400 484.050 555.600 ;
        RECT 460.950 553.950 463.050 554.400 ;
        RECT 481.950 553.950 484.050 554.400 ;
        RECT 550.950 555.600 553.050 556.050 ;
        RECT 610.950 555.600 613.050 556.050 ;
        RECT 664.950 555.600 667.050 556.050 ;
        RECT 550.950 554.400 667.050 555.600 ;
        RECT 550.950 553.950 553.050 554.400 ;
        RECT 610.950 553.950 613.050 554.400 ;
        RECT 664.950 553.950 667.050 554.400 ;
        RECT 685.950 555.600 688.050 556.050 ;
        RECT 700.950 555.600 703.050 556.050 ;
        RECT 685.950 554.400 703.050 555.600 ;
        RECT 685.950 553.950 688.050 554.400 ;
        RECT 700.950 553.950 703.050 554.400 ;
        RECT 760.950 555.600 763.050 556.050 ;
        RECT 865.950 555.600 868.050 556.050 ;
        RECT 760.950 554.400 868.050 555.600 ;
        RECT 760.950 553.950 763.050 554.400 ;
        RECT 865.950 553.950 868.050 554.400 ;
        RECT 871.950 555.600 874.050 556.050 ;
        RECT 913.950 555.600 916.050 556.050 ;
        RECT 871.950 554.400 916.050 555.600 ;
        RECT 871.950 553.950 874.050 554.400 ;
        RECT 913.950 553.950 916.050 554.400 ;
        RECT 940.950 555.600 943.050 556.050 ;
        RECT 970.950 555.600 973.050 556.050 ;
        RECT 940.950 554.400 973.050 555.600 ;
        RECT 940.950 553.950 943.050 554.400 ;
        RECT 970.950 553.950 973.050 554.400 ;
        RECT 202.950 552.600 205.050 553.050 ;
        RECT 244.950 552.600 247.050 553.050 ;
        RECT 202.950 551.400 247.050 552.600 ;
        RECT 202.950 550.950 205.050 551.400 ;
        RECT 244.950 550.950 247.050 551.400 ;
        RECT 277.950 552.600 280.050 553.050 ;
        RECT 355.950 552.600 358.050 553.050 ;
        RECT 277.950 551.400 358.050 552.600 ;
        RECT 277.950 550.950 280.050 551.400 ;
        RECT 355.950 550.950 358.050 551.400 ;
        RECT 547.950 552.600 550.050 553.050 ;
        RECT 580.950 552.600 583.050 553.050 ;
        RECT 547.950 551.400 583.050 552.600 ;
        RECT 547.950 550.950 550.050 551.400 ;
        RECT 580.950 550.950 583.050 551.400 ;
        RECT 667.950 552.600 670.050 553.050 ;
        RECT 706.950 552.600 709.050 553.050 ;
        RECT 667.950 551.400 709.050 552.600 ;
        RECT 667.950 550.950 670.050 551.400 ;
        RECT 706.950 550.950 709.050 551.400 ;
        RECT 772.950 552.600 775.050 553.050 ;
        RECT 784.950 552.600 787.050 553.050 ;
        RECT 772.950 551.400 787.050 552.600 ;
        RECT 772.950 550.950 775.050 551.400 ;
        RECT 784.950 550.950 787.050 551.400 ;
        RECT 847.950 552.600 850.050 553.050 ;
        RECT 919.950 552.600 922.050 553.050 ;
        RECT 925.800 552.600 927.900 553.050 ;
        RECT 847.950 551.400 906.600 552.600 ;
        RECT 847.950 550.950 850.050 551.400 ;
        RECT 295.950 549.600 298.050 550.050 ;
        RECT 325.950 549.600 328.050 550.050 ;
        RECT 394.950 549.600 397.050 550.050 ;
        RECT 295.950 548.400 328.050 549.600 ;
        RECT 295.950 547.950 298.050 548.400 ;
        RECT 325.950 547.950 328.050 548.400 ;
        RECT 329.400 548.400 397.050 549.600 ;
        RECT 16.950 546.600 19.050 547.050 ;
        RECT 64.950 546.600 67.050 547.050 ;
        RECT 70.950 546.600 73.050 547.050 ;
        RECT 16.950 545.400 73.050 546.600 ;
        RECT 16.950 544.950 19.050 545.400 ;
        RECT 64.950 544.950 67.050 545.400 ;
        RECT 70.950 544.950 73.050 545.400 ;
        RECT 76.950 546.600 79.050 547.050 ;
        RECT 193.950 546.600 196.050 547.050 ;
        RECT 76.950 545.400 196.050 546.600 ;
        RECT 76.950 544.950 79.050 545.400 ;
        RECT 193.950 544.950 196.050 545.400 ;
        RECT 259.950 546.600 262.050 547.050 ;
        RECT 329.400 546.600 330.600 548.400 ;
        RECT 394.950 547.950 397.050 548.400 ;
        RECT 415.950 549.600 418.050 550.050 ;
        RECT 436.950 549.600 439.050 550.050 ;
        RECT 415.950 548.400 439.050 549.600 ;
        RECT 415.950 547.950 418.050 548.400 ;
        RECT 436.950 547.950 439.050 548.400 ;
        RECT 481.950 549.600 484.050 550.050 ;
        RECT 520.950 549.600 523.050 550.050 ;
        RECT 541.950 549.600 544.050 550.050 ;
        RECT 589.950 549.600 592.050 550.050 ;
        RECT 649.950 549.600 652.050 550.050 ;
        RECT 481.950 548.400 652.050 549.600 ;
        RECT 481.950 547.950 484.050 548.400 ;
        RECT 520.950 547.950 523.050 548.400 ;
        RECT 541.950 547.950 544.050 548.400 ;
        RECT 589.950 547.950 592.050 548.400 ;
        RECT 649.950 547.950 652.050 548.400 ;
        RECT 667.950 549.600 670.050 549.900 ;
        RECT 703.950 549.600 706.050 550.050 ;
        RECT 667.950 548.400 706.050 549.600 ;
        RECT 667.950 547.800 670.050 548.400 ;
        RECT 703.950 547.950 706.050 548.400 ;
        RECT 709.950 549.600 712.050 550.050 ;
        RECT 727.950 549.600 730.050 550.050 ;
        RECT 859.950 549.600 862.050 550.050 ;
        RECT 709.950 548.400 730.050 549.600 ;
        RECT 709.950 547.950 712.050 548.400 ;
        RECT 727.950 547.950 730.050 548.400 ;
        RECT 800.400 548.400 862.050 549.600 ;
        RECT 800.400 547.050 801.600 548.400 ;
        RECT 859.950 547.950 862.050 548.400 ;
        RECT 877.950 549.600 880.050 550.050 ;
        RECT 898.950 549.600 901.050 550.050 ;
        RECT 877.950 548.400 901.050 549.600 ;
        RECT 905.400 549.600 906.600 551.400 ;
        RECT 919.950 551.400 927.900 552.600 ;
        RECT 919.950 550.950 922.050 551.400 ;
        RECT 925.800 550.950 927.900 551.400 ;
        RECT 928.950 552.600 931.050 553.050 ;
        RECT 943.950 552.600 946.050 553.050 ;
        RECT 928.950 551.400 946.050 552.600 ;
        RECT 928.950 550.950 931.050 551.400 ;
        RECT 943.950 550.950 946.050 551.400 ;
        RECT 970.950 552.600 973.050 552.900 ;
        RECT 997.950 552.600 1000.050 553.050 ;
        RECT 970.950 551.400 1000.050 552.600 ;
        RECT 970.950 550.800 973.050 551.400 ;
        RECT 997.950 550.950 1000.050 551.400 ;
        RECT 913.950 549.600 916.050 550.050 ;
        RECT 946.950 549.600 949.050 550.050 ;
        RECT 905.400 548.400 949.050 549.600 ;
        RECT 877.950 547.950 880.050 548.400 ;
        RECT 898.950 547.950 901.050 548.400 ;
        RECT 913.950 547.950 916.050 548.400 ;
        RECT 946.950 547.950 949.050 548.400 ;
        RECT 955.950 549.600 958.050 550.050 ;
        RECT 961.950 549.600 964.050 550.050 ;
        RECT 976.950 549.600 979.050 550.050 ;
        RECT 955.950 548.400 979.050 549.600 ;
        RECT 955.950 547.950 958.050 548.400 ;
        RECT 961.950 547.950 964.050 548.400 ;
        RECT 976.950 547.950 979.050 548.400 ;
        RECT 1000.950 549.600 1003.050 549.900 ;
        RECT 1024.950 549.600 1027.050 550.050 ;
        RECT 1000.950 548.400 1027.050 549.600 ;
        RECT 1000.950 547.800 1003.050 548.400 ;
        RECT 1024.950 547.950 1027.050 548.400 ;
        RECT 259.950 545.400 330.600 546.600 ;
        RECT 376.950 546.600 379.050 547.050 ;
        RECT 493.950 546.600 496.050 547.050 ;
        RECT 562.950 546.600 565.050 547.050 ;
        RECT 376.950 545.400 496.050 546.600 ;
        RECT 259.950 544.950 262.050 545.400 ;
        RECT 376.950 544.950 379.050 545.400 ;
        RECT 493.950 544.950 496.050 545.400 ;
        RECT 497.400 545.400 565.050 546.600 ;
        RECT 256.950 543.600 259.050 544.050 ;
        RECT 406.950 543.600 409.050 544.050 ;
        RECT 256.950 542.400 409.050 543.600 ;
        RECT 256.950 541.950 259.050 542.400 ;
        RECT 406.950 541.950 409.050 542.400 ;
        RECT 427.950 543.600 430.050 544.050 ;
        RECT 439.950 543.600 442.050 544.050 ;
        RECT 497.400 543.600 498.600 545.400 ;
        RECT 562.950 544.950 565.050 545.400 ;
        RECT 625.950 546.600 628.050 547.050 ;
        RECT 637.950 546.600 640.050 547.050 ;
        RECT 625.950 545.400 640.050 546.600 ;
        RECT 625.950 544.950 628.050 545.400 ;
        RECT 637.950 544.950 640.050 545.400 ;
        RECT 664.950 546.600 667.050 547.050 ;
        RECT 799.950 546.600 802.050 547.050 ;
        RECT 664.950 545.400 802.050 546.600 ;
        RECT 664.950 544.950 667.050 545.400 ;
        RECT 799.950 544.950 802.050 545.400 ;
        RECT 832.950 546.600 835.050 547.050 ;
        RECT 853.950 546.600 856.050 547.050 ;
        RECT 832.950 545.400 856.050 546.600 ;
        RECT 832.950 544.950 835.050 545.400 ;
        RECT 853.950 544.950 856.050 545.400 ;
        RECT 982.950 546.600 985.050 547.050 ;
        RECT 1033.950 546.600 1036.050 547.050 ;
        RECT 982.950 545.400 1036.050 546.600 ;
        RECT 982.950 544.950 985.050 545.400 ;
        RECT 1033.950 544.950 1036.050 545.400 ;
        RECT 427.950 542.400 498.600 543.600 ;
        RECT 520.950 543.600 523.050 544.050 ;
        RECT 544.950 543.600 547.050 544.050 ;
        RECT 520.950 542.400 547.050 543.600 ;
        RECT 427.950 541.950 430.050 542.400 ;
        RECT 439.950 541.950 442.050 542.400 ;
        RECT 520.950 541.950 523.050 542.400 ;
        RECT 544.950 541.950 547.050 542.400 ;
        RECT 574.950 543.600 577.050 544.050 ;
        RECT 586.950 543.600 589.050 544.050 ;
        RECT 574.950 542.400 589.050 543.600 ;
        RECT 574.950 541.950 577.050 542.400 ;
        RECT 586.950 541.950 589.050 542.400 ;
        RECT 610.950 543.600 613.050 544.050 ;
        RECT 661.950 543.600 664.050 544.050 ;
        RECT 610.950 542.400 664.050 543.600 ;
        RECT 610.950 541.950 613.050 542.400 ;
        RECT 661.950 541.950 664.050 542.400 ;
        RECT 676.950 543.600 679.050 544.050 ;
        RECT 697.950 543.600 700.050 544.050 ;
        RECT 676.950 542.400 700.050 543.600 ;
        RECT 676.950 541.950 679.050 542.400 ;
        RECT 697.950 541.950 700.050 542.400 ;
        RECT 703.950 543.600 706.050 544.050 ;
        RECT 709.950 543.600 712.050 544.050 ;
        RECT 775.950 543.600 778.050 544.050 ;
        RECT 886.950 543.600 889.050 544.050 ;
        RECT 703.950 542.400 712.050 543.600 ;
        RECT 703.950 541.950 706.050 542.400 ;
        RECT 709.950 541.950 712.050 542.400 ;
        RECT 716.400 542.400 778.050 543.600 ;
        RECT 73.950 540.600 76.050 541.050 ;
        RECT 88.950 540.600 91.050 541.050 ;
        RECT 73.950 539.400 91.050 540.600 ;
        RECT 73.950 538.950 76.050 539.400 ;
        RECT 88.950 538.950 91.050 539.400 ;
        RECT 103.950 540.600 106.050 541.050 ;
        RECT 112.950 540.600 115.050 541.050 ;
        RECT 103.950 539.400 115.050 540.600 ;
        RECT 103.950 538.950 106.050 539.400 ;
        RECT 112.950 538.950 115.050 539.400 ;
        RECT 124.950 540.600 127.050 541.050 ;
        RECT 133.950 540.600 136.050 541.050 ;
        RECT 124.950 539.400 136.050 540.600 ;
        RECT 124.950 538.950 127.050 539.400 ;
        RECT 133.950 538.950 136.050 539.400 ;
        RECT 193.950 540.600 196.050 540.900 ;
        RECT 208.950 540.600 211.050 541.050 ;
        RECT 457.950 540.600 460.050 541.050 ;
        RECT 526.950 540.600 529.050 541.050 ;
        RECT 193.950 539.400 211.050 540.600 ;
        RECT 193.950 538.800 196.050 539.400 ;
        RECT 208.950 538.950 211.050 539.400 ;
        RECT 401.400 539.400 529.050 540.600 ;
        RECT 401.400 538.050 402.600 539.400 ;
        RECT 457.950 538.950 460.050 539.400 ;
        RECT 526.950 538.950 529.050 539.400 ;
        RECT 616.950 540.600 619.050 541.050 ;
        RECT 661.950 540.600 664.050 540.900 ;
        RECT 616.950 539.400 664.050 540.600 ;
        RECT 616.950 538.950 619.050 539.400 ;
        RECT 661.950 538.800 664.050 539.400 ;
        RECT 706.950 540.600 709.050 541.050 ;
        RECT 716.400 540.600 717.600 542.400 ;
        RECT 775.950 541.950 778.050 542.400 ;
        RECT 827.400 542.400 889.050 543.600 ;
        RECT 706.950 539.400 717.600 540.600 ;
        RECT 769.950 540.600 772.050 541.050 ;
        RECT 827.400 540.600 828.600 542.400 ;
        RECT 886.950 541.950 889.050 542.400 ;
        RECT 769.950 539.400 828.600 540.600 ;
        RECT 835.950 540.600 838.050 541.050 ;
        RECT 844.950 540.600 847.050 541.050 ;
        RECT 871.950 540.600 874.050 541.050 ;
        RECT 835.950 539.400 874.050 540.600 ;
        RECT 706.950 538.950 709.050 539.400 ;
        RECT 769.950 538.950 772.050 539.400 ;
        RECT 835.950 538.950 838.050 539.400 ;
        RECT 844.950 538.950 847.050 539.400 ;
        RECT 871.950 538.950 874.050 539.400 ;
        RECT 916.950 540.600 919.050 541.050 ;
        RECT 922.950 540.600 925.050 541.050 ;
        RECT 916.950 539.400 925.050 540.600 ;
        RECT 916.950 538.950 919.050 539.400 ;
        RECT 922.950 538.950 925.050 539.400 ;
        RECT 100.950 537.600 103.050 538.050 ;
        RECT 26.400 537.000 103.050 537.600 ;
        RECT 25.950 536.400 103.050 537.000 ;
        RECT 25.950 532.950 28.050 536.400 ;
        RECT 100.950 535.950 103.050 536.400 ;
        RECT 163.950 537.600 166.050 538.050 ;
        RECT 172.950 537.600 175.050 538.050 ;
        RECT 208.950 537.600 211.050 537.900 ;
        RECT 163.950 536.400 211.050 537.600 ;
        RECT 163.950 535.950 166.050 536.400 ;
        RECT 172.950 535.950 175.050 536.400 ;
        RECT 208.950 535.800 211.050 536.400 ;
        RECT 262.950 537.600 265.050 538.050 ;
        RECT 319.950 537.600 322.050 538.050 ;
        RECT 262.950 536.400 322.050 537.600 ;
        RECT 262.950 535.950 265.050 536.400 ;
        RECT 319.950 535.950 322.050 536.400 ;
        RECT 391.950 537.600 394.050 538.050 ;
        RECT 400.950 537.600 403.050 538.050 ;
        RECT 391.950 536.400 403.050 537.600 ;
        RECT 391.950 535.950 394.050 536.400 ;
        RECT 400.950 535.950 403.050 536.400 ;
        RECT 628.950 537.600 631.050 538.050 ;
        RECT 670.950 537.600 673.050 538.050 ;
        RECT 628.950 536.400 673.050 537.600 ;
        RECT 628.950 535.950 631.050 536.400 ;
        RECT 670.950 535.950 673.050 536.400 ;
        RECT 715.950 537.600 718.050 538.050 ;
        RECT 733.950 537.600 736.050 538.050 ;
        RECT 754.950 537.600 757.050 538.050 ;
        RECT 715.950 536.400 757.050 537.600 ;
        RECT 715.950 535.950 718.050 536.400 ;
        RECT 733.950 535.950 736.050 536.400 ;
        RECT 754.950 535.950 757.050 536.400 ;
        RECT 811.950 537.600 814.050 538.050 ;
        RECT 829.950 537.600 832.050 538.050 ;
        RECT 877.950 537.600 880.050 538.050 ;
        RECT 811.950 536.400 880.050 537.600 ;
        RECT 811.950 535.950 814.050 536.400 ;
        RECT 829.950 535.950 832.050 536.400 ;
        RECT 877.950 535.950 880.050 536.400 ;
        RECT 937.950 537.600 940.050 538.050 ;
        RECT 955.950 537.600 958.050 538.050 ;
        RECT 937.950 536.400 958.050 537.600 ;
        RECT 937.950 535.950 940.050 536.400 ;
        RECT 955.950 535.950 958.050 536.400 ;
        RECT 112.950 534.600 115.050 535.050 ;
        RECT 130.950 534.600 133.050 535.050 ;
        RECT 136.950 534.600 139.050 535.050 ;
        RECT 112.950 533.400 139.050 534.600 ;
        RECT 112.950 532.950 115.050 533.400 ;
        RECT 130.950 532.950 133.050 533.400 ;
        RECT 136.950 532.950 139.050 533.400 ;
        RECT 421.950 534.600 424.050 535.050 ;
        RECT 433.950 534.600 436.050 535.050 ;
        RECT 421.950 533.400 436.050 534.600 ;
        RECT 421.950 532.950 424.050 533.400 ;
        RECT 433.950 532.950 436.050 533.400 ;
        RECT 487.950 534.600 490.050 535.050 ;
        RECT 502.950 534.600 505.050 535.050 ;
        RECT 487.950 533.400 505.050 534.600 ;
        RECT 487.950 532.950 490.050 533.400 ;
        RECT 502.950 532.950 505.050 533.400 ;
        RECT 655.950 534.600 658.050 535.050 ;
        RECT 679.950 534.600 682.050 535.050 ;
        RECT 655.950 533.400 682.050 534.600 ;
        RECT 655.950 532.950 658.050 533.400 ;
        RECT 679.950 532.950 682.050 533.400 ;
        RECT 718.950 534.600 721.050 535.050 ;
        RECT 730.800 534.600 732.900 535.050 ;
        RECT 718.950 533.400 732.900 534.600 ;
        RECT 718.950 532.950 721.050 533.400 ;
        RECT 730.800 532.950 732.900 533.400 ;
        RECT 733.950 534.600 736.050 534.900 ;
        RECT 769.950 534.600 772.050 535.050 ;
        RECT 733.950 533.400 772.050 534.600 ;
        RECT 733.950 532.800 736.050 533.400 ;
        RECT 769.950 532.950 772.050 533.400 ;
        RECT 832.950 534.600 835.050 535.050 ;
        RECT 850.950 534.600 853.050 535.050 ;
        RECT 871.950 534.600 874.050 535.050 ;
        RECT 889.950 534.600 892.050 535.050 ;
        RECT 832.950 533.400 892.050 534.600 ;
        RECT 832.950 532.950 835.050 533.400 ;
        RECT 850.950 532.950 853.050 533.400 ;
        RECT 871.950 532.950 874.050 533.400 ;
        RECT 889.950 532.950 892.050 533.400 ;
        RECT 901.950 534.600 904.050 535.050 ;
        RECT 910.950 534.600 913.050 535.050 ;
        RECT 901.950 533.400 913.050 534.600 ;
        RECT 901.950 532.950 904.050 533.400 ;
        RECT 910.950 532.950 913.050 533.400 ;
        RECT 4.950 531.600 7.050 532.200 ;
        RECT 13.950 531.600 16.050 532.050 ;
        RECT 4.950 530.400 16.050 531.600 ;
        RECT 4.950 530.100 7.050 530.400 ;
        RECT 13.950 529.950 16.050 530.400 ;
        RECT 238.950 531.600 241.050 532.050 ;
        RECT 256.950 531.600 259.050 532.050 ;
        RECT 238.950 530.400 259.050 531.600 ;
        RECT 238.950 529.950 241.050 530.400 ;
        RECT 256.950 529.950 259.050 530.400 ;
        RECT 277.950 531.600 280.050 532.050 ;
        RECT 283.950 531.600 286.050 532.050 ;
        RECT 277.950 530.400 286.050 531.600 ;
        RECT 277.950 529.950 280.050 530.400 ;
        RECT 283.950 529.950 286.050 530.400 ;
        RECT 298.950 531.600 301.050 532.050 ;
        RECT 337.950 531.600 340.050 532.050 ;
        RECT 364.950 531.600 367.050 532.050 ;
        RECT 394.950 531.600 397.050 532.050 ;
        RECT 298.950 530.400 315.600 531.600 ;
        RECT 298.950 529.950 301.050 530.400 ;
        RECT 28.950 525.600 31.050 529.050 ;
        RECT 94.950 528.600 97.050 529.200 ;
        RECT 115.950 528.600 118.050 529.200 ;
        RECT 94.950 527.400 118.050 528.600 ;
        RECT 94.950 527.100 97.050 527.400 ;
        RECT 115.950 527.100 118.050 527.400 ;
        RECT 142.950 528.750 145.050 529.200 ;
        RECT 148.950 528.750 151.050 529.200 ;
        RECT 142.950 527.550 151.050 528.750 ;
        RECT 142.950 527.100 145.050 527.550 ;
        RECT 148.950 527.100 151.050 527.550 ;
        RECT 163.950 528.600 166.050 529.200 ;
        RECT 175.950 528.600 178.050 529.050 ;
        RECT 187.950 528.600 190.050 529.200 ;
        RECT 163.950 527.400 190.050 528.600 ;
        RECT 163.950 527.100 166.050 527.400 ;
        RECT 175.950 526.950 178.050 527.400 ;
        RECT 187.950 527.100 190.050 527.400 ;
        RECT 199.950 528.750 202.050 529.200 ;
        RECT 214.950 528.750 217.050 529.200 ;
        RECT 199.950 527.550 217.050 528.750 ;
        RECT 199.950 527.100 202.050 527.550 ;
        RECT 214.950 527.100 217.050 527.550 ;
        RECT 229.950 528.600 232.050 529.050 ;
        RECT 250.950 528.600 253.050 529.050 ;
        RECT 229.950 527.400 253.050 528.600 ;
        RECT 314.400 528.600 315.600 530.400 ;
        RECT 337.950 530.400 397.050 531.600 ;
        RECT 337.950 529.950 340.050 530.400 ;
        RECT 364.950 529.950 367.050 530.400 ;
        RECT 394.950 529.950 397.050 530.400 ;
        RECT 409.950 531.600 412.050 532.050 ;
        RECT 418.950 531.600 421.050 531.900 ;
        RECT 454.950 531.600 457.050 532.050 ;
        RECT 409.950 530.400 457.050 531.600 ;
        RECT 409.950 529.950 412.050 530.400 ;
        RECT 418.950 529.800 421.050 530.400 ;
        RECT 454.950 529.950 457.050 530.400 ;
        RECT 460.950 531.600 463.050 532.050 ;
        RECT 466.950 531.600 469.050 532.050 ;
        RECT 475.950 531.600 478.050 532.050 ;
        RECT 460.950 530.400 478.050 531.600 ;
        RECT 460.950 529.950 463.050 530.400 ;
        RECT 466.950 529.950 469.050 530.400 ;
        RECT 475.950 529.950 478.050 530.400 ;
        RECT 496.950 531.600 499.050 532.050 ;
        RECT 547.950 531.600 550.050 532.050 ;
        RECT 496.950 530.400 504.600 531.600 ;
        RECT 496.950 529.950 499.050 530.400 ;
        RECT 316.950 528.600 319.050 529.200 ;
        RECT 314.400 527.400 319.050 528.600 ;
        RECT 229.950 526.950 232.050 527.400 ;
        RECT 250.950 526.950 253.050 527.400 ;
        RECT 316.950 527.100 319.050 527.400 ;
        RECT 373.950 528.600 376.050 529.200 ;
        RECT 382.950 528.600 385.050 529.050 ;
        RECT 373.950 527.400 385.050 528.600 ;
        RECT 373.950 527.100 376.050 527.400 ;
        RECT 382.950 526.950 385.050 527.400 ;
        RECT 424.950 528.600 427.050 529.200 ;
        RECT 448.950 528.600 451.050 529.200 ;
        RECT 424.950 527.400 451.050 528.600 ;
        RECT 424.950 527.100 427.050 527.400 ;
        RECT 448.950 527.100 451.050 527.400 ;
        RECT 469.950 527.100 472.050 529.200 ;
        RECT 52.950 525.600 55.050 526.050 ;
        RECT 331.950 525.600 334.050 526.050 ;
        RECT 28.950 525.000 55.050 525.600 ;
        RECT 29.400 524.400 55.050 525.000 ;
        RECT 52.950 523.950 55.050 524.400 ;
        RECT 326.400 524.400 334.050 525.600 ;
        RECT 79.950 522.600 82.050 523.050 ;
        RECT 85.950 522.600 88.050 522.900 ;
        RECT 79.950 521.400 88.050 522.600 ;
        RECT 79.950 520.950 82.050 521.400 ;
        RECT 85.950 520.800 88.050 521.400 ;
        RECT 100.950 522.600 103.050 523.050 ;
        RECT 133.950 522.600 136.050 522.900 ;
        RECT 100.950 521.400 136.050 522.600 ;
        RECT 100.950 520.950 103.050 521.400 ;
        RECT 133.950 520.800 136.050 521.400 ;
        RECT 205.950 522.600 208.050 522.900 ;
        RECT 223.950 522.600 226.050 523.050 ;
        RECT 205.950 521.400 226.050 522.600 ;
        RECT 205.950 520.800 208.050 521.400 ;
        RECT 223.950 520.950 226.050 521.400 ;
        RECT 271.950 522.600 274.050 523.050 ;
        RECT 280.950 522.600 283.050 523.050 ;
        RECT 271.950 521.400 283.050 522.600 ;
        RECT 271.950 520.950 274.050 521.400 ;
        RECT 280.950 520.950 283.050 521.400 ;
        RECT 313.950 522.600 316.050 522.900 ;
        RECT 326.400 522.600 327.600 524.400 ;
        RECT 331.950 523.950 334.050 524.400 ;
        RECT 313.950 521.400 327.600 522.600 ;
        RECT 406.950 522.600 409.050 523.050 ;
        RECT 421.950 522.600 424.050 522.900 ;
        RECT 406.950 521.400 424.050 522.600 ;
        RECT 313.950 520.800 316.050 521.400 ;
        RECT 406.950 520.950 409.050 521.400 ;
        RECT 421.950 520.800 424.050 521.400 ;
        RECT 427.950 522.450 430.050 522.900 ;
        RECT 433.950 522.450 436.050 522.900 ;
        RECT 427.950 521.250 436.050 522.450 ;
        RECT 427.950 520.800 430.050 521.250 ;
        RECT 433.950 520.800 436.050 521.250 ;
        RECT 439.950 522.450 442.050 522.900 ;
        RECT 445.950 522.450 448.050 522.900 ;
        RECT 439.950 521.250 448.050 522.450 ;
        RECT 439.950 520.800 442.050 521.250 ;
        RECT 445.950 520.800 448.050 521.250 ;
        RECT 454.950 522.600 457.050 523.050 ;
        RECT 466.950 522.600 469.050 522.900 ;
        RECT 454.950 521.400 469.050 522.600 ;
        RECT 454.950 520.950 457.050 521.400 ;
        RECT 466.950 520.800 469.050 521.400 ;
        RECT 470.400 520.050 471.600 527.100 ;
        RECT 472.950 522.450 475.050 522.900 ;
        RECT 478.800 522.450 480.900 522.900 ;
        RECT 472.950 521.250 480.900 522.450 ;
        RECT 472.950 520.800 475.050 521.250 ;
        RECT 478.800 520.800 480.900 521.250 ;
        RECT 481.950 522.600 484.050 523.050 ;
        RECT 490.950 522.600 493.050 523.050 ;
        RECT 503.400 522.900 504.600 530.400 ;
        RECT 539.400 530.400 550.050 531.600 ;
        RECT 535.950 525.600 538.050 525.900 ;
        RECT 539.400 525.600 540.600 530.400 ;
        RECT 547.950 529.950 550.050 530.400 ;
        RECT 595.950 531.750 598.050 532.200 ;
        RECT 601.950 531.750 604.050 532.200 ;
        RECT 595.950 530.550 604.050 531.750 ;
        RECT 595.950 530.100 598.050 530.550 ;
        RECT 601.950 530.100 604.050 530.550 ;
        RECT 610.950 528.600 613.050 529.050 ;
        RECT 631.950 528.600 634.050 529.200 ;
        RECT 610.950 527.400 634.050 528.600 ;
        RECT 610.950 526.950 613.050 527.400 ;
        RECT 631.950 527.100 634.050 527.400 ;
        RECT 640.950 528.600 643.050 529.050 ;
        RECT 658.950 528.600 661.050 532.050 ;
        RECT 673.950 531.600 676.050 532.050 ;
        RECT 682.950 531.600 685.050 532.050 ;
        RECT 718.950 531.600 721.050 531.900 ;
        RECT 673.950 530.400 685.050 531.600 ;
        RECT 673.950 529.950 676.050 530.400 ;
        RECT 682.950 529.950 685.050 530.400 ;
        RECT 713.400 530.400 721.050 531.600 ;
        RECT 703.950 528.600 706.050 529.050 ;
        RECT 709.950 528.600 712.050 529.200 ;
        RECT 713.400 528.600 714.600 530.400 ;
        RECT 718.950 529.800 721.050 530.400 ;
        RECT 757.950 531.600 760.050 532.050 ;
        RECT 772.950 531.600 775.050 532.050 ;
        RECT 757.950 530.400 775.050 531.600 ;
        RECT 757.950 529.950 760.050 530.400 ;
        RECT 772.950 529.950 775.050 530.400 ;
        RECT 823.950 531.600 826.050 532.050 ;
        RECT 841.950 531.600 844.050 532.050 ;
        RECT 868.950 531.600 871.050 532.050 ;
        RECT 823.950 530.400 871.050 531.600 ;
        RECT 823.950 529.950 826.050 530.400 ;
        RECT 841.950 529.950 844.050 530.400 ;
        RECT 868.950 529.950 871.050 530.400 ;
        RECT 640.950 527.400 693.600 528.600 ;
        RECT 640.950 526.950 643.050 527.400 ;
        RECT 550.950 525.750 553.050 526.200 ;
        RECT 571.950 525.750 574.050 526.200 ;
        RECT 518.400 525.000 549.600 525.600 ;
        RECT 517.950 524.400 549.600 525.000 ;
        RECT 481.950 521.400 493.050 522.600 ;
        RECT 481.950 520.950 484.050 521.400 ;
        RECT 490.950 520.950 493.050 521.400 ;
        RECT 502.950 520.800 505.050 522.900 ;
        RECT 517.950 520.950 520.050 524.400 ;
        RECT 535.950 523.800 538.050 524.400 ;
        RECT 548.400 522.600 549.600 524.400 ;
        RECT 550.950 524.550 574.050 525.750 ;
        RECT 550.950 524.100 553.050 524.550 ;
        RECT 571.950 524.100 574.050 524.550 ;
        RECT 692.400 526.050 693.600 527.400 ;
        RECT 703.950 527.400 714.600 528.600 ;
        RECT 727.950 528.750 730.050 529.200 ;
        RECT 736.950 528.750 739.050 529.200 ;
        RECT 727.950 528.600 739.050 528.750 ;
        RECT 778.950 528.600 781.050 529.200 ;
        RECT 727.950 527.550 781.050 528.600 ;
        RECT 703.950 526.950 706.050 527.400 ;
        RECT 709.950 527.100 712.050 527.400 ;
        RECT 727.950 527.100 730.050 527.550 ;
        RECT 736.950 527.400 781.050 527.550 ;
        RECT 736.950 527.100 739.050 527.400 ;
        RECT 778.950 527.100 781.050 527.400 ;
        RECT 784.950 528.600 787.050 529.050 ;
        RECT 793.950 528.600 796.050 529.050 ;
        RECT 784.950 527.400 796.050 528.600 ;
        RECT 784.950 526.950 787.050 527.400 ;
        RECT 793.950 526.950 796.050 527.400 ;
        RECT 805.950 528.600 808.050 529.050 ;
        RECT 811.950 528.600 814.050 529.050 ;
        RECT 832.800 528.600 834.900 529.050 ;
        RECT 805.950 527.400 814.050 528.600 ;
        RECT 805.950 526.950 808.050 527.400 ;
        RECT 811.950 526.950 814.050 527.400 ;
        RECT 827.400 527.400 834.900 528.600 ;
        RECT 692.400 524.400 697.050 526.050 ;
        RECT 693.000 523.950 697.050 524.400 ;
        RECT 787.950 525.600 790.050 526.050 ;
        RECT 814.950 525.600 817.050 526.050 ;
        RECT 787.950 524.400 817.050 525.600 ;
        RECT 787.950 523.950 790.050 524.400 ;
        RECT 814.950 523.950 817.050 524.400 ;
        RECT 610.950 522.600 613.050 523.050 ;
        RECT 616.950 522.600 619.050 522.900 ;
        RECT 548.400 521.400 588.600 522.600 ;
        RECT 112.950 519.600 115.050 520.050 ;
        RECT 151.950 519.600 154.050 520.050 ;
        RECT 199.950 519.600 202.050 520.050 ;
        RECT 112.950 518.400 154.050 519.600 ;
        RECT 112.950 517.950 115.050 518.400 ;
        RECT 151.950 517.950 154.050 518.400 ;
        RECT 161.400 518.400 202.050 519.600 ;
        RECT 161.400 517.050 162.600 518.400 ;
        RECT 199.950 517.950 202.050 518.400 ;
        RECT 328.950 519.600 331.050 520.050 ;
        RECT 340.950 519.600 343.050 520.050 ;
        RECT 328.950 518.400 343.050 519.600 ;
        RECT 328.950 517.950 331.050 518.400 ;
        RECT 340.950 517.950 343.050 518.400 ;
        RECT 397.950 519.600 400.050 520.050 ;
        RECT 412.950 519.600 415.050 520.050 ;
        RECT 397.950 518.400 415.050 519.600 ;
        RECT 397.950 517.950 400.050 518.400 ;
        RECT 412.950 517.950 415.050 518.400 ;
        RECT 469.950 517.950 472.050 520.050 ;
        RECT 481.950 519.600 484.050 519.900 ;
        RECT 496.950 519.600 499.050 520.050 ;
        RECT 481.950 518.400 499.050 519.600 ;
        RECT 58.950 516.600 61.050 517.050 ;
        RECT 64.950 516.600 67.050 517.050 ;
        RECT 124.950 516.600 127.050 517.050 ;
        RECT 160.950 516.600 163.050 517.050 ;
        RECT 58.950 515.400 163.050 516.600 ;
        RECT 200.400 516.600 201.600 517.950 ;
        RECT 481.950 517.800 484.050 518.400 ;
        RECT 496.950 517.950 499.050 518.400 ;
        RECT 511.950 519.600 514.050 520.050 ;
        RECT 523.950 519.600 526.050 520.050 ;
        RECT 511.950 518.400 526.050 519.600 ;
        RECT 587.400 519.600 588.600 521.400 ;
        RECT 610.950 521.400 619.050 522.600 ;
        RECT 610.950 520.950 613.050 521.400 ;
        RECT 616.950 520.800 619.050 521.400 ;
        RECT 697.950 522.450 700.050 523.050 ;
        RECT 827.400 522.900 828.600 527.400 ;
        RECT 832.800 526.950 834.900 527.400 ;
        RECT 835.950 528.600 838.050 528.900 ;
        RECT 844.950 528.600 847.050 529.050 ;
        RECT 874.950 528.600 877.050 532.050 ;
        RECT 895.950 531.600 898.050 532.050 ;
        RECT 919.950 531.600 922.050 532.050 ;
        RECT 942.000 531.600 946.050 532.050 ;
        RECT 895.950 530.400 922.050 531.600 ;
        RECT 895.950 529.950 898.050 530.400 ;
        RECT 919.950 529.950 922.050 530.400 ;
        RECT 941.400 529.950 946.050 531.600 ;
        RECT 949.950 531.600 952.050 532.200 ;
        RECT 981.000 531.600 985.050 532.050 ;
        RECT 949.950 531.000 972.600 531.600 ;
        RECT 949.950 530.400 973.050 531.000 ;
        RECT 949.950 530.100 952.050 530.400 ;
        RECT 835.950 527.400 847.050 528.600 ;
        RECT 835.950 526.800 838.050 527.400 ;
        RECT 844.950 526.950 847.050 527.400 ;
        RECT 872.400 528.000 877.050 528.600 ;
        RECT 901.950 528.750 904.050 529.200 ;
        RECT 910.950 528.750 913.050 529.200 ;
        RECT 872.400 527.400 876.600 528.000 ;
        RECT 901.950 527.550 913.050 528.750 ;
        RECT 872.400 525.600 873.600 527.400 ;
        RECT 901.950 527.100 904.050 527.550 ;
        RECT 910.950 527.100 913.050 527.550 ;
        RECT 854.400 524.400 873.600 525.600 ;
        RECT 941.400 525.600 942.600 529.950 ;
        RECT 943.950 528.600 946.050 528.900 ;
        RECT 949.950 528.600 952.050 529.050 ;
        RECT 960.000 528.600 964.050 529.050 ;
        RECT 943.950 527.400 952.050 528.600 ;
        RECT 943.950 526.800 946.050 527.400 ;
        RECT 949.950 526.950 952.050 527.400 ;
        RECT 959.400 526.950 964.050 528.600 ;
        RECT 970.950 526.950 973.050 530.400 ;
        RECT 980.400 529.950 985.050 531.600 ;
        RECT 980.400 529.050 981.600 529.950 ;
        RECT 979.950 526.950 982.050 529.050 ;
        RECT 1000.950 528.600 1003.050 529.050 ;
        RECT 992.400 527.400 1003.050 528.600 ;
        RECT 941.400 524.400 945.600 525.600 ;
        RECT 706.950 522.450 709.050 522.900 ;
        RECT 697.950 521.250 709.050 522.450 ;
        RECT 697.950 520.950 700.050 521.250 ;
        RECT 706.950 520.800 709.050 521.250 ;
        RECT 733.950 522.450 736.050 522.900 ;
        RECT 751.950 522.450 754.050 522.900 ;
        RECT 733.950 521.250 754.050 522.450 ;
        RECT 733.950 520.800 736.050 521.250 ;
        RECT 751.950 520.800 754.050 521.250 ;
        RECT 793.950 522.450 796.050 522.900 ;
        RECT 802.950 522.450 805.050 522.900 ;
        RECT 793.950 521.250 805.050 522.450 ;
        RECT 793.950 520.800 796.050 521.250 ;
        RECT 802.950 520.800 805.050 521.250 ;
        RECT 826.950 520.800 829.050 522.900 ;
        RECT 832.950 522.600 835.050 523.050 ;
        RECT 854.400 522.600 855.600 524.400 ;
        RECT 832.950 521.400 855.600 522.600 ;
        RECT 856.950 522.600 859.050 523.050 ;
        RECT 874.950 522.600 877.050 522.900 ;
        RECT 856.950 521.400 877.050 522.600 ;
        RECT 832.950 520.950 835.050 521.400 ;
        RECT 856.950 520.950 859.050 521.400 ;
        RECT 874.950 520.800 877.050 521.400 ;
        RECT 880.950 522.450 883.050 522.900 ;
        RECT 898.950 522.450 901.050 522.900 ;
        RECT 880.950 521.250 901.050 522.450 ;
        RECT 880.950 520.800 883.050 521.250 ;
        RECT 898.950 520.800 901.050 521.250 ;
        RECT 910.950 522.600 913.050 523.050 ;
        RECT 922.950 522.600 925.050 522.900 ;
        RECT 910.950 521.400 925.050 522.600 ;
        RECT 910.950 520.950 913.050 521.400 ;
        RECT 922.950 520.800 925.050 521.400 ;
        RECT 928.950 522.450 931.050 522.900 ;
        RECT 934.950 522.450 937.050 522.900 ;
        RECT 928.950 521.250 937.050 522.450 ;
        RECT 928.950 520.800 931.050 521.250 ;
        RECT 934.950 520.800 937.050 521.250 ;
        RECT 607.950 519.600 610.050 520.050 ;
        RECT 658.950 519.600 661.050 520.050 ;
        RECT 587.400 518.400 661.050 519.600 ;
        RECT 511.950 517.950 514.050 518.400 ;
        RECT 523.950 517.950 526.050 518.400 ;
        RECT 607.950 517.950 610.050 518.400 ;
        RECT 658.950 517.950 661.050 518.400 ;
        RECT 670.950 519.600 673.050 520.050 ;
        RECT 697.950 519.600 700.050 519.900 ;
        RECT 670.950 518.400 700.050 519.600 ;
        RECT 670.950 517.950 673.050 518.400 ;
        RECT 697.950 517.800 700.050 518.400 ;
        RECT 754.950 519.600 757.050 520.050 ;
        RECT 784.950 519.600 787.050 520.050 ;
        RECT 754.950 518.400 787.050 519.600 ;
        RECT 754.950 517.950 757.050 518.400 ;
        RECT 784.950 517.950 787.050 518.400 ;
        RECT 796.950 519.600 799.050 520.050 ;
        RECT 820.950 519.600 823.050 520.050 ;
        RECT 796.950 518.400 823.050 519.600 ;
        RECT 944.400 519.600 945.600 524.400 ;
        RECT 946.950 522.600 949.050 523.050 ;
        RECT 959.400 522.900 960.600 526.950 ;
        RECT 992.400 523.050 993.600 527.400 ;
        RECT 1000.950 526.950 1003.050 527.400 ;
        RECT 1027.950 526.950 1030.050 529.050 ;
        RECT 1039.800 528.000 1041.900 529.050 ;
        RECT 1039.800 526.950 1042.050 528.000 ;
        RECT 952.950 522.600 955.050 522.900 ;
        RECT 946.950 521.400 955.050 522.600 ;
        RECT 946.950 520.950 949.050 521.400 ;
        RECT 952.950 520.800 955.050 521.400 ;
        RECT 958.950 520.800 961.050 522.900 ;
        RECT 988.950 521.400 993.600 523.050 ;
        RECT 1009.950 522.600 1012.050 522.900 ;
        RECT 1028.400 522.600 1029.600 526.950 ;
        RECT 1039.950 526.050 1042.050 526.950 ;
        RECT 1039.950 525.900 1044.000 526.050 ;
        RECT 1039.950 525.000 1045.050 525.900 ;
        RECT 1040.400 524.400 1045.050 525.000 ;
        RECT 1041.000 523.950 1045.050 524.400 ;
        RECT 1042.950 523.800 1045.050 523.950 ;
        RECT 1033.950 522.600 1036.050 522.900 ;
        RECT 1009.950 521.400 1036.050 522.600 ;
        RECT 988.950 520.950 993.000 521.400 ;
        RECT 1009.950 520.800 1012.050 521.400 ;
        RECT 1033.950 520.800 1036.050 521.400 ;
        RECT 955.950 519.600 958.050 520.050 ;
        RECT 944.400 518.400 958.050 519.600 ;
        RECT 796.950 517.950 799.050 518.400 ;
        RECT 820.950 517.950 823.050 518.400 ;
        RECT 955.950 517.950 958.050 518.400 ;
        RECT 1012.950 519.600 1015.050 520.050 ;
        RECT 1024.950 519.600 1027.050 520.050 ;
        RECT 1012.950 518.400 1027.050 519.600 ;
        RECT 1012.950 517.950 1015.050 518.400 ;
        RECT 1024.950 517.950 1027.050 518.400 ;
        RECT 259.950 516.600 262.050 517.050 ;
        RECT 200.400 515.400 262.050 516.600 ;
        RECT 58.950 514.950 61.050 515.400 ;
        RECT 64.950 514.950 67.050 515.400 ;
        RECT 124.950 514.950 127.050 515.400 ;
        RECT 160.950 514.950 163.050 515.400 ;
        RECT 259.950 514.950 262.050 515.400 ;
        RECT 325.950 516.600 328.050 517.050 ;
        RECT 370.950 516.600 373.050 517.050 ;
        RECT 325.950 515.400 373.050 516.600 ;
        RECT 325.950 514.950 328.050 515.400 ;
        RECT 370.950 514.950 373.050 515.400 ;
        RECT 538.950 516.600 541.050 517.050 ;
        RECT 640.950 516.600 643.050 517.050 ;
        RECT 538.950 515.400 643.050 516.600 ;
        RECT 538.950 514.950 541.050 515.400 ;
        RECT 640.950 514.950 643.050 515.400 ;
        RECT 652.950 516.600 655.050 517.050 ;
        RECT 667.950 516.600 670.050 517.050 ;
        RECT 652.950 515.400 670.050 516.600 ;
        RECT 652.950 514.950 655.050 515.400 ;
        RECT 667.950 514.950 670.050 515.400 ;
        RECT 688.950 516.600 691.050 517.050 ;
        RECT 712.950 516.600 715.050 517.050 ;
        RECT 688.950 515.400 715.050 516.600 ;
        RECT 688.950 514.950 691.050 515.400 ;
        RECT 712.950 514.950 715.050 515.400 ;
        RECT 808.950 516.600 811.050 517.050 ;
        RECT 832.950 516.600 835.050 517.050 ;
        RECT 808.950 515.400 835.050 516.600 ;
        RECT 808.950 514.950 811.050 515.400 ;
        RECT 832.950 514.950 835.050 515.400 ;
        RECT 889.950 516.600 892.050 517.050 ;
        RECT 922.950 516.600 925.050 517.050 ;
        RECT 889.950 515.400 925.050 516.600 ;
        RECT 889.950 514.950 892.050 515.400 ;
        RECT 922.950 514.950 925.050 515.400 ;
        RECT 964.950 516.600 967.050 517.050 ;
        RECT 1003.950 516.600 1006.050 517.050 ;
        RECT 964.950 515.400 1006.050 516.600 ;
        RECT 964.950 514.950 967.050 515.400 ;
        RECT 1003.950 514.950 1006.050 515.400 ;
        RECT 1009.950 516.600 1012.050 517.050 ;
        RECT 1042.950 516.600 1045.050 517.050 ;
        RECT 1009.950 515.400 1045.050 516.600 ;
        RECT 1009.950 514.950 1012.050 515.400 ;
        RECT 1042.950 514.950 1045.050 515.400 ;
        RECT 70.950 513.600 73.050 514.050 ;
        RECT 112.950 513.600 115.050 514.050 ;
        RECT 70.950 512.400 115.050 513.600 ;
        RECT 70.950 511.950 73.050 512.400 ;
        RECT 112.950 511.950 115.050 512.400 ;
        RECT 139.950 513.600 142.050 514.050 ;
        RECT 211.950 513.600 214.050 514.050 ;
        RECT 139.950 512.400 214.050 513.600 ;
        RECT 139.950 511.950 142.050 512.400 ;
        RECT 211.950 511.950 214.050 512.400 ;
        RECT 292.950 513.600 295.050 514.050 ;
        RECT 409.950 513.600 412.050 514.050 ;
        RECT 292.950 512.400 412.050 513.600 ;
        RECT 292.950 511.950 295.050 512.400 ;
        RECT 409.950 511.950 412.050 512.400 ;
        RECT 448.950 513.600 451.050 514.050 ;
        RECT 490.950 513.600 493.050 514.050 ;
        RECT 448.950 512.400 493.050 513.600 ;
        RECT 448.950 511.950 451.050 512.400 ;
        RECT 490.950 511.950 493.050 512.400 ;
        RECT 529.950 513.600 532.050 514.050 ;
        RECT 610.800 513.600 612.900 514.050 ;
        RECT 529.950 512.400 612.900 513.600 ;
        RECT 529.950 511.950 532.050 512.400 ;
        RECT 610.800 511.950 612.900 512.400 ;
        RECT 613.950 513.600 616.050 514.050 ;
        RECT 622.950 513.600 625.050 514.050 ;
        RECT 613.950 512.400 625.050 513.600 ;
        RECT 613.950 511.950 616.050 512.400 ;
        RECT 622.950 511.950 625.050 512.400 ;
        RECT 643.950 513.600 646.050 514.050 ;
        RECT 682.950 513.600 685.050 514.050 ;
        RECT 709.950 513.600 712.050 514.050 ;
        RECT 643.950 512.400 685.050 513.600 ;
        RECT 643.950 511.950 646.050 512.400 ;
        RECT 682.950 511.950 685.050 512.400 ;
        RECT 686.400 512.400 712.050 513.600 ;
        RECT 148.950 510.600 151.050 511.050 ;
        RECT 184.950 510.600 187.050 511.050 ;
        RECT 148.950 509.400 187.050 510.600 ;
        RECT 148.950 508.950 151.050 509.400 ;
        RECT 184.950 508.950 187.050 509.400 ;
        RECT 220.950 510.600 223.050 511.050 ;
        RECT 232.950 510.600 235.050 511.050 ;
        RECT 271.950 510.600 274.050 511.050 ;
        RECT 220.950 509.400 274.050 510.600 ;
        RECT 220.950 508.950 223.050 509.400 ;
        RECT 232.950 508.950 235.050 509.400 ;
        RECT 271.950 508.950 274.050 509.400 ;
        RECT 319.950 510.600 322.050 511.050 ;
        RECT 331.950 510.600 334.050 511.050 ;
        RECT 346.950 510.600 349.050 511.050 ;
        RECT 319.950 509.400 349.050 510.600 ;
        RECT 319.950 508.950 322.050 509.400 ;
        RECT 331.950 508.950 334.050 509.400 ;
        RECT 346.950 508.950 349.050 509.400 ;
        RECT 502.950 510.600 505.050 511.050 ;
        RECT 514.950 510.600 517.050 511.050 ;
        RECT 502.950 509.400 517.050 510.600 ;
        RECT 502.950 508.950 505.050 509.400 ;
        RECT 514.950 508.950 517.050 509.400 ;
        RECT 637.950 510.600 640.050 511.050 ;
        RECT 686.400 510.600 687.600 512.400 ;
        RECT 709.950 511.950 712.050 512.400 ;
        RECT 784.950 513.600 787.050 514.050 ;
        RECT 799.950 513.600 802.050 514.050 ;
        RECT 784.950 512.400 802.050 513.600 ;
        RECT 784.950 511.950 787.050 512.400 ;
        RECT 799.950 511.950 802.050 512.400 ;
        RECT 841.950 513.600 844.050 514.050 ;
        RECT 850.950 513.600 853.050 514.050 ;
        RECT 841.950 512.400 853.050 513.600 ;
        RECT 841.950 511.950 844.050 512.400 ;
        RECT 850.950 511.950 853.050 512.400 ;
        RECT 913.950 513.600 916.050 514.050 ;
        RECT 931.950 513.600 934.050 514.050 ;
        RECT 913.950 512.400 934.050 513.600 ;
        RECT 913.950 511.950 916.050 512.400 ;
        RECT 931.950 511.950 934.050 512.400 ;
        RECT 943.950 513.600 946.050 514.050 ;
        RECT 976.950 513.600 979.050 514.050 ;
        RECT 943.950 512.400 979.050 513.600 ;
        RECT 943.950 511.950 946.050 512.400 ;
        RECT 976.950 511.950 979.050 512.400 ;
        RECT 997.950 513.600 1000.050 514.050 ;
        RECT 1015.950 513.600 1018.050 514.050 ;
        RECT 997.950 512.400 1018.050 513.600 ;
        RECT 997.950 511.950 1000.050 512.400 ;
        RECT 1015.950 511.950 1018.050 512.400 ;
        RECT 721.950 510.600 724.050 511.050 ;
        RECT 745.950 510.600 748.050 511.050 ;
        RECT 637.950 509.400 687.600 510.600 ;
        RECT 689.400 509.400 748.050 510.600 ;
        RECT 637.950 508.950 640.050 509.400 ;
        RECT 61.950 507.600 64.050 508.050 ;
        RECT 97.950 507.600 100.050 508.050 ;
        RECT 61.950 506.400 100.050 507.600 ;
        RECT 61.950 505.950 64.050 506.400 ;
        RECT 97.950 505.950 100.050 506.400 ;
        RECT 427.950 507.600 430.050 508.050 ;
        RECT 457.950 507.600 460.050 508.050 ;
        RECT 427.950 506.400 460.050 507.600 ;
        RECT 427.950 505.950 430.050 506.400 ;
        RECT 457.950 505.950 460.050 506.400 ;
        RECT 586.950 507.600 589.050 508.050 ;
        RECT 598.950 507.600 601.050 508.050 ;
        RECT 586.950 506.400 601.050 507.600 ;
        RECT 586.950 505.950 589.050 506.400 ;
        RECT 598.950 505.950 601.050 506.400 ;
        RECT 652.950 507.600 655.050 508.050 ;
        RECT 670.950 507.600 673.050 508.050 ;
        RECT 652.950 506.400 673.050 507.600 ;
        RECT 652.950 505.950 655.050 506.400 ;
        RECT 670.950 505.950 673.050 506.400 ;
        RECT 676.950 507.600 679.050 508.050 ;
        RECT 689.400 507.600 690.600 509.400 ;
        RECT 721.950 508.950 724.050 509.400 ;
        RECT 745.950 508.950 748.050 509.400 ;
        RECT 790.950 510.600 793.050 511.050 ;
        RECT 808.950 510.600 811.050 511.050 ;
        RECT 790.950 509.400 811.050 510.600 ;
        RECT 790.950 508.950 793.050 509.400 ;
        RECT 808.950 508.950 811.050 509.400 ;
        RECT 841.950 510.600 844.050 510.900 ;
        RECT 865.950 510.600 868.050 511.050 ;
        RECT 841.950 509.400 868.050 510.600 ;
        RECT 841.950 508.800 844.050 509.400 ;
        RECT 865.950 508.950 868.050 509.400 ;
        RECT 958.950 510.600 961.050 511.050 ;
        RECT 988.950 510.600 991.050 511.050 ;
        RECT 958.950 509.400 991.050 510.600 ;
        RECT 958.950 508.950 961.050 509.400 ;
        RECT 988.950 508.950 991.050 509.400 ;
        RECT 676.950 506.400 690.600 507.600 ;
        RECT 694.950 507.600 697.050 508.050 ;
        RECT 718.950 507.600 721.050 508.050 ;
        RECT 823.950 507.600 826.050 508.050 ;
        RECT 862.950 507.600 865.050 508.050 ;
        RECT 694.950 506.400 721.050 507.600 ;
        RECT 676.950 505.950 679.050 506.400 ;
        RECT 694.950 505.950 697.050 506.400 ;
        RECT 718.950 505.950 721.050 506.400 ;
        RECT 725.400 506.400 744.600 507.600 ;
        RECT 196.950 504.600 199.050 505.050 ;
        RECT 202.950 504.600 205.050 505.050 ;
        RECT 196.950 503.400 205.050 504.600 ;
        RECT 196.950 502.950 199.050 503.400 ;
        RECT 202.950 502.950 205.050 503.400 ;
        RECT 229.950 504.600 232.050 505.050 ;
        RECT 265.950 504.600 268.050 505.050 ;
        RECT 229.950 503.400 268.050 504.600 ;
        RECT 229.950 502.950 232.050 503.400 ;
        RECT 265.950 502.950 268.050 503.400 ;
        RECT 715.950 504.600 718.050 505.050 ;
        RECT 725.400 504.600 726.600 506.400 ;
        RECT 715.950 503.400 726.600 504.600 ;
        RECT 743.400 504.600 744.600 506.400 ;
        RECT 823.950 506.400 865.050 507.600 ;
        RECT 823.950 505.950 826.050 506.400 ;
        RECT 862.950 505.950 865.050 506.400 ;
        RECT 904.950 507.600 907.050 508.050 ;
        RECT 913.950 507.600 916.050 508.050 ;
        RECT 904.950 506.400 916.050 507.600 ;
        RECT 904.950 505.950 907.050 506.400 ;
        RECT 913.950 505.950 916.050 506.400 ;
        RECT 943.950 507.600 946.050 508.050 ;
        RECT 973.950 507.600 976.050 508.050 ;
        RECT 943.950 506.400 976.050 507.600 ;
        RECT 943.950 505.950 946.050 506.400 ;
        RECT 973.950 505.950 976.050 506.400 ;
        RECT 1000.950 507.600 1003.050 508.050 ;
        RECT 1015.950 507.600 1018.050 508.050 ;
        RECT 1000.950 506.400 1018.050 507.600 ;
        RECT 1000.950 505.950 1003.050 506.400 ;
        RECT 1015.950 505.950 1018.050 506.400 ;
        RECT 1021.950 507.600 1024.050 508.050 ;
        RECT 1030.950 507.600 1033.050 508.050 ;
        RECT 1021.950 506.400 1033.050 507.600 ;
        RECT 1021.950 505.950 1024.050 506.400 ;
        RECT 1030.950 505.950 1033.050 506.400 ;
        RECT 811.950 504.600 814.050 505.050 ;
        RECT 743.400 503.400 814.050 504.600 ;
        RECT 715.950 502.950 718.050 503.400 ;
        RECT 811.950 502.950 814.050 503.400 ;
        RECT 838.950 504.600 841.050 505.050 ;
        RECT 850.950 504.600 853.050 505.050 ;
        RECT 838.950 503.400 853.050 504.600 ;
        RECT 838.950 502.950 841.050 503.400 ;
        RECT 850.950 502.950 853.050 503.400 ;
        RECT 55.950 501.600 58.050 502.050 ;
        RECT 70.950 501.600 73.050 502.050 ;
        RECT 55.950 500.400 73.050 501.600 ;
        RECT 55.950 499.950 58.050 500.400 ;
        RECT 70.950 499.950 73.050 500.400 ;
        RECT 178.950 501.600 181.050 502.050 ;
        RECT 334.950 501.600 337.050 502.050 ;
        RECT 340.950 501.600 343.050 502.050 ;
        RECT 358.950 501.600 361.050 502.050 ;
        RECT 178.950 500.400 189.600 501.600 ;
        RECT 178.950 499.950 181.050 500.400 ;
        RECT 175.950 498.600 178.050 499.050 ;
        RECT 175.950 497.400 183.600 498.600 ;
        RECT 175.950 496.950 178.050 497.400 ;
        RECT 16.950 495.750 19.050 496.200 ;
        RECT 25.950 495.750 28.050 496.200 ;
        RECT 16.950 494.550 28.050 495.750 ;
        RECT 16.950 494.100 19.050 494.550 ;
        RECT 25.950 494.100 28.050 494.550 ;
        RECT 40.950 495.600 43.050 496.200 ;
        RECT 82.950 495.600 85.050 496.200 ;
        RECT 40.950 494.400 85.050 495.600 ;
        RECT 40.950 494.100 43.050 494.400 ;
        RECT 82.950 494.100 85.050 494.400 ;
        RECT 88.950 495.600 91.050 496.200 ;
        RECT 109.950 495.600 112.050 496.200 ;
        RECT 88.950 494.400 112.050 495.600 ;
        RECT 88.950 494.100 91.050 494.400 ;
        RECT 109.950 494.100 112.050 494.400 ;
        RECT 115.950 495.750 118.050 496.200 ;
        RECT 124.950 495.750 127.050 496.200 ;
        RECT 115.950 494.550 127.050 495.750 ;
        RECT 115.950 494.100 118.050 494.550 ;
        RECT 124.950 494.100 127.050 494.550 ;
        RECT 139.950 495.600 142.050 496.200 ;
        RECT 182.400 496.050 183.600 497.400 ;
        RECT 148.950 495.600 151.050 496.050 ;
        RECT 139.950 494.400 151.050 495.600 ;
        RECT 182.400 494.400 187.050 496.050 ;
        RECT 139.950 494.100 142.050 494.400 ;
        RECT 148.950 493.950 151.050 494.400 ;
        RECT 183.000 493.950 187.050 494.400 ;
        RECT 188.400 493.050 189.600 500.400 ;
        RECT 334.950 500.400 361.050 501.600 ;
        RECT 334.950 499.950 337.050 500.400 ;
        RECT 340.950 499.950 343.050 500.400 ;
        RECT 358.950 499.950 361.050 500.400 ;
        RECT 379.950 501.600 382.050 502.050 ;
        RECT 397.950 501.600 400.050 502.050 ;
        RECT 379.950 500.400 400.050 501.600 ;
        RECT 379.950 499.950 382.050 500.400 ;
        RECT 397.950 499.950 400.050 500.400 ;
        RECT 454.950 501.600 457.050 502.050 ;
        RECT 487.950 501.600 490.050 502.050 ;
        RECT 454.950 500.400 490.050 501.600 ;
        RECT 454.950 499.950 457.050 500.400 ;
        RECT 487.950 499.950 490.050 500.400 ;
        RECT 496.950 501.600 499.050 502.050 ;
        RECT 514.950 501.600 517.050 502.050 ;
        RECT 496.950 500.400 517.050 501.600 ;
        RECT 496.950 499.950 499.050 500.400 ;
        RECT 514.950 499.950 517.050 500.400 ;
        RECT 526.950 501.600 529.050 502.050 ;
        RECT 544.950 501.600 547.050 502.050 ;
        RECT 526.950 500.400 547.050 501.600 ;
        RECT 526.950 499.950 529.050 500.400 ;
        RECT 544.950 499.950 547.050 500.400 ;
        RECT 550.950 501.600 553.050 502.050 ;
        RECT 631.950 501.600 634.050 502.050 ;
        RECT 550.950 500.400 634.050 501.600 ;
        RECT 550.950 499.950 553.050 500.400 ;
        RECT 631.950 499.950 634.050 500.400 ;
        RECT 829.950 501.600 832.050 502.050 ;
        RECT 835.950 501.600 838.050 502.050 ;
        RECT 829.950 500.400 838.050 501.600 ;
        RECT 829.950 499.950 832.050 500.400 ;
        RECT 835.950 499.950 838.050 500.400 ;
        RECT 916.950 501.600 919.050 502.050 ;
        RECT 964.950 501.600 967.050 502.050 ;
        RECT 916.950 500.400 967.050 501.600 ;
        RECT 916.950 499.950 919.050 500.400 ;
        RECT 964.950 499.950 967.050 500.400 ;
        RECT 970.950 501.600 973.050 502.050 ;
        RECT 982.950 501.600 985.050 501.900 ;
        RECT 970.950 500.400 985.050 501.600 ;
        RECT 970.950 499.950 973.050 500.400 ;
        RECT 982.950 499.800 985.050 500.400 ;
        RECT 241.950 498.600 244.050 499.050 ;
        RECT 227.400 497.400 244.050 498.600 ;
        RECT 196.950 495.600 199.050 496.050 ;
        RECT 205.950 495.600 208.050 496.050 ;
        RECT 220.950 495.600 223.050 496.200 ;
        RECT 196.950 494.400 223.050 495.600 ;
        RECT 196.950 493.950 199.050 494.400 ;
        RECT 205.950 493.950 208.050 494.400 ;
        RECT 220.950 494.100 223.050 494.400 ;
        RECT 188.400 491.400 193.050 493.050 ;
        RECT 189.000 490.950 193.050 491.400 ;
        RECT 227.400 490.050 228.600 497.400 ;
        RECT 241.950 496.950 244.050 497.400 ;
        RECT 253.950 498.600 256.050 498.900 ;
        RECT 277.950 498.600 280.050 499.050 ;
        RECT 253.950 497.400 280.050 498.600 ;
        RECT 253.950 496.800 256.050 497.400 ;
        RECT 277.950 496.950 280.050 497.400 ;
        RECT 295.950 498.600 298.050 499.050 ;
        RECT 304.950 498.600 307.050 499.050 ;
        RECT 295.950 497.400 307.050 498.600 ;
        RECT 295.950 496.950 298.050 497.400 ;
        RECT 304.950 496.950 307.050 497.400 ;
        RECT 604.950 498.600 607.050 499.050 ;
        RECT 616.950 498.600 619.050 499.050 ;
        RECT 763.950 498.600 766.050 499.050 ;
        RECT 604.950 497.400 619.050 498.600 ;
        RECT 604.950 496.950 607.050 497.400 ;
        RECT 616.950 496.950 619.050 497.400 ;
        RECT 743.400 497.400 766.050 498.600 ;
        RECT 235.950 495.750 238.050 496.200 ;
        RECT 244.950 495.750 247.050 496.200 ;
        RECT 235.950 494.550 247.050 495.750 ;
        RECT 235.950 494.100 238.050 494.550 ;
        RECT 244.950 494.100 247.050 494.550 ;
        RECT 265.950 494.100 268.050 496.200 ;
        RECT 289.950 495.600 292.050 496.200 ;
        RECT 307.950 495.600 310.050 496.050 ;
        RECT 289.950 494.400 310.050 495.600 ;
        RECT 289.950 494.100 292.050 494.400 ;
        RECT 266.400 492.600 267.600 494.100 ;
        RECT 307.950 493.950 310.050 494.400 ;
        RECT 346.950 495.600 349.050 496.200 ;
        RECT 355.950 495.600 358.050 496.050 ;
        RECT 346.950 494.400 358.050 495.600 ;
        RECT 346.950 494.100 349.050 494.400 ;
        RECT 355.950 493.950 358.050 494.400 ;
        RECT 367.950 495.750 370.050 496.200 ;
        RECT 385.950 495.750 388.050 496.200 ;
        RECT 367.950 494.550 388.050 495.750 ;
        RECT 367.950 494.100 370.050 494.550 ;
        RECT 385.950 494.100 388.050 494.550 ;
        RECT 409.950 495.750 412.050 496.200 ;
        RECT 415.950 495.750 418.050 496.200 ;
        RECT 409.950 494.550 418.050 495.750 ;
        RECT 409.950 494.100 412.050 494.550 ;
        RECT 415.950 494.100 418.050 494.550 ;
        RECT 421.950 495.750 424.050 496.200 ;
        RECT 436.950 495.750 439.050 496.200 ;
        RECT 421.950 494.550 439.050 495.750 ;
        RECT 421.950 494.100 424.050 494.550 ;
        RECT 436.950 494.100 439.050 494.550 ;
        RECT 442.950 495.600 445.050 496.200 ;
        RECT 457.950 495.600 460.050 496.050 ;
        RECT 442.950 494.400 460.050 495.600 ;
        RECT 442.950 494.100 445.050 494.400 ;
        RECT 457.950 493.950 460.050 494.400 ;
        RECT 472.950 494.100 475.050 496.200 ;
        RECT 502.950 495.600 505.050 496.200 ;
        RECT 520.950 495.600 523.050 496.200 ;
        RECT 743.400 496.050 744.600 497.400 ;
        RECT 763.950 496.950 766.050 497.400 ;
        RECT 811.950 498.600 814.050 499.050 ;
        RECT 820.950 498.600 823.050 499.050 ;
        RECT 811.950 497.400 823.050 498.600 ;
        RECT 811.950 496.950 814.050 497.400 ;
        RECT 820.950 496.950 823.050 497.400 ;
        RECT 919.950 498.600 922.050 499.050 ;
        RECT 934.950 498.600 937.050 499.050 ;
        RECT 919.950 497.400 937.050 498.600 ;
        RECT 919.950 496.950 922.050 497.400 ;
        RECT 934.950 496.950 937.050 497.400 ;
        RECT 985.950 498.600 988.050 499.050 ;
        RECT 994.950 498.600 997.050 499.050 ;
        RECT 985.950 497.400 997.050 498.600 ;
        RECT 985.950 496.950 988.050 497.400 ;
        RECT 994.950 496.950 997.050 497.400 ;
        RECT 502.950 494.400 523.050 495.600 ;
        RECT 502.950 494.100 505.050 494.400 ;
        RECT 520.950 494.100 523.050 494.400 ;
        RECT 544.950 495.600 547.050 496.050 ;
        RECT 556.950 495.600 559.050 496.050 ;
        RECT 544.950 494.400 559.050 495.600 ;
        RECT 263.400 492.000 267.600 492.600 ;
        RECT 262.950 491.400 267.600 492.000 ;
        RECT 473.400 492.600 474.600 494.100 ;
        RECT 544.950 493.950 547.050 494.400 ;
        RECT 556.950 493.950 559.050 494.400 ;
        RECT 643.950 495.600 648.000 496.050 ;
        RECT 730.950 495.600 733.050 496.050 ;
        RECT 643.950 493.950 648.600 495.600 ;
        RECT 665.400 495.000 733.050 495.600 ;
        RECT 484.950 492.600 487.050 493.050 ;
        RECT 473.400 491.400 487.050 492.600 ;
        RECT 85.950 489.450 88.050 489.900 ;
        RECT 97.950 489.450 100.050 489.900 ;
        RECT 85.950 488.250 100.050 489.450 ;
        RECT 85.950 487.800 88.050 488.250 ;
        RECT 97.950 487.800 100.050 488.250 ;
        RECT 124.950 489.600 127.050 490.050 ;
        RECT 136.950 489.600 139.050 489.900 ;
        RECT 124.950 488.400 139.050 489.600 ;
        RECT 124.950 487.950 127.050 488.400 ;
        RECT 136.950 487.800 139.050 488.400 ;
        RECT 142.950 489.600 145.050 489.900 ;
        RECT 160.950 489.600 163.050 489.900 ;
        RECT 142.950 488.400 163.050 489.600 ;
        RECT 142.950 487.800 145.050 488.400 ;
        RECT 160.950 487.800 163.050 488.400 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 241.950 489.450 244.050 489.900 ;
        RECT 253.950 489.450 256.050 489.900 ;
        RECT 241.950 488.250 256.050 489.450 ;
        RECT 241.950 487.800 244.050 488.250 ;
        RECT 253.950 487.800 256.050 488.250 ;
        RECT 262.950 487.950 265.050 491.400 ;
        RECT 484.950 490.950 487.050 491.400 ;
        RECT 580.950 492.600 583.050 493.050 ;
        RECT 598.950 492.600 601.050 493.050 ;
        RECT 580.950 491.400 601.050 492.600 ;
        RECT 580.950 490.950 583.050 491.400 ;
        RECT 598.950 490.950 601.050 491.400 ;
        RECT 268.950 489.600 271.050 489.900 ;
        RECT 268.950 488.400 324.600 489.600 ;
        RECT 268.950 487.800 271.050 488.400 ;
        RECT 19.950 486.600 22.050 487.050 ;
        RECT 49.950 486.600 52.050 487.050 ;
        RECT 58.950 486.600 61.050 487.050 ;
        RECT 19.950 485.400 61.050 486.600 ;
        RECT 19.950 484.950 22.050 485.400 ;
        RECT 49.950 484.950 52.050 485.400 ;
        RECT 58.950 484.950 61.050 485.400 ;
        RECT 91.950 486.600 94.050 487.050 ;
        RECT 103.950 486.600 106.050 487.050 ;
        RECT 115.950 486.600 118.050 487.050 ;
        RECT 91.950 485.400 118.050 486.600 ;
        RECT 91.950 484.950 94.050 485.400 ;
        RECT 103.950 484.950 106.050 485.400 ;
        RECT 115.950 484.950 118.050 485.400 ;
        RECT 121.950 486.600 124.050 487.050 ;
        RECT 142.950 486.600 145.050 487.050 ;
        RECT 121.950 485.400 145.050 486.600 ;
        RECT 323.400 486.600 324.600 488.400 ;
        RECT 355.950 489.450 358.050 489.900 ;
        RECT 364.950 489.450 367.050 489.900 ;
        RECT 355.950 488.250 367.050 489.450 ;
        RECT 355.950 487.800 358.050 488.250 ;
        RECT 364.950 487.800 367.050 488.250 ;
        RECT 418.950 489.600 421.050 489.900 ;
        RECT 439.950 489.600 442.050 489.900 ;
        RECT 418.950 488.400 442.050 489.600 ;
        RECT 418.950 487.800 421.050 488.400 ;
        RECT 439.950 487.800 442.050 488.400 ;
        RECT 457.950 489.450 460.050 489.900 ;
        RECT 469.950 489.450 472.050 489.900 ;
        RECT 457.950 488.250 472.050 489.450 ;
        RECT 457.950 487.800 460.050 488.250 ;
        RECT 469.950 487.800 472.050 488.250 ;
        RECT 487.950 489.450 490.050 489.900 ;
        RECT 493.950 489.450 496.050 489.900 ;
        RECT 487.950 488.250 496.050 489.450 ;
        RECT 487.950 487.800 490.050 488.250 ;
        RECT 493.950 487.800 496.050 488.250 ;
        RECT 535.950 487.800 538.050 489.900 ;
        RECT 556.950 489.600 559.050 490.050 ;
        RECT 577.950 489.600 580.050 490.050 ;
        RECT 556.950 488.400 580.050 489.600 ;
        RECT 556.950 487.950 559.050 488.400 ;
        RECT 577.950 487.950 580.050 488.400 ;
        RECT 325.950 486.600 328.050 487.050 ;
        RECT 343.950 486.600 346.050 487.050 ;
        RECT 323.400 485.400 346.050 486.600 ;
        RECT 121.950 484.950 124.050 485.400 ;
        RECT 142.950 484.950 145.050 485.400 ;
        RECT 325.950 484.950 328.050 485.400 ;
        RECT 343.950 484.950 346.050 485.400 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 409.950 486.600 412.050 487.050 ;
        RECT 370.950 485.400 412.050 486.600 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 409.950 484.950 412.050 485.400 ;
        RECT 478.950 486.600 481.050 487.050 ;
        RECT 499.950 486.600 502.050 487.050 ;
        RECT 478.950 485.400 502.050 486.600 ;
        RECT 536.400 486.600 537.600 487.800 ;
        RECT 647.400 487.050 648.600 493.950 ;
        RECT 664.950 494.400 733.050 495.000 ;
        RECT 664.950 490.950 667.050 494.400 ;
        RECT 730.950 493.950 733.050 494.400 ;
        RECT 739.950 494.400 744.600 496.050 ;
        RECT 814.950 495.600 817.050 496.050 ;
        RECT 826.950 495.600 829.050 496.050 ;
        RECT 814.950 494.400 829.050 495.600 ;
        RECT 739.950 493.950 744.000 494.400 ;
        RECT 814.950 493.950 817.050 494.400 ;
        RECT 826.950 493.950 829.050 494.400 ;
        RECT 841.950 493.950 844.050 496.050 ;
        RECT 862.950 495.750 865.050 496.200 ;
        RECT 913.950 495.750 916.050 496.050 ;
        RECT 862.950 494.550 916.050 495.750 ;
        RECT 862.950 494.100 865.050 494.550 ;
        RECT 913.950 493.950 916.050 494.550 ;
        RECT 937.950 495.600 940.050 496.050 ;
        RECT 952.950 495.600 955.050 496.200 ;
        RECT 990.000 495.600 994.050 496.050 ;
        RECT 937.950 494.400 955.050 495.600 ;
        RECT 937.950 493.950 940.050 494.400 ;
        RECT 952.950 494.100 955.050 494.400 ;
        RECT 989.400 493.950 994.050 495.600 ;
        RECT 1003.950 495.600 1006.050 496.200 ;
        RECT 1021.950 495.600 1024.050 496.200 ;
        RECT 1003.950 494.400 1024.050 495.600 ;
        RECT 1003.950 494.100 1006.050 494.400 ;
        RECT 1021.950 494.100 1024.050 494.400 ;
        RECT 1027.950 495.600 1030.050 496.050 ;
        RECT 1036.950 495.600 1039.050 496.050 ;
        RECT 1027.950 494.400 1039.050 495.600 ;
        RECT 1027.950 493.950 1030.050 494.400 ;
        RECT 1036.950 493.950 1039.050 494.400 ;
        RECT 757.950 489.600 760.050 493.050 ;
        RECT 763.950 492.450 766.050 492.900 ;
        RECT 778.950 492.450 781.050 492.900 ;
        RECT 763.950 491.250 781.050 492.450 ;
        RECT 763.950 490.800 766.050 491.250 ;
        RECT 778.950 490.800 781.050 491.250 ;
        RECT 805.950 492.750 808.050 493.200 ;
        RECT 817.950 492.750 820.050 492.900 ;
        RECT 805.950 491.550 820.050 492.750 ;
        RECT 805.950 491.100 808.050 491.550 ;
        RECT 817.950 490.800 820.050 491.550 ;
        RECT 842.400 490.050 843.600 493.950 ;
        RECT 913.950 492.600 916.050 492.900 ;
        RECT 919.950 492.600 922.050 493.200 ;
        RECT 890.400 491.400 922.050 492.600 ;
        RECT 757.950 489.000 762.600 489.600 ;
        RECT 758.400 488.400 762.600 489.000 ;
        RECT 761.400 487.050 762.600 488.400 ;
        RECT 841.950 487.950 844.050 490.050 ;
        RECT 853.950 489.600 856.050 490.050 ;
        RECT 890.400 489.600 891.600 491.400 ;
        RECT 913.950 490.800 916.050 491.400 ;
        RECT 919.950 491.100 922.050 491.400 ;
        RECT 925.950 490.950 928.050 493.050 ;
        RECT 934.950 492.600 937.050 493.050 ;
        RECT 964.950 492.600 967.050 493.050 ;
        RECT 989.400 492.600 990.600 493.950 ;
        RECT 934.950 492.000 948.600 492.600 ;
        RECT 934.950 491.400 949.050 492.000 ;
        RECT 934.950 490.950 937.050 491.400 ;
        RECT 853.950 488.400 891.600 489.600 ;
        RECT 853.950 487.950 856.050 488.400 ;
        RECT 926.400 487.050 927.600 490.950 ;
        RECT 946.950 487.950 949.050 491.400 ;
        RECT 964.950 491.400 990.600 492.600 ;
        RECT 964.950 490.950 967.050 491.400 ;
        RECT 989.400 490.050 990.600 491.400 ;
        RECT 989.400 488.400 994.050 490.050 ;
        RECT 990.000 487.950 994.050 488.400 ;
        RECT 1000.950 489.450 1003.050 489.900 ;
        RECT 1009.950 489.450 1012.050 489.900 ;
        RECT 1000.950 488.250 1012.050 489.450 ;
        RECT 1000.950 487.800 1003.050 488.250 ;
        RECT 1009.950 487.800 1012.050 488.250 ;
        RECT 544.950 486.600 547.050 487.050 ;
        RECT 536.400 485.400 547.050 486.600 ;
        RECT 478.950 484.950 481.050 485.400 ;
        RECT 499.950 484.950 502.050 485.400 ;
        RECT 544.950 484.950 547.050 485.400 ;
        RECT 646.950 484.950 649.050 487.050 ;
        RECT 688.950 486.600 691.050 487.050 ;
        RECT 727.950 486.600 730.050 487.050 ;
        RECT 757.950 486.600 760.050 487.050 ;
        RECT 688.950 485.400 760.050 486.600 ;
        RECT 761.400 485.400 766.050 487.050 ;
        RECT 688.950 484.950 691.050 485.400 ;
        RECT 727.950 484.950 730.050 485.400 ;
        RECT 757.950 484.950 760.050 485.400 ;
        RECT 762.000 484.950 766.050 485.400 ;
        RECT 799.950 486.600 802.050 487.050 ;
        RECT 856.950 486.600 859.050 487.050 ;
        RECT 799.950 485.400 843.600 486.600 ;
        RECT 799.950 484.950 802.050 485.400 ;
        RECT 259.950 483.600 262.050 484.050 ;
        RECT 292.950 483.600 295.050 484.050 ;
        RECT 259.950 482.400 295.050 483.600 ;
        RECT 259.950 481.950 262.050 482.400 ;
        RECT 292.950 481.950 295.050 482.400 ;
        RECT 310.950 483.600 313.050 484.050 ;
        RECT 316.950 483.600 319.050 484.050 ;
        RECT 322.950 483.600 325.050 484.050 ;
        RECT 310.950 482.400 325.050 483.600 ;
        RECT 310.950 481.950 313.050 482.400 ;
        RECT 316.950 481.950 319.050 482.400 ;
        RECT 322.950 481.950 325.050 482.400 ;
        RECT 508.950 483.600 511.050 484.050 ;
        RECT 541.950 483.600 544.050 484.050 ;
        RECT 508.950 482.400 544.050 483.600 ;
        RECT 508.950 481.950 511.050 482.400 ;
        RECT 541.950 481.950 544.050 482.400 ;
        RECT 649.950 483.600 652.050 484.050 ;
        RECT 664.950 483.600 667.050 484.050 ;
        RECT 778.950 483.600 781.050 484.050 ;
        RECT 649.950 482.400 667.050 483.600 ;
        RECT 649.950 481.950 652.050 482.400 ;
        RECT 664.950 481.950 667.050 482.400 ;
        RECT 731.400 482.400 781.050 483.600 ;
        RECT 25.950 480.600 28.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 25.950 479.400 121.050 480.600 ;
        RECT 25.950 478.950 28.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 157.950 480.600 160.050 481.050 ;
        RECT 175.950 480.600 178.050 481.050 ;
        RECT 157.950 479.400 178.050 480.600 ;
        RECT 157.950 478.950 160.050 479.400 ;
        RECT 175.950 478.950 178.050 479.400 ;
        RECT 247.950 480.600 250.050 481.050 ;
        RECT 268.950 480.600 271.050 481.050 ;
        RECT 247.950 479.400 271.050 480.600 ;
        RECT 247.950 478.950 250.050 479.400 ;
        RECT 268.950 478.950 271.050 479.400 ;
        RECT 280.950 480.600 283.050 481.050 ;
        RECT 292.950 480.600 295.050 480.900 ;
        RECT 280.950 479.400 295.050 480.600 ;
        RECT 280.950 478.950 283.050 479.400 ;
        RECT 292.950 478.800 295.050 479.400 ;
        RECT 403.950 480.600 406.050 481.050 ;
        RECT 502.950 480.600 505.050 481.050 ;
        RECT 403.950 479.400 505.050 480.600 ;
        RECT 403.950 478.950 406.050 479.400 ;
        RECT 502.950 478.950 505.050 479.400 ;
        RECT 514.950 480.600 517.050 481.050 ;
        RECT 619.950 480.600 622.050 481.050 ;
        RECT 514.950 479.400 622.050 480.600 ;
        RECT 514.950 478.950 517.050 479.400 ;
        RECT 619.950 478.950 622.050 479.400 ;
        RECT 277.950 477.600 280.050 478.050 ;
        RECT 298.950 477.600 301.050 478.050 ;
        RECT 337.950 477.600 340.050 478.050 ;
        RECT 460.950 477.600 463.050 478.050 ;
        RECT 277.950 476.400 340.050 477.600 ;
        RECT 277.950 475.950 280.050 476.400 ;
        RECT 298.950 475.950 301.050 476.400 ;
        RECT 337.950 475.950 340.050 476.400 ;
        RECT 434.400 476.400 463.050 477.600 ;
        RECT 190.950 474.600 193.050 475.050 ;
        RECT 199.950 474.600 202.050 475.050 ;
        RECT 190.950 473.400 202.050 474.600 ;
        RECT 190.950 472.950 193.050 473.400 ;
        RECT 199.950 472.950 202.050 473.400 ;
        RECT 211.950 474.600 214.050 475.050 ;
        RECT 434.400 474.600 435.600 476.400 ;
        RECT 460.950 475.950 463.050 476.400 ;
        RECT 670.950 477.600 673.050 478.050 ;
        RECT 731.400 477.600 732.600 482.400 ;
        RECT 778.950 481.950 781.050 482.400 ;
        RECT 799.950 483.600 802.050 483.900 ;
        RECT 808.800 483.600 810.900 484.050 ;
        RECT 799.950 482.400 810.900 483.600 ;
        RECT 799.950 481.800 802.050 482.400 ;
        RECT 808.800 481.950 810.900 482.400 ;
        RECT 811.950 483.600 814.050 484.050 ;
        RECT 832.950 483.600 835.050 484.050 ;
        RECT 838.950 483.600 841.050 484.050 ;
        RECT 811.950 482.400 841.050 483.600 ;
        RECT 842.400 483.600 843.600 485.400 ;
        RECT 856.950 485.400 882.600 486.600 ;
        RECT 856.950 484.950 859.050 485.400 ;
        RECT 877.950 483.600 880.050 484.050 ;
        RECT 842.400 482.400 880.050 483.600 ;
        RECT 881.400 483.600 882.600 485.400 ;
        RECT 925.950 484.950 928.050 487.050 ;
        RECT 919.950 483.600 922.050 484.050 ;
        RECT 881.400 482.400 922.050 483.600 ;
        RECT 811.950 481.950 814.050 482.400 ;
        RECT 832.950 481.950 835.050 482.400 ;
        RECT 838.950 481.950 841.050 482.400 ;
        RECT 877.950 481.950 880.050 482.400 ;
        RECT 919.950 481.950 922.050 482.400 ;
        RECT 976.950 483.600 979.050 484.050 ;
        RECT 982.950 483.600 985.050 484.050 ;
        RECT 976.950 482.400 985.050 483.600 ;
        RECT 976.950 481.950 979.050 482.400 ;
        RECT 982.950 481.950 985.050 482.400 ;
        RECT 817.950 480.600 820.050 481.050 ;
        RECT 853.800 480.600 855.900 481.050 ;
        RECT 817.950 479.400 855.900 480.600 ;
        RECT 817.950 478.950 820.050 479.400 ;
        RECT 853.800 478.950 855.900 479.400 ;
        RECT 856.950 480.600 859.050 481.050 ;
        RECT 913.950 480.600 916.050 481.050 ;
        RECT 856.950 479.400 916.050 480.600 ;
        RECT 856.950 478.950 859.050 479.400 ;
        RECT 913.950 478.950 916.050 479.400 ;
        RECT 940.950 480.600 943.050 481.050 ;
        RECT 973.950 480.600 976.050 481.050 ;
        RECT 940.950 479.400 976.050 480.600 ;
        RECT 940.950 478.950 943.050 479.400 ;
        RECT 973.950 478.950 976.050 479.400 ;
        RECT 994.950 480.600 997.050 481.050 ;
        RECT 1000.950 480.600 1003.050 481.050 ;
        RECT 994.950 479.400 1003.050 480.600 ;
        RECT 994.950 478.950 997.050 479.400 ;
        RECT 1000.950 478.950 1003.050 479.400 ;
        RECT 670.950 476.400 732.600 477.600 ;
        RECT 802.950 477.600 805.050 478.050 ;
        RECT 808.950 477.600 811.050 478.050 ;
        RECT 802.950 476.400 811.050 477.600 ;
        RECT 670.950 475.950 673.050 476.400 ;
        RECT 802.950 475.950 805.050 476.400 ;
        RECT 808.950 475.950 811.050 476.400 ;
        RECT 814.950 477.600 817.050 478.050 ;
        RECT 865.950 477.600 868.050 478.050 ;
        RECT 814.950 476.400 868.050 477.600 ;
        RECT 814.950 475.950 817.050 476.400 ;
        RECT 865.950 475.950 868.050 476.400 ;
        RECT 874.950 477.600 877.050 478.050 ;
        RECT 892.950 477.600 895.050 478.050 ;
        RECT 874.950 476.400 895.050 477.600 ;
        RECT 874.950 475.950 877.050 476.400 ;
        RECT 892.950 475.950 895.050 476.400 ;
        RECT 946.950 477.600 949.050 478.050 ;
        RECT 982.950 477.600 985.050 478.050 ;
        RECT 946.950 476.400 985.050 477.600 ;
        RECT 946.950 475.950 949.050 476.400 ;
        RECT 982.950 475.950 985.050 476.400 ;
        RECT 1003.950 477.600 1006.050 478.050 ;
        RECT 1012.950 477.600 1015.050 478.050 ;
        RECT 1003.950 476.400 1015.050 477.600 ;
        RECT 1003.950 475.950 1006.050 476.400 ;
        RECT 1012.950 475.950 1015.050 476.400 ;
        RECT 211.950 473.400 435.600 474.600 ;
        RECT 625.950 474.600 628.050 475.050 ;
        RECT 652.950 474.600 655.050 475.050 ;
        RECT 625.950 473.400 655.050 474.600 ;
        RECT 211.950 472.950 214.050 473.400 ;
        RECT 625.950 472.950 628.050 473.400 ;
        RECT 652.950 472.950 655.050 473.400 ;
        RECT 757.950 474.600 760.050 475.050 ;
        RECT 811.950 474.600 814.050 475.050 ;
        RECT 757.950 473.400 814.050 474.600 ;
        RECT 757.950 472.950 760.050 473.400 ;
        RECT 811.950 472.950 814.050 473.400 ;
        RECT 919.950 474.600 922.050 475.050 ;
        RECT 934.950 474.600 937.050 475.050 ;
        RECT 970.800 474.600 972.900 475.050 ;
        RECT 919.950 473.400 972.900 474.600 ;
        RECT 919.950 472.950 922.050 473.400 ;
        RECT 934.950 472.950 937.050 473.400 ;
        RECT 970.800 472.950 972.900 473.400 ;
        RECT 973.950 474.600 976.050 475.050 ;
        RECT 988.950 474.600 991.050 475.050 ;
        RECT 973.950 473.400 991.050 474.600 ;
        RECT 973.950 472.950 976.050 473.400 ;
        RECT 988.950 472.950 991.050 473.400 ;
        RECT 256.950 471.600 259.050 472.050 ;
        RECT 358.950 471.600 361.050 472.050 ;
        RECT 382.950 471.600 385.050 472.050 ;
        RECT 424.950 471.600 427.050 472.050 ;
        RECT 256.950 470.400 427.050 471.600 ;
        RECT 256.950 469.950 259.050 470.400 ;
        RECT 358.950 469.950 361.050 470.400 ;
        RECT 382.950 469.950 385.050 470.400 ;
        RECT 424.950 469.950 427.050 470.400 ;
        RECT 439.950 471.600 442.050 472.050 ;
        RECT 511.950 471.600 514.050 472.050 ;
        RECT 439.950 470.400 514.050 471.600 ;
        RECT 439.950 469.950 442.050 470.400 ;
        RECT 511.950 469.950 514.050 470.400 ;
        RECT 526.950 471.600 529.050 472.050 ;
        RECT 547.950 471.600 550.050 472.050 ;
        RECT 526.950 470.400 550.050 471.600 ;
        RECT 526.950 469.950 529.050 470.400 ;
        RECT 547.950 469.950 550.050 470.400 ;
        RECT 604.950 471.600 607.050 472.050 ;
        RECT 667.950 471.600 670.050 472.050 ;
        RECT 604.950 470.400 670.050 471.600 ;
        RECT 604.950 469.950 607.050 470.400 ;
        RECT 667.950 469.950 670.050 470.400 ;
        RECT 685.950 471.600 688.050 472.050 ;
        RECT 718.950 471.600 721.050 472.050 ;
        RECT 685.950 470.400 721.050 471.600 ;
        RECT 685.950 469.950 688.050 470.400 ;
        RECT 718.950 469.950 721.050 470.400 ;
        RECT 778.950 471.600 781.050 472.050 ;
        RECT 838.950 471.600 841.050 472.050 ;
        RECT 778.950 470.400 841.050 471.600 ;
        RECT 778.950 469.950 781.050 470.400 ;
        RECT 838.950 469.950 841.050 470.400 ;
        RECT 844.950 471.600 847.050 472.050 ;
        RECT 850.950 471.600 853.050 472.050 ;
        RECT 844.950 470.400 853.050 471.600 ;
        RECT 844.950 469.950 847.050 470.400 ;
        RECT 850.950 469.950 853.050 470.400 ;
        RECT 913.950 471.600 916.050 472.050 ;
        RECT 928.950 471.600 931.050 472.050 ;
        RECT 913.950 470.400 931.050 471.600 ;
        RECT 913.950 469.950 916.050 470.400 ;
        RECT 928.950 469.950 931.050 470.400 ;
        RECT 964.950 471.600 967.050 472.050 ;
        RECT 994.950 471.600 997.050 472.050 ;
        RECT 964.950 470.400 997.050 471.600 ;
        RECT 964.950 469.950 967.050 470.400 ;
        RECT 994.950 469.950 997.050 470.400 ;
        RECT 1003.950 471.600 1006.050 472.050 ;
        RECT 1015.950 471.600 1018.050 472.050 ;
        RECT 1003.950 470.400 1018.050 471.600 ;
        RECT 1003.950 469.950 1006.050 470.400 ;
        RECT 1015.950 469.950 1018.050 470.400 ;
        RECT 28.950 468.600 31.050 469.050 ;
        RECT 37.950 468.600 40.050 469.050 ;
        RECT 28.950 467.400 40.050 468.600 ;
        RECT 28.950 466.950 31.050 467.400 ;
        RECT 37.950 466.950 40.050 467.400 ;
        RECT 64.950 468.600 67.050 469.050 ;
        RECT 148.950 468.600 151.050 469.050 ;
        RECT 64.950 467.400 151.050 468.600 ;
        RECT 64.950 466.950 67.050 467.400 ;
        RECT 148.950 466.950 151.050 467.400 ;
        RECT 199.950 468.600 202.050 469.050 ;
        RECT 223.950 468.600 226.050 469.050 ;
        RECT 199.950 467.400 226.050 468.600 ;
        RECT 199.950 466.950 202.050 467.400 ;
        RECT 223.950 466.950 226.050 467.400 ;
        RECT 394.950 468.600 397.050 469.050 ;
        RECT 415.950 468.600 418.050 469.050 ;
        RECT 394.950 467.400 418.050 468.600 ;
        RECT 394.950 466.950 397.050 467.400 ;
        RECT 415.950 466.950 418.050 467.400 ;
        RECT 445.950 468.600 448.050 469.050 ;
        RECT 475.950 468.600 478.050 469.050 ;
        RECT 445.950 467.400 478.050 468.600 ;
        RECT 445.950 466.950 448.050 467.400 ;
        RECT 475.950 466.950 478.050 467.400 ;
        RECT 682.950 468.600 685.050 469.050 ;
        RECT 724.950 468.600 727.050 469.050 ;
        RECT 682.950 467.400 727.050 468.600 ;
        RECT 682.950 466.950 685.050 467.400 ;
        RECT 724.950 466.950 727.050 467.400 ;
        RECT 754.950 468.600 757.050 469.050 ;
        RECT 784.950 468.600 787.050 469.050 ;
        RECT 754.950 467.400 787.050 468.600 ;
        RECT 754.950 466.950 757.050 467.400 ;
        RECT 784.950 466.950 787.050 467.400 ;
        RECT 811.950 468.600 814.050 469.050 ;
        RECT 817.950 468.600 820.050 469.050 ;
        RECT 811.950 467.400 820.050 468.600 ;
        RECT 811.950 466.950 814.050 467.400 ;
        RECT 817.950 466.950 820.050 467.400 ;
        RECT 853.950 468.600 856.050 469.050 ;
        RECT 859.950 468.600 862.050 469.050 ;
        RECT 853.950 467.400 862.050 468.600 ;
        RECT 853.950 466.950 856.050 467.400 ;
        RECT 859.950 466.950 862.050 467.400 ;
        RECT 865.950 468.600 868.050 469.050 ;
        RECT 919.950 468.600 922.050 469.050 ;
        RECT 865.950 467.400 922.050 468.600 ;
        RECT 929.400 468.600 930.600 469.950 ;
        RECT 949.950 468.600 952.050 469.050 ;
        RECT 929.400 467.400 952.050 468.600 ;
        RECT 865.950 466.950 868.050 467.400 ;
        RECT 919.950 466.950 922.050 467.400 ;
        RECT 949.950 466.950 952.050 467.400 ;
        RECT 970.950 468.600 973.050 469.050 ;
        RECT 1024.950 468.600 1027.050 469.050 ;
        RECT 970.950 467.400 1027.050 468.600 ;
        RECT 970.950 466.950 973.050 467.400 ;
        RECT 1024.950 466.950 1027.050 467.400 ;
        RECT 601.950 465.600 604.050 466.050 ;
        RECT 607.950 465.600 610.050 466.050 ;
        RECT 643.950 465.600 646.050 466.050 ;
        RECT 755.400 465.600 756.600 466.950 ;
        RECT 601.950 464.400 756.600 465.600 ;
        RECT 763.950 465.600 766.050 466.050 ;
        RECT 775.950 465.600 778.050 466.050 ;
        RECT 763.950 464.400 778.050 465.600 ;
        RECT 601.950 463.950 604.050 464.400 ;
        RECT 607.950 463.950 610.050 464.400 ;
        RECT 643.950 463.950 646.050 464.400 ;
        RECT 763.950 463.950 766.050 464.400 ;
        RECT 775.950 463.950 778.050 464.400 ;
        RECT 793.950 465.600 796.050 466.050 ;
        RECT 808.950 465.600 811.050 466.050 ;
        RECT 793.950 464.400 811.050 465.600 ;
        RECT 793.950 463.950 796.050 464.400 ;
        RECT 808.950 463.950 811.050 464.400 ;
        RECT 817.950 465.600 820.050 465.900 ;
        RECT 826.950 465.600 829.050 466.050 ;
        RECT 844.950 465.600 847.050 466.050 ;
        RECT 817.950 464.400 847.050 465.600 ;
        RECT 817.950 463.800 820.050 464.400 ;
        RECT 826.950 463.950 829.050 464.400 ;
        RECT 844.950 463.950 847.050 464.400 ;
        RECT 889.950 465.600 892.050 466.050 ;
        RECT 946.950 465.600 949.050 466.050 ;
        RECT 889.950 464.400 949.050 465.600 ;
        RECT 889.950 463.950 892.050 464.400 ;
        RECT 946.950 463.950 949.050 464.400 ;
        RECT 991.950 465.600 994.050 466.050 ;
        RECT 1033.950 465.600 1036.050 466.050 ;
        RECT 991.950 464.400 1036.050 465.600 ;
        RECT 991.950 463.950 994.050 464.400 ;
        RECT 1033.950 463.950 1036.050 464.400 ;
        RECT 229.950 462.600 232.050 463.050 ;
        RECT 361.950 462.600 364.050 463.050 ;
        RECT 229.950 461.400 364.050 462.600 ;
        RECT 229.950 460.950 232.050 461.400 ;
        RECT 361.950 460.950 364.050 461.400 ;
        RECT 373.950 462.600 376.050 463.050 ;
        RECT 397.950 462.600 400.050 463.050 ;
        RECT 373.950 461.400 400.050 462.600 ;
        RECT 373.950 460.950 376.050 461.400 ;
        RECT 397.950 460.950 400.050 461.400 ;
        RECT 610.950 462.600 613.050 463.050 ;
        RECT 670.950 462.600 673.050 463.050 ;
        RECT 610.950 461.400 673.050 462.600 ;
        RECT 610.950 460.950 613.050 461.400 ;
        RECT 670.950 460.950 673.050 461.400 ;
        RECT 784.950 462.600 787.050 463.050 ;
        RECT 859.950 462.600 862.050 463.050 ;
        RECT 784.950 461.400 862.050 462.600 ;
        RECT 784.950 460.950 787.050 461.400 ;
        RECT 859.950 460.950 862.050 461.400 ;
        RECT 910.950 462.600 913.050 463.050 ;
        RECT 916.800 462.600 918.900 463.050 ;
        RECT 910.950 461.400 918.900 462.600 ;
        RECT 910.950 460.950 913.050 461.400 ;
        RECT 916.800 460.950 918.900 461.400 ;
        RECT 919.950 462.600 922.050 463.050 ;
        RECT 958.950 462.600 961.050 463.050 ;
        RECT 919.950 461.400 961.050 462.600 ;
        RECT 919.950 460.950 922.050 461.400 ;
        RECT 958.950 460.950 961.050 461.400 ;
        RECT 967.950 462.600 970.050 463.050 ;
        RECT 1018.950 462.600 1021.050 463.050 ;
        RECT 967.950 461.400 1021.050 462.600 ;
        RECT 967.950 460.950 970.050 461.400 ;
        RECT 1018.950 460.950 1021.050 461.400 ;
        RECT 58.950 459.600 61.050 460.050 ;
        RECT 115.950 459.600 118.050 460.050 ;
        RECT 58.950 458.400 118.050 459.600 ;
        RECT 58.950 457.950 61.050 458.400 ;
        RECT 115.950 457.950 118.050 458.400 ;
        RECT 172.950 459.600 175.050 460.050 ;
        RECT 211.950 459.600 214.050 460.050 ;
        RECT 172.950 458.400 214.050 459.600 ;
        RECT 172.950 457.950 175.050 458.400 ;
        RECT 211.950 457.950 214.050 458.400 ;
        RECT 511.950 459.600 514.050 460.050 ;
        RECT 532.950 459.600 535.050 460.050 ;
        RECT 511.950 458.400 535.050 459.600 ;
        RECT 511.950 457.950 514.050 458.400 ;
        RECT 532.950 457.950 535.050 458.400 ;
        RECT 541.950 459.600 544.050 460.050 ;
        RECT 601.950 459.600 604.050 460.050 ;
        RECT 712.950 459.600 715.050 460.050 ;
        RECT 541.950 458.400 604.050 459.600 ;
        RECT 541.950 457.950 544.050 458.400 ;
        RECT 601.950 457.950 604.050 458.400 ;
        RECT 689.400 458.400 715.050 459.600 ;
        RECT 70.950 456.600 73.050 457.050 ;
        RECT 400.950 456.600 403.050 457.050 ;
        RECT 538.950 456.600 541.050 457.050 ;
        RECT 70.950 455.400 403.050 456.600 ;
        RECT 70.950 454.950 73.050 455.400 ;
        RECT 400.950 454.950 403.050 455.400 ;
        RECT 506.400 455.400 541.050 456.600 ;
        RECT 4.950 453.600 7.050 454.200 ;
        RECT 13.950 453.600 16.050 454.050 ;
        RECT 4.950 452.400 16.050 453.600 ;
        RECT 4.950 452.100 7.050 452.400 ;
        RECT 13.950 451.950 16.050 452.400 ;
        RECT 187.950 453.600 190.050 454.050 ;
        RECT 196.950 453.600 199.050 454.050 ;
        RECT 187.950 452.400 199.050 453.600 ;
        RECT 187.950 451.950 190.050 452.400 ;
        RECT 196.950 451.950 199.050 452.400 ;
        RECT 268.950 453.600 271.050 454.050 ;
        RECT 283.950 453.600 286.050 454.050 ;
        RECT 268.950 452.400 286.050 453.600 ;
        RECT 268.950 451.950 271.050 452.400 ;
        RECT 283.950 451.950 286.050 452.400 ;
        RECT 349.950 453.600 352.050 454.050 ;
        RECT 358.950 453.600 361.050 454.050 ;
        RECT 349.950 452.400 361.050 453.600 ;
        RECT 349.950 451.950 352.050 452.400 ;
        RECT 358.950 451.950 361.050 452.400 ;
        RECT 439.950 453.600 442.050 454.050 ;
        RECT 445.950 453.600 448.050 454.050 ;
        RECT 439.950 452.400 448.050 453.600 ;
        RECT 439.950 451.950 442.050 452.400 ;
        RECT 445.950 451.950 448.050 452.400 ;
        RECT 88.950 450.600 91.050 451.200 ;
        RECT 100.950 450.600 103.050 451.050 ;
        RECT 88.950 449.400 103.050 450.600 ;
        RECT 88.950 449.100 91.050 449.400 ;
        RECT 100.950 448.950 103.050 449.400 ;
        RECT 109.950 449.100 112.050 451.200 ;
        RECT 145.950 450.750 148.050 451.200 ;
        RECT 157.950 450.750 160.050 451.200 ;
        RECT 145.950 449.550 160.050 450.750 ;
        RECT 145.950 449.100 148.050 449.550 ;
        RECT 157.950 449.100 160.050 449.550 ;
        RECT 163.950 449.100 166.050 451.200 ;
        RECT 175.950 450.750 178.050 451.200 ;
        RECT 184.950 450.750 187.050 451.200 ;
        RECT 175.950 449.550 187.050 450.750 ;
        RECT 175.950 449.100 178.050 449.550 ;
        RECT 184.950 449.100 187.050 449.550 ;
        RECT 217.950 450.750 220.050 451.200 ;
        RECT 223.950 450.750 226.050 451.200 ;
        RECT 217.950 449.550 226.050 450.750 ;
        RECT 217.950 449.100 220.050 449.550 ;
        RECT 223.950 449.100 226.050 449.550 ;
        RECT 241.950 449.100 244.050 451.200 ;
        RECT 247.950 450.750 250.050 451.200 ;
        RECT 256.950 450.750 259.050 451.200 ;
        RECT 247.950 449.550 259.050 450.750 ;
        RECT 247.950 449.100 250.050 449.550 ;
        RECT 256.950 449.100 259.050 449.550 ;
        RECT 262.950 450.600 265.050 451.050 ;
        RECT 283.950 450.600 286.050 450.900 ;
        RECT 262.950 449.400 286.050 450.600 ;
        RECT 110.400 447.600 111.600 449.100 ;
        RECT 110.400 446.400 138.600 447.600 ;
        RECT 10.950 444.600 13.050 445.050 ;
        RECT 49.950 444.600 52.050 445.050 ;
        RECT 10.950 443.400 52.050 444.600 ;
        RECT 10.950 442.950 13.050 443.400 ;
        RECT 49.950 442.950 52.050 443.400 ;
        RECT 64.950 444.600 67.050 445.050 ;
        RECT 76.950 444.600 79.050 445.050 ;
        RECT 64.950 443.400 79.050 444.600 ;
        RECT 64.950 442.950 67.050 443.400 ;
        RECT 76.950 442.950 79.050 443.400 ;
        RECT 85.950 444.600 88.050 444.900 ;
        RECT 106.950 444.600 109.050 444.900 ;
        RECT 85.950 443.400 109.050 444.600 ;
        RECT 85.950 442.800 88.050 443.400 ;
        RECT 106.950 442.800 109.050 443.400 ;
        RECT 118.950 444.450 121.050 444.900 ;
        RECT 133.950 444.450 136.050 444.900 ;
        RECT 118.950 443.250 136.050 444.450 ;
        RECT 137.400 444.600 138.600 446.400 ;
        RECT 160.950 444.600 163.050 444.900 ;
        RECT 137.400 443.400 163.050 444.600 ;
        RECT 164.400 444.600 165.600 449.100 ;
        RECT 169.950 444.600 172.050 445.050 ;
        RECT 187.950 444.600 190.050 444.900 ;
        RECT 164.400 443.400 190.050 444.600 ;
        RECT 242.400 444.600 243.600 449.100 ;
        RECT 262.950 448.950 265.050 449.400 ;
        RECT 283.950 448.800 286.050 449.400 ;
        RECT 322.950 448.950 325.050 451.050 ;
        RECT 340.950 450.600 343.050 451.200 ;
        RECT 364.950 450.600 367.050 451.200 ;
        RECT 388.950 450.600 391.050 451.200 ;
        RECT 409.950 450.600 412.050 451.200 ;
        RECT 340.950 449.400 412.050 450.600 ;
        RECT 340.950 449.100 343.050 449.400 ;
        RECT 364.950 449.100 367.050 449.400 ;
        RECT 388.950 449.100 391.050 449.400 ;
        RECT 409.950 449.100 412.050 449.400 ;
        RECT 427.950 450.600 430.050 450.900 ;
        RECT 436.950 450.600 439.050 451.200 ;
        RECT 427.950 449.400 439.050 450.600 ;
        RECT 323.400 445.050 324.600 448.950 ;
        RECT 427.950 448.800 430.050 449.400 ;
        RECT 436.950 449.100 439.050 449.400 ;
        RECT 448.950 450.600 451.050 451.050 ;
        RECT 454.950 450.600 457.050 451.050 ;
        RECT 448.950 449.400 457.050 450.600 ;
        RECT 448.950 448.950 451.050 449.400 ;
        RECT 454.950 448.950 457.050 449.400 ;
        RECT 475.950 450.750 478.050 451.200 ;
        RECT 484.950 450.750 487.050 451.200 ;
        RECT 475.950 449.550 487.050 450.750 ;
        RECT 475.950 449.100 478.050 449.550 ;
        RECT 484.950 449.100 487.050 449.550 ;
        RECT 490.950 450.600 493.050 451.200 ;
        RECT 502.950 450.600 505.050 451.050 ;
        RECT 506.400 450.600 507.600 455.400 ;
        RECT 538.950 454.950 541.050 455.400 ;
        RECT 553.950 456.600 556.050 457.050 ;
        RECT 610.950 456.600 613.050 457.050 ;
        RECT 553.950 455.400 613.050 456.600 ;
        RECT 553.950 454.950 556.050 455.400 ;
        RECT 610.950 454.950 613.050 455.400 ;
        RECT 631.950 456.600 634.050 457.050 ;
        RECT 689.400 456.600 690.600 458.400 ;
        RECT 712.950 457.950 715.050 458.400 ;
        RECT 721.950 459.600 724.050 460.050 ;
        RECT 796.950 459.600 799.050 460.050 ;
        RECT 826.950 459.600 829.050 460.050 ;
        RECT 721.950 458.400 777.600 459.600 ;
        RECT 721.950 457.950 724.050 458.400 ;
        RECT 631.950 455.400 690.600 456.600 ;
        RECT 718.950 456.600 721.050 457.050 ;
        RECT 776.400 456.600 777.600 458.400 ;
        RECT 796.950 458.400 829.050 459.600 ;
        RECT 796.950 457.950 799.050 458.400 ;
        RECT 826.950 457.950 829.050 458.400 ;
        RECT 838.950 459.600 841.050 460.050 ;
        RECT 856.950 459.600 859.050 460.050 ;
        RECT 838.950 458.400 859.050 459.600 ;
        RECT 838.950 457.950 841.050 458.400 ;
        RECT 856.950 457.950 859.050 458.400 ;
        RECT 934.950 459.600 937.050 460.050 ;
        RECT 961.950 459.600 964.050 460.050 ;
        RECT 934.950 458.400 964.050 459.600 ;
        RECT 934.950 457.950 937.050 458.400 ;
        RECT 961.950 457.950 964.050 458.400 ;
        RECT 982.800 459.000 984.900 460.050 ;
        RECT 985.950 459.600 988.050 460.050 ;
        RECT 1000.950 459.600 1003.050 460.050 ;
        RECT 982.800 457.950 985.050 459.000 ;
        RECT 985.950 458.400 1003.050 459.600 ;
        RECT 985.950 457.950 988.050 458.400 ;
        RECT 1000.950 457.950 1003.050 458.400 ;
        RECT 820.950 456.600 823.050 456.900 ;
        RECT 718.950 455.400 741.600 456.600 ;
        RECT 776.400 455.400 823.050 456.600 ;
        RECT 631.950 454.950 634.050 455.400 ;
        RECT 718.950 454.950 721.050 455.400 ;
        RECT 580.950 453.600 583.050 454.050 ;
        RECT 613.950 453.600 616.050 454.050 ;
        RECT 580.950 452.400 616.050 453.600 ;
        RECT 580.950 451.950 583.050 452.400 ;
        RECT 613.950 451.950 616.050 452.400 ;
        RECT 691.950 453.600 694.050 454.050 ;
        RECT 697.950 453.600 700.050 454.050 ;
        RECT 715.950 453.600 718.050 454.050 ;
        RECT 691.950 452.400 718.050 453.600 ;
        RECT 691.950 451.950 694.050 452.400 ;
        RECT 697.950 451.950 700.050 452.400 ;
        RECT 715.950 451.950 718.050 452.400 ;
        RECT 727.950 453.600 732.000 454.050 ;
        RECT 727.950 451.950 732.600 453.600 ;
        RECT 736.950 451.950 739.050 454.050 ;
        RECT 740.400 453.600 741.600 455.400 ;
        RECT 820.950 454.800 823.050 455.400 ;
        RECT 859.950 456.600 862.050 457.050 ;
        RECT 865.950 456.600 868.050 457.050 ;
        RECT 859.950 455.400 868.050 456.600 ;
        RECT 859.950 454.950 862.050 455.400 ;
        RECT 865.950 454.950 868.050 455.400 ;
        RECT 919.950 456.600 922.050 457.050 ;
        RECT 964.950 456.600 967.050 457.050 ;
        RECT 919.950 455.400 967.050 456.600 ;
        RECT 982.950 456.600 985.050 457.950 ;
        RECT 1027.950 456.600 1030.050 457.050 ;
        RECT 982.950 456.000 1030.050 456.600 ;
        RECT 983.400 455.400 1030.050 456.000 ;
        RECT 919.950 454.950 922.050 455.400 ;
        RECT 964.950 454.950 967.050 455.400 ;
        RECT 1027.950 454.950 1030.050 455.400 ;
        RECT 805.950 453.600 808.050 454.050 ;
        RECT 740.400 452.400 808.050 453.600 ;
        RECT 805.950 451.950 808.050 452.400 ;
        RECT 841.950 453.600 844.050 454.050 ;
        RECT 853.950 453.600 856.050 454.050 ;
        RECT 841.950 452.400 856.050 453.600 ;
        RECT 841.950 451.950 844.050 452.400 ;
        RECT 853.950 451.950 856.050 452.400 ;
        RECT 490.950 449.400 507.600 450.600 ;
        RECT 514.950 450.750 517.050 451.200 ;
        RECT 520.800 450.750 522.900 451.200 ;
        RECT 514.950 449.550 522.900 450.750 ;
        RECT 490.950 449.100 493.050 449.400 ;
        RECT 502.950 448.950 505.050 449.400 ;
        RECT 514.950 449.100 517.050 449.550 ;
        RECT 520.800 449.100 522.900 449.550 ;
        RECT 523.950 450.750 526.050 451.200 ;
        RECT 538.950 450.750 541.050 451.200 ;
        RECT 523.950 449.550 541.050 450.750 ;
        RECT 523.950 449.100 526.050 449.550 ;
        RECT 538.950 449.100 541.050 449.550 ;
        RECT 559.950 449.100 562.050 451.200 ;
        RECT 565.950 450.750 568.050 451.200 ;
        RECT 574.950 450.750 577.050 451.200 ;
        RECT 565.950 449.550 577.050 450.750 ;
        RECT 565.950 449.100 568.050 449.550 ;
        RECT 574.950 449.100 577.050 449.550 ;
        RECT 589.950 450.600 592.050 451.200 ;
        RECT 598.950 450.600 601.050 451.050 ;
        RECT 589.950 449.400 601.050 450.600 ;
        RECT 589.950 449.100 592.050 449.400 ;
        RECT 325.950 447.600 328.050 448.050 ;
        RECT 349.950 447.600 352.050 448.050 ;
        RECT 325.950 446.400 352.050 447.600 ;
        RECT 325.950 445.950 328.050 446.400 ;
        RECT 349.950 445.950 352.050 446.400 ;
        RECT 250.950 444.600 253.050 445.050 ;
        RECT 242.400 443.400 253.050 444.600 ;
        RECT 118.950 442.800 121.050 443.250 ;
        RECT 133.950 442.800 136.050 443.250 ;
        RECT 160.950 442.800 163.050 443.400 ;
        RECT 169.950 442.950 172.050 443.400 ;
        RECT 187.950 442.800 190.050 443.400 ;
        RECT 250.950 442.950 253.050 443.400 ;
        RECT 265.950 444.450 268.050 444.900 ;
        RECT 298.950 444.450 301.050 444.900 ;
        RECT 265.950 443.250 301.050 444.450 ;
        RECT 265.950 442.800 268.050 443.250 ;
        RECT 298.950 442.800 301.050 443.250 ;
        RECT 307.950 444.450 310.050 444.900 ;
        RECT 313.950 444.450 316.050 444.900 ;
        RECT 307.950 443.250 316.050 444.450 ;
        RECT 307.950 442.800 310.050 443.250 ;
        RECT 313.950 442.800 316.050 443.250 ;
        RECT 322.950 442.950 325.050 445.050 ;
        RECT 331.950 444.600 334.050 445.050 ;
        RECT 343.950 444.600 346.050 445.050 ;
        RECT 331.950 443.400 346.050 444.600 ;
        RECT 331.950 442.950 334.050 443.400 ;
        RECT 343.950 442.950 346.050 443.400 ;
        RECT 361.950 444.600 364.050 444.900 ;
        RECT 370.800 444.600 372.900 445.050 ;
        RECT 361.950 443.400 372.900 444.600 ;
        RECT 361.950 442.800 364.050 443.400 ;
        RECT 370.800 442.950 372.900 443.400 ;
        RECT 373.950 444.450 376.050 444.900 ;
        RECT 385.950 444.450 388.050 444.900 ;
        RECT 373.950 443.250 388.050 444.450 ;
        RECT 373.950 442.800 376.050 443.250 ;
        RECT 385.950 442.800 388.050 443.250 ;
        RECT 412.950 444.600 415.050 444.900 ;
        RECT 433.950 444.600 436.050 444.900 ;
        RECT 412.950 443.400 436.050 444.600 ;
        RECT 412.950 442.800 415.050 443.400 ;
        RECT 433.950 442.800 436.050 443.400 ;
        RECT 463.950 444.600 466.050 444.900 ;
        RECT 478.950 444.600 481.050 445.050 ;
        RECT 463.950 443.400 481.050 444.600 ;
        RECT 463.950 442.800 466.050 443.400 ;
        RECT 478.950 442.950 481.050 443.400 ;
        RECT 493.950 444.600 496.050 445.050 ;
        RECT 526.950 444.600 529.050 445.050 ;
        RECT 493.950 443.400 529.050 444.600 ;
        RECT 493.950 442.950 496.050 443.400 ;
        RECT 526.950 442.950 529.050 443.400 ;
        RECT 541.950 444.600 544.050 444.900 ;
        RECT 547.950 444.600 550.050 445.050 ;
        RECT 541.950 443.400 550.050 444.600 ;
        RECT 541.950 442.800 544.050 443.400 ;
        RECT 547.950 442.950 550.050 443.400 ;
        RECT 560.400 442.050 561.600 449.100 ;
        RECT 598.950 448.950 601.050 449.400 ;
        RECT 640.950 450.600 643.050 451.200 ;
        RECT 646.950 450.600 649.050 450.900 ;
        RECT 640.950 449.400 649.050 450.600 ;
        RECT 640.950 449.100 643.050 449.400 ;
        RECT 646.950 448.800 649.050 449.400 ;
        RECT 652.950 450.750 655.050 451.200 ;
        RECT 664.950 450.750 667.050 451.200 ;
        RECT 652.950 449.550 667.050 450.750 ;
        RECT 721.950 450.600 724.050 451.050 ;
        RECT 652.950 449.100 655.050 449.550 ;
        RECT 664.950 449.100 667.050 449.550 ;
        RECT 689.400 449.400 724.050 450.600 ;
        RECT 731.400 450.600 732.600 451.950 ;
        RECT 731.400 449.400 735.600 450.600 ;
        RECT 689.400 447.600 690.600 449.400 ;
        RECT 721.950 448.950 724.050 449.400 ;
        RECT 734.400 447.900 735.600 449.400 ;
        RECT 737.400 448.050 738.600 451.950 ;
        RECT 823.950 450.600 826.050 451.050 ;
        RECT 794.400 449.400 826.050 450.600 ;
        RECT 593.400 446.400 690.600 447.600 ;
        RECT 593.400 444.900 594.600 446.400 ;
        RECT 733.800 445.800 735.900 447.900 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 760.950 446.100 763.050 448.200 ;
        RECT 580.950 444.450 583.050 444.900 ;
        RECT 586.950 444.450 589.050 444.900 ;
        RECT 580.950 443.250 589.050 444.450 ;
        RECT 580.950 442.800 583.050 443.250 ;
        RECT 586.950 442.800 589.050 443.250 ;
        RECT 592.950 442.800 595.050 444.900 ;
        RECT 598.950 444.450 601.050 444.900 ;
        RECT 619.950 444.600 622.050 444.900 ;
        RECT 637.950 444.600 640.050 444.900 ;
        RECT 619.950 444.450 640.050 444.600 ;
        RECT 598.950 443.400 640.050 444.450 ;
        RECT 598.950 443.250 622.050 443.400 ;
        RECT 598.950 442.800 601.050 443.250 ;
        RECT 619.950 442.800 622.050 443.250 ;
        RECT 637.950 442.800 640.050 443.400 ;
        RECT 646.950 444.450 649.050 444.900 ;
        RECT 661.950 444.450 664.050 444.900 ;
        RECT 646.950 443.250 664.050 444.450 ;
        RECT 646.950 442.800 649.050 443.250 ;
        RECT 661.950 442.800 664.050 443.250 ;
        RECT 697.950 444.450 700.050 444.900 ;
        RECT 715.950 444.450 718.050 444.900 ;
        RECT 697.950 443.250 718.050 444.450 ;
        RECT 697.950 442.800 700.050 443.250 ;
        RECT 715.950 442.800 718.050 443.250 ;
        RECT 133.950 441.600 136.050 442.050 ;
        RECT 166.950 441.600 169.050 442.050 ;
        RECT 133.950 440.400 169.050 441.600 ;
        RECT 133.950 439.950 136.050 440.400 ;
        RECT 166.950 439.950 169.050 440.400 ;
        RECT 220.950 441.600 223.050 442.050 ;
        RECT 256.950 441.600 259.050 442.050 ;
        RECT 418.950 441.600 421.050 442.050 ;
        RECT 220.950 440.400 259.050 441.600 ;
        RECT 220.950 439.950 223.050 440.400 ;
        RECT 256.950 439.950 259.050 440.400 ;
        RECT 296.400 440.400 421.050 441.600 ;
        RECT 55.950 438.600 58.050 439.050 ;
        RECT 70.950 438.600 73.050 439.050 ;
        RECT 106.950 438.600 109.050 439.050 ;
        RECT 55.950 437.400 109.050 438.600 ;
        RECT 55.950 436.950 58.050 437.400 ;
        RECT 70.950 436.950 73.050 437.400 ;
        RECT 106.950 436.950 109.050 437.400 ;
        RECT 151.950 438.600 154.050 439.050 ;
        RECT 296.400 438.600 297.600 440.400 ;
        RECT 418.950 439.950 421.050 440.400 ;
        RECT 481.950 441.600 484.050 442.050 ;
        RECT 487.950 441.600 490.050 442.050 ;
        RECT 517.950 441.600 520.050 442.050 ;
        RECT 481.950 440.400 490.050 441.600 ;
        RECT 481.950 439.950 484.050 440.400 ;
        RECT 487.950 439.950 490.050 440.400 ;
        RECT 509.400 440.400 520.050 441.600 ;
        RECT 151.950 437.400 297.600 438.600 ;
        RECT 298.950 438.600 301.050 439.050 ;
        RECT 337.950 438.600 340.050 439.050 ;
        RECT 298.950 437.400 340.050 438.600 ;
        RECT 151.950 436.950 154.050 437.400 ;
        RECT 298.950 436.950 301.050 437.400 ;
        RECT 337.950 436.950 340.050 437.400 ;
        RECT 451.950 438.600 454.050 439.050 ;
        RECT 463.950 438.600 466.050 439.050 ;
        RECT 451.950 437.400 466.050 438.600 ;
        RECT 451.950 436.950 454.050 437.400 ;
        RECT 463.950 436.950 466.050 437.400 ;
        RECT 472.950 438.600 475.050 438.900 ;
        RECT 509.400 438.600 510.600 440.400 ;
        RECT 517.950 439.950 520.050 440.400 ;
        RECT 559.950 439.950 562.050 442.050 ;
        RECT 727.950 441.600 730.050 442.050 ;
        RECT 739.950 441.600 742.050 442.050 ;
        RECT 727.950 440.400 742.050 441.600 ;
        RECT 761.400 441.600 762.600 446.100 ;
        RECT 784.950 444.600 787.050 445.050 ;
        RECT 794.400 444.600 795.600 449.400 ;
        RECT 823.950 448.950 826.050 449.400 ;
        RECT 961.950 450.750 964.050 451.200 ;
        RECT 967.950 450.750 970.050 451.200 ;
        RECT 961.950 449.550 970.050 450.750 ;
        RECT 961.950 449.100 964.050 449.550 ;
        RECT 967.950 449.100 970.050 449.550 ;
        RECT 1006.950 450.750 1009.050 451.200 ;
        RECT 1012.950 450.750 1015.050 451.200 ;
        RECT 1006.950 449.550 1015.050 450.750 ;
        RECT 1006.950 449.100 1009.050 449.550 ;
        RECT 1012.950 449.100 1015.050 449.550 ;
        RECT 868.950 447.600 871.050 448.050 ;
        RECT 886.800 447.600 888.900 448.050 ;
        RECT 868.950 446.400 888.900 447.600 ;
        RECT 868.950 445.950 871.050 446.400 ;
        RECT 886.800 445.950 888.900 446.400 ;
        RECT 889.950 446.100 892.050 448.200 ;
        RECT 910.950 447.450 913.050 447.900 ;
        RECT 916.950 447.450 919.050 447.900 ;
        RECT 910.950 446.250 919.050 447.450 ;
        RECT 784.950 443.400 795.600 444.600 ;
        RECT 808.950 444.450 811.050 444.900 ;
        RECT 814.950 444.600 817.050 445.050 ;
        RECT 835.950 444.600 838.050 444.900 ;
        RECT 814.950 444.450 838.050 444.600 ;
        RECT 808.950 443.400 838.050 444.450 ;
        RECT 784.950 442.950 787.050 443.400 ;
        RECT 808.950 443.250 817.050 443.400 ;
        RECT 808.950 442.800 811.050 443.250 ;
        RECT 814.950 442.950 817.050 443.250 ;
        RECT 835.950 442.800 838.050 443.400 ;
        RECT 781.950 441.600 784.050 442.050 ;
        RECT 761.400 440.400 784.050 441.600 ;
        RECT 727.950 439.950 730.050 440.400 ;
        RECT 739.950 439.950 742.050 440.400 ;
        RECT 781.950 439.950 784.050 440.400 ;
        RECT 472.950 437.400 510.600 438.600 ;
        RECT 511.950 438.600 514.050 439.050 ;
        RECT 523.950 438.600 526.050 439.050 ;
        RECT 511.950 437.400 526.050 438.600 ;
        RECT 472.950 436.800 475.050 437.400 ;
        RECT 511.950 436.950 514.050 437.400 ;
        RECT 523.950 436.950 526.050 437.400 ;
        RECT 535.950 438.600 538.050 439.050 ;
        RECT 562.950 438.600 565.050 439.050 ;
        RECT 652.950 438.600 655.050 439.050 ;
        RECT 535.950 437.400 565.050 438.600 ;
        RECT 535.950 436.950 538.050 437.400 ;
        RECT 562.950 436.950 565.050 437.400 ;
        RECT 608.400 437.400 655.050 438.600 ;
        RECT 112.950 435.600 115.050 436.050 ;
        RECT 148.950 435.600 151.050 436.050 ;
        RECT 112.950 434.400 151.050 435.600 ;
        RECT 112.950 433.950 115.050 434.400 ;
        RECT 148.950 433.950 151.050 434.400 ;
        RECT 217.950 435.600 220.050 436.050 ;
        RECT 319.950 435.600 322.050 436.050 ;
        RECT 217.950 434.400 322.050 435.600 ;
        RECT 217.950 433.950 220.050 434.400 ;
        RECT 319.950 433.950 322.050 434.400 ;
        RECT 400.950 435.600 403.050 436.050 ;
        RECT 493.950 435.600 496.050 436.050 ;
        RECT 608.400 435.600 609.600 437.400 ;
        RECT 652.950 436.950 655.050 437.400 ;
        RECT 664.950 438.600 667.050 439.050 ;
        RECT 724.950 438.600 727.050 439.050 ;
        RECT 664.950 437.400 727.050 438.600 ;
        RECT 664.950 436.950 667.050 437.400 ;
        RECT 724.950 436.950 727.050 437.400 ;
        RECT 811.950 438.600 814.050 439.050 ;
        RECT 853.950 438.600 856.050 439.050 ;
        RECT 811.950 437.400 856.050 438.600 ;
        RECT 811.950 436.950 814.050 437.400 ;
        RECT 853.950 436.950 856.050 437.400 ;
        RECT 400.950 434.400 496.050 435.600 ;
        RECT 400.950 433.950 403.050 434.400 ;
        RECT 493.950 433.950 496.050 434.400 ;
        RECT 548.400 434.400 609.600 435.600 ;
        RECT 610.950 435.600 613.050 436.050 ;
        RECT 649.950 435.600 652.050 436.050 ;
        RECT 787.950 435.600 790.050 436.050 ;
        RECT 610.950 434.400 652.050 435.600 ;
        RECT 184.950 432.600 187.050 433.050 ;
        RECT 265.950 432.600 268.050 433.050 ;
        RECT 184.950 431.400 268.050 432.600 ;
        RECT 184.950 430.950 187.050 431.400 ;
        RECT 265.950 430.950 268.050 431.400 ;
        RECT 313.950 432.600 316.050 433.050 ;
        RECT 328.950 432.600 331.050 433.050 ;
        RECT 313.950 431.400 331.050 432.600 ;
        RECT 313.950 430.950 316.050 431.400 ;
        RECT 328.950 430.950 331.050 431.400 ;
        RECT 397.950 432.600 400.050 433.050 ;
        RECT 439.950 432.600 442.050 433.050 ;
        RECT 397.950 431.400 442.050 432.600 ;
        RECT 397.950 430.950 400.050 431.400 ;
        RECT 439.950 430.950 442.050 431.400 ;
        RECT 457.950 432.600 460.050 433.050 ;
        RECT 466.950 432.600 469.050 433.050 ;
        RECT 457.950 431.400 469.050 432.600 ;
        RECT 457.950 430.950 460.050 431.400 ;
        RECT 466.950 430.950 469.050 431.400 ;
        RECT 517.950 432.600 520.050 433.050 ;
        RECT 548.400 432.600 549.600 434.400 ;
        RECT 610.950 433.950 613.050 434.400 ;
        RECT 649.950 433.950 652.050 434.400 ;
        RECT 758.400 434.400 790.050 435.600 ;
        RECT 571.950 432.600 574.050 433.050 ;
        RECT 517.950 431.400 549.600 432.600 ;
        RECT 551.400 431.400 574.050 432.600 ;
        RECT 517.950 430.950 520.050 431.400 ;
        RECT 208.950 429.600 211.050 430.050 ;
        RECT 247.950 429.600 250.050 430.050 ;
        RECT 208.950 428.400 250.050 429.600 ;
        RECT 208.950 427.950 211.050 428.400 ;
        RECT 247.950 427.950 250.050 428.400 ;
        RECT 256.950 429.600 259.050 430.050 ;
        RECT 271.950 429.600 274.050 430.050 ;
        RECT 256.950 428.400 274.050 429.600 ;
        RECT 256.950 427.950 259.050 428.400 ;
        RECT 271.950 427.950 274.050 428.400 ;
        RECT 403.950 429.600 406.050 430.050 ;
        RECT 424.950 429.600 427.050 430.050 ;
        RECT 403.950 428.400 427.050 429.600 ;
        RECT 403.950 427.950 406.050 428.400 ;
        RECT 424.950 427.950 427.050 428.400 ;
        RECT 502.950 429.600 505.050 430.050 ;
        RECT 514.950 429.600 517.050 430.050 ;
        RECT 502.950 428.400 517.050 429.600 ;
        RECT 502.950 427.950 505.050 428.400 ;
        RECT 514.950 427.950 517.050 428.400 ;
        RECT 544.950 429.600 547.050 430.050 ;
        RECT 551.400 429.600 552.600 431.400 ;
        RECT 571.950 430.950 574.050 431.400 ;
        RECT 613.950 432.600 616.050 433.050 ;
        RECT 631.950 432.600 634.050 433.050 ;
        RECT 613.950 431.400 634.050 432.600 ;
        RECT 613.950 430.950 616.050 431.400 ;
        RECT 631.950 430.950 634.050 431.400 ;
        RECT 667.950 432.600 670.050 433.050 ;
        RECT 724.950 432.600 727.050 433.050 ;
        RECT 667.950 431.400 727.050 432.600 ;
        RECT 667.950 430.950 670.050 431.400 ;
        RECT 724.950 430.950 727.050 431.400 ;
        RECT 544.950 428.400 552.600 429.600 ;
        RECT 577.950 429.600 580.050 430.050 ;
        RECT 589.950 429.600 592.050 430.050 ;
        RECT 577.950 428.400 592.050 429.600 ;
        RECT 544.950 427.950 547.050 428.400 ;
        RECT 577.950 427.950 580.050 428.400 ;
        RECT 589.950 427.950 592.050 428.400 ;
        RECT 601.950 429.600 604.050 430.050 ;
        RECT 640.950 429.600 643.050 430.050 ;
        RECT 601.950 428.400 643.050 429.600 ;
        RECT 601.950 427.950 604.050 428.400 ;
        RECT 640.950 427.950 643.050 428.400 ;
        RECT 751.950 429.600 754.050 430.050 ;
        RECT 758.400 429.600 759.600 434.400 ;
        RECT 787.950 433.950 790.050 434.400 ;
        RECT 793.950 435.600 796.050 436.050 ;
        RECT 823.950 435.600 826.050 436.050 ;
        RECT 793.950 434.400 826.050 435.600 ;
        RECT 793.950 433.950 796.050 434.400 ;
        RECT 823.950 433.950 826.050 434.400 ;
        RECT 763.950 432.600 766.050 433.050 ;
        RECT 796.950 432.600 799.050 433.050 ;
        RECT 763.950 431.400 799.050 432.600 ;
        RECT 763.950 430.950 766.050 431.400 ;
        RECT 796.950 430.950 799.050 431.400 ;
        RECT 802.950 432.600 805.050 433.050 ;
        RECT 817.950 432.600 820.050 433.050 ;
        RECT 802.950 431.400 820.050 432.600 ;
        RECT 802.950 430.950 805.050 431.400 ;
        RECT 817.950 430.950 820.050 431.400 ;
        RECT 829.950 432.600 832.050 433.050 ;
        RECT 838.950 432.600 841.050 433.050 ;
        RECT 829.950 431.400 841.050 432.600 ;
        RECT 829.950 430.950 832.050 431.400 ;
        RECT 838.950 430.950 841.050 431.400 ;
        RECT 868.950 432.600 871.050 433.050 ;
        RECT 883.950 432.600 886.050 433.050 ;
        RECT 868.950 431.400 886.050 432.600 ;
        RECT 890.400 432.600 891.600 446.100 ;
        RECT 910.950 445.800 913.050 446.250 ;
        RECT 916.950 445.800 919.050 446.250 ;
        RECT 946.950 444.600 949.050 444.900 ;
        RECT 946.950 443.400 951.600 444.600 ;
        RECT 946.950 442.800 949.050 443.400 ;
        RECT 925.950 441.600 928.050 442.050 ;
        RECT 943.950 441.600 946.050 442.050 ;
        RECT 925.950 440.400 946.050 441.600 ;
        RECT 950.400 441.600 951.600 443.400 ;
        RECT 964.950 444.450 967.050 444.900 ;
        RECT 979.950 444.450 982.050 444.900 ;
        RECT 964.950 443.250 982.050 444.450 ;
        RECT 964.950 442.800 967.050 443.250 ;
        RECT 979.950 442.800 982.050 443.250 ;
        RECT 1021.950 444.450 1024.050 444.900 ;
        RECT 1027.950 444.450 1030.050 444.900 ;
        RECT 1021.950 443.250 1030.050 444.450 ;
        RECT 1021.950 442.800 1024.050 443.250 ;
        RECT 1027.950 442.800 1030.050 443.250 ;
        RECT 961.950 441.600 964.050 442.050 ;
        RECT 950.400 440.400 964.050 441.600 ;
        RECT 925.950 439.950 928.050 440.400 ;
        RECT 943.950 439.950 946.050 440.400 ;
        RECT 961.950 439.950 964.050 440.400 ;
        RECT 1006.950 441.600 1009.050 442.050 ;
        RECT 1012.950 441.600 1015.050 442.050 ;
        RECT 1006.950 440.400 1015.050 441.600 ;
        RECT 1006.950 439.950 1009.050 440.400 ;
        RECT 1012.950 439.950 1015.050 440.400 ;
        RECT 910.950 438.600 913.050 439.050 ;
        RECT 922.950 438.600 925.050 439.050 ;
        RECT 910.950 437.400 925.050 438.600 ;
        RECT 910.950 436.950 913.050 437.400 ;
        RECT 922.950 436.950 925.050 437.400 ;
        RECT 928.950 435.600 931.050 436.050 ;
        RECT 985.950 435.600 988.050 436.050 ;
        RECT 928.950 434.400 988.050 435.600 ;
        RECT 928.950 433.950 931.050 434.400 ;
        RECT 985.950 433.950 988.050 434.400 ;
        RECT 997.950 435.600 1000.050 436.050 ;
        RECT 1015.950 435.600 1018.050 436.050 ;
        RECT 997.950 434.400 1018.050 435.600 ;
        RECT 997.950 433.950 1000.050 434.400 ;
        RECT 1015.950 433.950 1018.050 434.400 ;
        RECT 895.950 432.600 898.050 433.050 ;
        RECT 890.400 431.400 898.050 432.600 ;
        RECT 868.950 430.950 871.050 431.400 ;
        RECT 883.950 430.950 886.050 431.400 ;
        RECT 895.950 430.950 898.050 431.400 ;
        RECT 961.950 432.600 964.050 433.050 ;
        RECT 967.950 432.600 970.050 433.050 ;
        RECT 961.950 431.400 970.050 432.600 ;
        RECT 961.950 430.950 964.050 431.400 ;
        RECT 967.950 430.950 970.050 431.400 ;
        RECT 751.950 428.400 759.600 429.600 ;
        RECT 823.950 429.600 826.050 430.050 ;
        RECT 919.950 429.600 922.050 430.050 ;
        RECT 823.950 428.400 922.050 429.600 ;
        RECT 751.950 427.950 754.050 428.400 ;
        RECT 823.950 427.950 826.050 428.400 ;
        RECT 919.950 427.950 922.050 428.400 ;
        RECT 970.950 429.600 973.050 430.050 ;
        RECT 1006.950 429.600 1009.050 430.050 ;
        RECT 970.950 428.400 1009.050 429.600 ;
        RECT 970.950 427.950 973.050 428.400 ;
        RECT 1006.950 427.950 1009.050 428.400 ;
        RECT 61.950 426.600 64.050 427.050 ;
        RECT 121.950 426.600 124.050 427.050 ;
        RECT 130.950 426.600 133.050 427.050 ;
        RECT 163.950 426.600 166.050 427.050 ;
        RECT 61.950 425.400 166.050 426.600 ;
        RECT 61.950 424.950 64.050 425.400 ;
        RECT 121.950 424.950 124.050 425.400 ;
        RECT 130.950 424.950 133.050 425.400 ;
        RECT 163.950 424.950 166.050 425.400 ;
        RECT 214.950 426.600 217.050 427.050 ;
        RECT 241.950 426.600 244.050 427.050 ;
        RECT 253.950 426.600 256.050 427.050 ;
        RECT 214.950 425.400 256.050 426.600 ;
        RECT 214.950 424.950 217.050 425.400 ;
        RECT 241.950 424.950 244.050 425.400 ;
        RECT 253.950 424.950 256.050 425.400 ;
        RECT 289.950 426.600 292.050 427.050 ;
        RECT 334.950 426.600 337.050 427.050 ;
        RECT 289.950 425.400 337.050 426.600 ;
        RECT 289.950 424.950 292.050 425.400 ;
        RECT 334.950 424.950 337.050 425.400 ;
        RECT 388.950 426.600 391.050 427.050 ;
        RECT 400.950 426.600 403.050 427.050 ;
        RECT 388.950 425.400 403.050 426.600 ;
        RECT 388.950 424.950 391.050 425.400 ;
        RECT 400.950 424.950 403.050 425.400 ;
        RECT 415.950 426.600 418.050 427.050 ;
        RECT 421.950 426.600 424.050 427.050 ;
        RECT 415.950 425.400 424.050 426.600 ;
        RECT 415.950 424.950 418.050 425.400 ;
        RECT 421.950 424.950 424.050 425.400 ;
        RECT 436.950 426.600 439.050 427.050 ;
        RECT 460.950 426.600 463.050 427.050 ;
        RECT 436.950 425.400 463.050 426.600 ;
        RECT 436.950 424.950 439.050 425.400 ;
        RECT 460.950 424.950 463.050 425.400 ;
        RECT 475.950 426.600 478.050 427.050 ;
        RECT 520.950 426.600 523.050 427.050 ;
        RECT 535.950 426.600 538.050 427.050 ;
        RECT 568.950 426.600 571.050 427.050 ;
        RECT 664.950 426.600 667.050 427.050 ;
        RECT 475.950 425.400 667.050 426.600 ;
        RECT 475.950 424.950 478.050 425.400 ;
        RECT 520.950 424.950 523.050 425.400 ;
        RECT 535.950 424.950 538.050 425.400 ;
        RECT 568.950 424.950 571.050 425.400 ;
        RECT 664.950 424.950 667.050 425.400 ;
        RECT 691.950 426.600 694.050 427.050 ;
        RECT 700.950 426.600 703.050 427.050 ;
        RECT 691.950 425.400 703.050 426.600 ;
        RECT 691.950 424.950 694.050 425.400 ;
        RECT 700.950 424.950 703.050 425.400 ;
        RECT 766.950 426.600 769.050 427.050 ;
        RECT 775.950 426.600 778.050 427.050 ;
        RECT 766.950 425.400 778.050 426.600 ;
        RECT 766.950 424.950 769.050 425.400 ;
        RECT 775.950 424.950 778.050 425.400 ;
        RECT 820.950 426.600 823.050 427.050 ;
        RECT 829.950 426.600 832.050 427.050 ;
        RECT 820.950 425.400 832.050 426.600 ;
        RECT 820.950 424.950 823.050 425.400 ;
        RECT 829.950 424.950 832.050 425.400 ;
        RECT 904.950 426.600 907.050 427.050 ;
        RECT 910.950 426.600 913.050 427.050 ;
        RECT 904.950 425.400 913.050 426.600 ;
        RECT 904.950 424.950 907.050 425.400 ;
        RECT 910.950 424.950 913.050 425.400 ;
        RECT 943.950 426.600 946.050 427.050 ;
        RECT 958.950 426.600 961.050 427.050 ;
        RECT 943.950 425.400 961.050 426.600 ;
        RECT 943.950 424.950 946.050 425.400 ;
        RECT 958.950 424.950 961.050 425.400 ;
        RECT 13.950 423.600 16.050 424.050 ;
        RECT 28.950 423.600 31.050 424.050 ;
        RECT 13.950 422.400 31.050 423.600 ;
        RECT 13.950 421.950 16.050 422.400 ;
        RECT 28.950 421.950 31.050 422.400 ;
        RECT 139.950 423.600 142.050 424.050 ;
        RECT 145.950 423.600 148.050 424.050 ;
        RECT 139.950 422.400 148.050 423.600 ;
        RECT 139.950 421.950 142.050 422.400 ;
        RECT 145.950 421.950 148.050 422.400 ;
        RECT 175.950 423.600 178.050 424.050 ;
        RECT 235.950 423.600 238.050 424.050 ;
        RECT 175.950 422.400 238.050 423.600 ;
        RECT 175.950 421.950 178.050 422.400 ;
        RECT 235.950 421.950 238.050 422.400 ;
        RECT 253.950 423.600 256.050 423.900 ;
        RECT 259.950 423.600 262.050 424.050 ;
        RECT 325.950 423.600 328.050 424.050 ;
        RECT 253.950 422.400 328.050 423.600 ;
        RECT 253.950 421.800 256.050 422.400 ;
        RECT 259.950 421.950 262.050 422.400 ;
        RECT 325.950 421.950 328.050 422.400 ;
        RECT 427.950 423.600 430.050 424.050 ;
        RECT 469.950 423.600 472.050 424.050 ;
        RECT 427.950 422.400 472.050 423.600 ;
        RECT 427.950 421.950 430.050 422.400 ;
        RECT 469.950 421.950 472.050 422.400 ;
        RECT 478.950 423.600 481.050 424.050 ;
        RECT 502.950 423.600 505.050 424.050 ;
        RECT 478.950 422.400 505.050 423.600 ;
        RECT 478.950 421.950 481.050 422.400 ;
        RECT 502.950 421.950 505.050 422.400 ;
        RECT 571.950 423.600 574.050 424.050 ;
        RECT 625.950 423.600 628.050 424.050 ;
        RECT 571.950 422.400 628.050 423.600 ;
        RECT 571.950 421.950 574.050 422.400 ;
        RECT 625.950 421.950 628.050 422.400 ;
        RECT 715.950 423.600 718.050 424.050 ;
        RECT 724.950 423.600 727.050 424.050 ;
        RECT 763.950 423.600 766.050 424.050 ;
        RECT 715.950 422.400 766.050 423.600 ;
        RECT 715.950 421.950 718.050 422.400 ;
        RECT 724.950 421.950 727.050 422.400 ;
        RECT 763.950 421.950 766.050 422.400 ;
        RECT 847.950 423.600 850.050 424.050 ;
        RECT 871.950 423.600 874.050 423.900 ;
        RECT 847.950 422.400 874.050 423.600 ;
        RECT 847.950 421.950 850.050 422.400 ;
        RECT 871.950 421.800 874.050 422.400 ;
        RECT 892.950 423.600 895.050 424.050 ;
        RECT 916.950 423.600 919.050 424.050 ;
        RECT 892.950 422.400 919.050 423.600 ;
        RECT 892.950 421.950 895.050 422.400 ;
        RECT 916.950 421.950 919.050 422.400 ;
        RECT 928.950 423.600 931.050 424.050 ;
        RECT 970.950 423.600 973.050 424.050 ;
        RECT 928.950 422.400 973.050 423.600 ;
        RECT 928.950 421.950 931.050 422.400 ;
        RECT 970.950 421.950 973.050 422.400 ;
        RECT 232.950 418.950 235.050 421.050 ;
        RECT 553.950 420.600 556.050 421.050 ;
        RECT 565.950 420.600 568.050 421.050 ;
        RECT 553.950 419.400 568.050 420.600 ;
        RECT 553.950 418.950 556.050 419.400 ;
        RECT 565.950 418.950 568.050 419.400 ;
        RECT 652.950 420.600 655.050 421.050 ;
        RECT 673.950 420.600 676.050 421.050 ;
        RECT 652.950 419.400 676.050 420.600 ;
        RECT 652.950 418.950 655.050 419.400 ;
        RECT 673.950 418.950 676.050 419.400 ;
        RECT 679.950 420.600 682.050 421.050 ;
        RECT 685.950 420.600 688.050 421.050 ;
        RECT 679.950 419.400 688.050 420.600 ;
        RECT 679.950 418.950 682.050 419.400 ;
        RECT 685.950 418.950 688.050 419.400 ;
        RECT 769.950 420.600 772.050 421.050 ;
        RECT 784.950 420.600 787.050 421.050 ;
        RECT 769.950 419.400 787.050 420.600 ;
        RECT 769.950 418.950 772.050 419.400 ;
        RECT 784.950 418.950 787.050 419.400 ;
        RECT 862.950 420.600 865.050 421.050 ;
        RECT 925.950 420.600 928.050 421.050 ;
        RECT 862.950 419.400 928.050 420.600 ;
        RECT 862.950 418.950 865.050 419.400 ;
        RECT 925.950 418.950 928.050 419.400 ;
        RECT 16.950 416.100 19.050 418.200 ;
        RECT 22.950 417.750 25.050 418.200 ;
        RECT 31.950 417.750 34.050 418.200 ;
        RECT 22.950 416.550 34.050 417.750 ;
        RECT 22.950 416.100 25.050 416.550 ;
        RECT 31.950 416.100 34.050 416.550 ;
        RECT 40.950 416.100 43.050 418.200 ;
        RECT 46.950 416.100 49.050 418.200 ;
        RECT 115.950 417.600 118.050 418.050 ;
        RECT 127.950 417.750 130.050 418.200 ;
        RECT 136.950 417.750 139.050 418.200 ;
        RECT 127.950 417.600 139.050 417.750 ;
        RECT 115.950 416.550 139.050 417.600 ;
        RECT 115.950 416.400 130.050 416.550 ;
        RECT 17.400 409.050 18.600 416.100 ;
        RECT 41.400 412.050 42.600 416.100 ;
        RECT 47.400 414.600 48.600 416.100 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 127.950 416.100 130.050 416.400 ;
        RECT 136.950 416.100 139.050 416.550 ;
        RECT 148.950 417.750 151.050 418.200 ;
        RECT 157.950 417.750 160.050 418.200 ;
        RECT 148.950 416.550 160.050 417.750 ;
        RECT 148.950 416.100 151.050 416.550 ;
        RECT 157.950 416.100 160.050 416.550 ;
        RECT 217.950 415.950 220.050 418.050 ;
        RECT 223.950 417.600 226.050 417.900 ;
        RECT 229.950 417.600 232.050 418.050 ;
        RECT 223.950 416.400 232.050 417.600 ;
        RECT 58.950 414.600 61.050 415.050 ;
        RECT 37.950 410.400 42.600 412.050 ;
        RECT 44.400 413.400 48.600 414.600 ;
        RECT 50.400 413.400 61.050 414.600 ;
        RECT 37.950 409.950 42.000 410.400 ;
        RECT 44.400 409.050 45.600 413.400 ;
        RECT 50.400 411.900 51.600 413.400 ;
        RECT 58.950 412.950 61.050 413.400 ;
        RECT 79.950 414.450 82.050 414.900 ;
        RECT 103.950 414.450 106.050 414.900 ;
        RECT 79.950 413.250 106.050 414.450 ;
        RECT 79.950 412.800 82.050 413.250 ;
        RECT 103.950 412.800 106.050 413.250 ;
        RECT 218.400 412.050 219.600 415.950 ;
        RECT 223.950 415.800 226.050 416.400 ;
        RECT 229.950 415.950 232.050 416.400 ;
        RECT 49.950 409.800 52.050 411.900 ;
        RECT 139.950 411.600 142.050 411.900 ;
        RECT 145.950 411.600 148.050 412.050 ;
        RECT 139.950 410.400 148.050 411.600 ;
        RECT 139.950 409.800 142.050 410.400 ;
        RECT 145.950 409.950 148.050 410.400 ;
        RECT 160.950 411.600 163.050 411.900 ;
        RECT 187.950 411.600 190.050 411.900 ;
        RECT 211.950 411.600 214.050 411.900 ;
        RECT 160.950 410.400 214.050 411.600 ;
        RECT 160.950 409.800 163.050 410.400 ;
        RECT 187.950 409.800 190.050 410.400 ;
        RECT 211.950 409.800 214.050 410.400 ;
        RECT 217.950 409.950 220.050 412.050 ;
        RECT 233.400 411.900 234.600 418.950 ;
        RECT 265.950 417.750 268.050 418.200 ;
        RECT 274.950 417.750 277.050 418.200 ;
        RECT 265.950 416.550 277.050 417.750 ;
        RECT 265.950 416.100 268.050 416.550 ;
        RECT 274.950 416.100 277.050 416.550 ;
        RECT 292.950 417.750 295.050 418.200 ;
        RECT 319.950 417.750 322.050 418.200 ;
        RECT 292.950 416.550 322.050 417.750 ;
        RECT 292.950 416.100 295.050 416.550 ;
        RECT 319.950 416.100 322.050 416.550 ;
        RECT 331.950 417.600 334.050 418.050 ;
        RECT 373.950 417.600 376.050 418.200 ;
        RECT 331.950 416.400 376.050 417.600 ;
        RECT 331.950 415.950 334.050 416.400 ;
        RECT 373.950 416.100 376.050 416.400 ;
        RECT 421.950 417.750 424.050 418.200 ;
        RECT 430.950 417.750 433.050 418.200 ;
        RECT 421.950 416.550 433.050 417.750 ;
        RECT 421.950 416.100 424.050 416.550 ;
        RECT 430.950 416.100 433.050 416.550 ;
        RECT 448.950 417.750 451.050 418.200 ;
        RECT 457.950 417.750 460.050 418.200 ;
        RECT 448.950 416.550 460.050 417.750 ;
        RECT 448.950 416.100 451.050 416.550 ;
        RECT 457.950 416.100 460.050 416.550 ;
        RECT 496.950 417.750 499.050 418.200 ;
        RECT 520.950 417.750 523.050 418.200 ;
        RECT 496.950 416.550 523.050 417.750 ;
        RECT 496.950 416.100 499.050 416.550 ;
        RECT 520.950 416.100 523.050 416.550 ;
        RECT 529.950 417.750 532.050 418.200 ;
        RECT 541.950 417.750 544.050 418.200 ;
        RECT 529.950 416.550 544.050 417.750 ;
        RECT 529.950 416.100 532.050 416.550 ;
        RECT 541.950 416.100 544.050 416.550 ;
        RECT 559.950 417.600 562.050 418.200 ;
        RECT 574.950 417.600 577.050 418.200 ;
        RECT 559.950 416.400 577.050 417.600 ;
        RECT 559.950 416.100 562.050 416.400 ;
        RECT 572.400 412.050 573.600 416.400 ;
        RECT 574.950 416.100 577.050 416.400 ;
        RECT 586.950 417.600 589.050 418.050 ;
        RECT 607.950 417.600 610.050 418.050 ;
        RECT 586.950 416.400 610.050 417.600 ;
        RECT 586.950 415.950 589.050 416.400 ;
        RECT 607.950 415.950 610.050 416.400 ;
        RECT 625.950 416.100 628.050 418.200 ;
        RECT 643.950 417.600 646.050 418.050 ;
        RECT 694.950 417.600 697.050 418.050 ;
        RECT 643.950 416.400 697.050 417.600 ;
        RECT 626.400 414.600 627.600 416.100 ;
        RECT 643.950 415.950 646.050 416.400 ;
        RECT 694.950 415.950 697.050 416.400 ;
        RECT 703.950 417.750 706.050 418.200 ;
        RECT 712.950 417.750 715.050 418.050 ;
        RECT 733.950 417.750 736.050 418.200 ;
        RECT 703.950 416.550 736.050 417.750 ;
        RECT 703.950 416.100 706.050 416.550 ;
        RECT 712.950 415.950 715.050 416.550 ;
        RECT 733.950 416.100 736.050 416.550 ;
        RECT 757.950 416.100 760.050 418.200 ;
        RECT 766.950 417.600 769.050 418.050 ;
        RECT 799.950 417.600 802.050 418.050 ;
        RECT 766.950 416.400 802.050 417.600 ;
        RECT 637.950 414.600 640.050 415.050 ;
        RECT 626.400 413.400 640.050 414.600 ;
        RECT 637.950 412.950 640.050 413.400 ;
        RECT 232.950 409.800 235.050 411.900 ;
        RECT 238.950 411.600 241.050 411.900 ;
        RECT 250.950 411.600 253.050 412.050 ;
        RECT 262.950 411.600 265.050 411.900 ;
        RECT 238.950 410.400 265.050 411.600 ;
        RECT 238.950 409.800 241.050 410.400 ;
        RECT 250.950 409.950 253.050 410.400 ;
        RECT 262.950 409.800 265.050 410.400 ;
        RECT 274.950 411.600 277.050 412.050 ;
        RECT 286.950 411.600 289.050 411.900 ;
        RECT 274.950 410.400 289.050 411.600 ;
        RECT 274.950 409.950 277.050 410.400 ;
        RECT 286.950 409.800 289.050 410.400 ;
        RECT 298.950 411.450 301.050 411.900 ;
        RECT 304.950 411.450 307.050 411.900 ;
        RECT 352.950 411.600 355.050 411.900 ;
        RECT 298.950 410.250 307.050 411.450 ;
        RECT 298.950 409.800 301.050 410.250 ;
        RECT 304.950 409.800 307.050 410.250 ;
        RECT 344.400 410.400 355.050 411.600 ;
        RECT 16.950 406.950 19.050 409.050 ;
        RECT 40.950 407.400 45.600 409.050 ;
        RECT 58.950 408.600 61.050 409.050 ;
        RECT 64.950 408.600 67.050 409.050 ;
        RECT 58.950 407.400 67.050 408.600 ;
        RECT 40.950 406.950 45.000 407.400 ;
        RECT 58.950 406.950 61.050 407.400 ;
        RECT 64.950 406.950 67.050 407.400 ;
        RECT 331.950 408.600 334.050 409.050 ;
        RECT 344.400 408.600 345.600 410.400 ;
        RECT 352.950 409.800 355.050 410.400 ;
        RECT 385.950 411.450 388.050 411.900 ;
        RECT 397.950 411.450 400.050 411.900 ;
        RECT 385.950 410.250 400.050 411.450 ;
        RECT 385.950 409.800 388.050 410.250 ;
        RECT 397.950 409.800 400.050 410.250 ;
        RECT 418.950 411.450 421.050 411.900 ;
        RECT 433.950 411.450 436.050 411.900 ;
        RECT 418.950 410.250 436.050 411.450 ;
        RECT 418.950 409.800 421.050 410.250 ;
        RECT 433.950 409.800 436.050 410.250 ;
        RECT 442.950 411.600 445.050 412.050 ;
        RECT 466.950 411.600 469.050 412.050 ;
        RECT 475.950 411.600 478.050 411.900 ;
        RECT 442.950 410.400 478.050 411.600 ;
        RECT 442.950 409.950 445.050 410.400 ;
        RECT 466.950 409.950 469.050 410.400 ;
        RECT 475.950 409.800 478.050 410.400 ;
        RECT 571.950 409.950 574.050 412.050 ;
        RECT 628.950 411.600 631.050 411.900 ;
        RECT 649.950 411.600 652.050 411.900 ;
        RECT 628.950 410.400 652.050 411.600 ;
        RECT 628.950 409.800 631.050 410.400 ;
        RECT 649.950 409.800 652.050 410.400 ;
        RECT 676.950 411.450 679.050 411.900 ;
        RECT 691.950 411.450 694.050 411.900 ;
        RECT 676.950 410.250 694.050 411.450 ;
        RECT 676.950 409.800 679.050 410.250 ;
        RECT 691.950 409.800 694.050 410.250 ;
        RECT 700.950 411.600 703.050 411.900 ;
        RECT 706.950 411.600 709.050 412.050 ;
        RECT 700.950 410.400 709.050 411.600 ;
        RECT 700.950 409.800 703.050 410.400 ;
        RECT 706.950 409.950 709.050 410.400 ;
        RECT 712.950 411.450 715.050 411.900 ;
        RECT 718.950 411.450 721.050 411.900 ;
        RECT 712.950 410.250 721.050 411.450 ;
        RECT 712.950 409.800 715.050 410.250 ;
        RECT 718.950 409.800 721.050 410.250 ;
        RECT 748.950 411.600 751.050 412.050 ;
        RECT 758.400 411.600 759.600 416.100 ;
        RECT 766.950 415.950 769.050 416.400 ;
        RECT 799.950 415.950 802.050 416.400 ;
        RECT 817.950 417.600 820.050 418.050 ;
        RECT 823.950 417.600 826.050 418.200 ;
        RECT 835.950 417.600 838.050 418.050 ;
        RECT 817.950 416.400 826.050 417.600 ;
        RECT 817.950 415.950 820.050 416.400 ;
        RECT 823.950 416.100 826.050 416.400 ;
        RECT 827.400 416.400 838.050 417.600 ;
        RECT 827.400 414.600 828.600 416.400 ;
        RECT 835.950 415.950 838.050 416.400 ;
        RECT 853.950 416.100 856.050 418.200 ;
        RECT 910.950 416.100 913.050 418.200 ;
        RECT 809.400 413.400 828.600 414.600 ;
        RECT 854.400 414.600 855.600 416.100 ;
        RECT 907.950 414.600 910.050 415.050 ;
        RECT 854.400 413.400 910.050 414.600 ;
        RECT 911.400 414.600 912.600 416.100 ;
        RECT 940.950 415.950 943.050 418.050 ;
        RECT 946.950 416.100 949.050 418.200 ;
        RECT 970.950 417.600 973.050 418.200 ;
        RECT 991.950 417.600 994.050 418.200 ;
        RECT 970.950 416.400 994.050 417.600 ;
        RECT 970.950 416.100 973.050 416.400 ;
        RECT 991.950 416.100 994.050 416.400 ;
        RECT 1018.950 416.100 1021.050 418.200 ;
        RECT 928.950 414.600 931.050 415.050 ;
        RECT 911.400 413.400 931.050 414.600 ;
        RECT 748.950 410.400 759.600 411.600 ;
        RECT 763.950 411.450 766.050 411.900 ;
        RECT 772.950 411.450 775.050 412.050 ;
        RECT 778.950 411.450 781.050 411.900 ;
        RECT 748.950 409.950 751.050 410.400 ;
        RECT 763.950 410.250 781.050 411.450 ;
        RECT 763.950 409.800 766.050 410.250 ;
        RECT 772.950 409.950 775.050 410.250 ;
        RECT 778.950 409.800 781.050 410.250 ;
        RECT 805.950 411.600 808.050 411.900 ;
        RECT 809.400 411.600 810.600 413.400 ;
        RECT 907.950 412.950 910.050 413.400 ;
        RECT 928.950 412.950 931.050 413.400 ;
        RECT 941.400 412.050 942.600 415.950 ;
        RECT 805.950 410.400 810.600 411.600 ;
        RECT 832.950 411.450 835.050 411.900 ;
        RECT 841.950 411.450 844.050 411.900 ;
        RECT 805.950 409.800 808.050 410.400 ;
        RECT 832.950 410.250 844.050 411.450 ;
        RECT 832.950 409.800 835.050 410.250 ;
        RECT 841.950 409.800 844.050 410.250 ;
        RECT 889.950 411.600 892.050 411.900 ;
        RECT 895.950 411.600 898.050 412.050 ;
        RECT 889.950 410.400 898.050 411.600 ;
        RECT 889.950 409.800 892.050 410.400 ;
        RECT 895.950 409.950 898.050 410.400 ;
        RECT 940.950 409.950 943.050 412.050 ;
        RECT 947.400 411.600 948.600 416.100 ;
        RECT 955.950 411.600 958.050 412.050 ;
        RECT 1015.950 411.600 1018.050 411.900 ;
        RECT 947.400 410.400 954.600 411.600 ;
        RECT 331.950 407.400 345.600 408.600 ;
        RECT 568.950 408.600 571.050 409.050 ;
        RECT 577.950 408.600 580.050 409.050 ;
        RECT 568.950 407.400 580.050 408.600 ;
        RECT 331.950 406.950 334.050 407.400 ;
        RECT 568.950 406.950 571.050 407.400 ;
        RECT 577.950 406.950 580.050 407.400 ;
        RECT 757.950 408.600 760.050 409.050 ;
        RECT 766.950 408.600 769.050 409.050 ;
        RECT 757.950 407.400 769.050 408.600 ;
        RECT 757.950 406.950 760.050 407.400 ;
        RECT 766.950 406.950 769.050 407.400 ;
        RECT 850.950 408.600 853.050 409.050 ;
        RECT 880.950 408.600 883.050 409.050 ;
        RECT 850.950 407.400 883.050 408.600 ;
        RECT 953.400 408.600 954.600 410.400 ;
        RECT 955.950 410.400 1018.050 411.600 ;
        RECT 955.950 409.950 958.050 410.400 ;
        RECT 1015.950 409.800 1018.050 410.400 ;
        RECT 973.950 408.600 976.050 409.050 ;
        RECT 988.950 408.600 991.050 409.050 ;
        RECT 1019.400 408.600 1020.600 416.100 ;
        RECT 1024.950 415.950 1027.050 418.050 ;
        RECT 1025.400 412.050 1026.600 415.950 ;
        RECT 1024.950 409.950 1027.050 412.050 ;
        RECT 953.400 407.400 1020.600 408.600 ;
        RECT 850.950 406.950 853.050 407.400 ;
        RECT 880.950 406.950 883.050 407.400 ;
        RECT 973.950 406.950 976.050 407.400 ;
        RECT 988.950 406.950 991.050 407.400 ;
        RECT 10.950 405.600 13.050 406.050 ;
        RECT 19.950 405.600 22.050 406.050 ;
        RECT 10.950 404.400 22.050 405.600 ;
        RECT 10.950 403.950 13.050 404.400 ;
        RECT 19.950 403.950 22.050 404.400 ;
        RECT 28.950 405.600 31.050 406.050 ;
        RECT 55.950 405.600 58.050 406.050 ;
        RECT 28.950 404.400 58.050 405.600 ;
        RECT 28.950 403.950 31.050 404.400 ;
        RECT 55.950 403.950 58.050 404.400 ;
        RECT 190.950 405.600 193.050 406.050 ;
        RECT 253.950 405.600 256.050 406.050 ;
        RECT 190.950 404.400 256.050 405.600 ;
        RECT 190.950 403.950 193.050 404.400 ;
        RECT 253.950 403.950 256.050 404.400 ;
        RECT 274.950 405.600 277.050 406.050 ;
        RECT 298.950 405.600 301.050 406.050 ;
        RECT 274.950 404.400 301.050 405.600 ;
        RECT 274.950 403.950 277.050 404.400 ;
        RECT 298.950 403.950 301.050 404.400 ;
        RECT 334.950 405.600 337.050 406.050 ;
        RECT 403.950 405.600 406.050 406.050 ;
        RECT 334.950 404.400 406.050 405.600 ;
        RECT 334.950 403.950 337.050 404.400 ;
        RECT 403.950 403.950 406.050 404.400 ;
        RECT 541.950 405.600 544.050 406.050 ;
        RECT 700.950 405.600 703.050 406.050 ;
        RECT 541.950 404.400 703.050 405.600 ;
        RECT 541.950 403.950 544.050 404.400 ;
        RECT 700.950 403.950 703.050 404.400 ;
        RECT 928.950 405.600 931.050 406.050 ;
        RECT 955.950 405.600 958.050 406.050 ;
        RECT 928.950 404.400 958.050 405.600 ;
        RECT 928.950 403.950 931.050 404.400 ;
        RECT 955.950 403.950 958.050 404.400 ;
        RECT 994.950 405.600 997.050 406.050 ;
        RECT 1009.950 405.600 1012.050 406.050 ;
        RECT 1021.950 405.600 1024.050 406.050 ;
        RECT 994.950 404.400 1024.050 405.600 ;
        RECT 994.950 403.950 997.050 404.400 ;
        RECT 1009.950 403.950 1012.050 404.400 ;
        RECT 1021.950 403.950 1024.050 404.400 ;
        RECT 265.950 402.600 268.050 403.050 ;
        RECT 271.950 402.600 274.050 403.050 ;
        RECT 265.950 401.400 274.050 402.600 ;
        RECT 265.950 400.950 268.050 401.400 ;
        RECT 271.950 400.950 274.050 401.400 ;
        RECT 565.950 402.600 568.050 403.050 ;
        RECT 595.950 402.600 598.050 403.050 ;
        RECT 643.950 402.600 646.050 403.050 ;
        RECT 757.950 402.600 760.050 403.050 ;
        RECT 565.950 401.400 760.050 402.600 ;
        RECT 565.950 400.950 568.050 401.400 ;
        RECT 595.950 400.950 598.050 401.400 ;
        RECT 643.950 400.950 646.050 401.400 ;
        RECT 757.950 400.950 760.050 401.400 ;
        RECT 763.950 402.600 766.050 403.050 ;
        RECT 784.950 402.600 787.050 403.050 ;
        RECT 829.950 402.600 832.050 403.050 ;
        RECT 763.950 401.400 832.050 402.600 ;
        RECT 763.950 400.950 766.050 401.400 ;
        RECT 784.950 400.950 787.050 401.400 ;
        RECT 829.950 400.950 832.050 401.400 ;
        RECT 871.950 402.600 874.050 403.050 ;
        RECT 919.950 402.600 922.050 403.050 ;
        RECT 871.950 401.400 922.050 402.600 ;
        RECT 871.950 400.950 874.050 401.400 ;
        RECT 919.950 400.950 922.050 401.400 ;
        RECT 961.950 402.600 964.050 403.050 ;
        RECT 1030.950 402.600 1033.050 403.050 ;
        RECT 961.950 401.400 1033.050 402.600 ;
        RECT 961.950 400.950 964.050 401.400 ;
        RECT 1030.950 400.950 1033.050 401.400 ;
        RECT 16.950 399.600 19.050 400.050 ;
        RECT 25.950 399.600 28.050 400.050 ;
        RECT 16.950 398.400 28.050 399.600 ;
        RECT 16.950 397.950 19.050 398.400 ;
        RECT 25.950 397.950 28.050 398.400 ;
        RECT 184.950 399.600 187.050 400.050 ;
        RECT 232.950 399.600 235.050 400.050 ;
        RECT 184.950 398.400 235.050 399.600 ;
        RECT 184.950 397.950 187.050 398.400 ;
        RECT 232.950 397.950 235.050 398.400 ;
        RECT 286.950 399.600 289.050 400.050 ;
        RECT 301.950 399.600 304.050 400.050 ;
        RECT 349.950 399.600 352.050 400.050 ;
        RECT 370.950 399.600 373.050 400.050 ;
        RECT 286.950 398.400 373.050 399.600 ;
        RECT 286.950 397.950 289.050 398.400 ;
        RECT 301.950 397.950 304.050 398.400 ;
        RECT 349.950 397.950 352.050 398.400 ;
        RECT 370.950 397.950 373.050 398.400 ;
        RECT 430.950 399.600 433.050 400.050 ;
        RECT 463.950 399.600 466.050 400.050 ;
        RECT 586.950 399.600 589.050 400.050 ;
        RECT 430.950 398.400 589.050 399.600 ;
        RECT 430.950 397.950 433.050 398.400 ;
        RECT 463.950 397.950 466.050 398.400 ;
        RECT 586.950 397.950 589.050 398.400 ;
        RECT 637.950 399.600 640.050 400.050 ;
        RECT 655.950 399.600 658.050 400.050 ;
        RECT 637.950 398.400 658.050 399.600 ;
        RECT 637.950 397.950 640.050 398.400 ;
        RECT 655.950 397.950 658.050 398.400 ;
        RECT 682.950 399.600 685.050 400.050 ;
        RECT 712.950 399.600 715.050 400.050 ;
        RECT 682.950 398.400 715.050 399.600 ;
        RECT 682.950 397.950 685.050 398.400 ;
        RECT 712.950 397.950 715.050 398.400 ;
        RECT 718.950 399.600 721.050 400.050 ;
        RECT 736.950 399.600 739.050 400.050 ;
        RECT 718.950 398.400 739.050 399.600 ;
        RECT 718.950 397.950 721.050 398.400 ;
        RECT 736.950 397.950 739.050 398.400 ;
        RECT 874.950 399.600 877.050 400.050 ;
        RECT 889.800 399.600 891.900 400.050 ;
        RECT 874.950 398.400 891.900 399.600 ;
        RECT 874.950 397.950 877.050 398.400 ;
        RECT 889.800 397.950 891.900 398.400 ;
        RECT 892.950 399.600 895.050 400.050 ;
        RECT 943.950 399.600 946.050 400.050 ;
        RECT 892.950 398.400 946.050 399.600 ;
        RECT 892.950 397.950 895.050 398.400 ;
        RECT 943.950 397.950 946.050 398.400 ;
        RECT 949.950 399.600 952.050 400.050 ;
        RECT 1042.950 399.600 1045.050 400.050 ;
        RECT 949.950 398.400 1045.050 399.600 ;
        RECT 949.950 397.950 952.050 398.400 ;
        RECT 1042.950 397.950 1045.050 398.400 ;
        RECT 31.950 396.600 34.050 397.050 ;
        RECT 127.950 396.600 130.050 397.050 ;
        RECT 31.950 395.400 130.050 396.600 ;
        RECT 31.950 394.950 34.050 395.400 ;
        RECT 127.950 394.950 130.050 395.400 ;
        RECT 250.950 396.600 253.050 397.050 ;
        RECT 292.950 396.600 295.050 397.050 ;
        RECT 250.950 395.400 295.050 396.600 ;
        RECT 250.950 394.950 253.050 395.400 ;
        RECT 292.950 394.950 295.050 395.400 ;
        RECT 304.950 396.600 307.050 397.050 ;
        RECT 331.950 396.600 334.050 397.050 ;
        RECT 304.950 395.400 334.050 396.600 ;
        RECT 304.950 394.950 307.050 395.400 ;
        RECT 331.950 394.950 334.050 395.400 ;
        RECT 739.950 396.600 742.050 397.050 ;
        RECT 793.950 396.600 796.050 397.050 ;
        RECT 739.950 395.400 796.050 396.600 ;
        RECT 739.950 394.950 742.050 395.400 ;
        RECT 793.950 394.950 796.050 395.400 ;
        RECT 802.950 396.600 805.050 397.050 ;
        RECT 814.950 396.600 817.050 397.050 ;
        RECT 913.950 396.600 916.050 397.050 ;
        RECT 976.950 396.600 979.050 397.050 ;
        RECT 802.950 395.400 817.050 396.600 ;
        RECT 802.950 394.950 805.050 395.400 ;
        RECT 814.950 394.950 817.050 395.400 ;
        RECT 878.400 395.400 885.600 396.600 ;
        RECT 43.950 393.600 46.050 394.050 ;
        RECT 169.950 393.600 172.050 394.050 ;
        RECT 43.950 392.400 172.050 393.600 ;
        RECT 43.950 391.950 46.050 392.400 ;
        RECT 169.950 391.950 172.050 392.400 ;
        RECT 571.950 393.600 574.050 394.050 ;
        RECT 748.950 393.600 751.050 394.050 ;
        RECT 790.950 393.600 793.050 394.050 ;
        RECT 571.950 392.400 751.050 393.600 ;
        RECT 571.950 391.950 574.050 392.400 ;
        RECT 748.950 391.950 751.050 392.400 ;
        RECT 764.400 392.400 793.050 393.600 ;
        RECT 67.950 390.600 70.050 391.050 ;
        RECT 181.950 390.600 184.050 391.050 ;
        RECT 67.950 389.400 184.050 390.600 ;
        RECT 67.950 388.950 70.050 389.400 ;
        RECT 181.950 388.950 184.050 389.400 ;
        RECT 247.950 390.600 250.050 391.050 ;
        RECT 376.950 390.600 379.050 391.050 ;
        RECT 247.950 389.400 379.050 390.600 ;
        RECT 247.950 388.950 250.050 389.400 ;
        RECT 376.950 388.950 379.050 389.400 ;
        RECT 508.950 390.600 511.050 391.050 ;
        RECT 556.950 390.600 559.050 391.050 ;
        RECT 508.950 389.400 559.050 390.600 ;
        RECT 508.950 388.950 511.050 389.400 ;
        RECT 556.950 388.950 559.050 389.400 ;
        RECT 574.950 390.600 577.050 391.050 ;
        RECT 601.950 390.600 604.050 391.050 ;
        RECT 574.950 389.400 604.050 390.600 ;
        RECT 574.950 388.950 577.050 389.400 ;
        RECT 601.950 388.950 604.050 389.400 ;
        RECT 643.950 390.600 646.050 391.050 ;
        RECT 682.950 390.600 685.050 391.050 ;
        RECT 643.950 389.400 685.050 390.600 ;
        RECT 643.950 388.950 646.050 389.400 ;
        RECT 682.950 388.950 685.050 389.400 ;
        RECT 688.950 390.600 691.050 391.050 ;
        RECT 709.950 390.600 712.050 391.050 ;
        RECT 688.950 389.400 712.050 390.600 ;
        RECT 688.950 388.950 691.050 389.400 ;
        RECT 709.950 388.950 712.050 389.400 ;
        RECT 727.950 390.600 730.050 391.050 ;
        RECT 764.400 390.600 765.600 392.400 ;
        RECT 790.950 391.950 793.050 392.400 ;
        RECT 826.950 393.600 829.050 394.050 ;
        RECT 878.400 393.600 879.600 395.400 ;
        RECT 826.950 392.400 879.600 393.600 ;
        RECT 884.400 393.600 885.600 395.400 ;
        RECT 913.950 395.400 979.050 396.600 ;
        RECT 913.950 394.950 916.050 395.400 ;
        RECT 976.950 394.950 979.050 395.400 ;
        RECT 991.950 396.600 994.050 397.050 ;
        RECT 1015.950 396.600 1018.050 397.050 ;
        RECT 991.950 395.400 1018.050 396.600 ;
        RECT 991.950 394.950 994.050 395.400 ;
        RECT 1015.950 394.950 1018.050 395.400 ;
        RECT 892.950 393.600 895.050 394.050 ;
        RECT 884.400 392.400 895.050 393.600 ;
        RECT 826.950 391.950 829.050 392.400 ;
        RECT 892.950 391.950 895.050 392.400 ;
        RECT 943.950 393.600 946.050 394.050 ;
        RECT 958.950 393.600 961.050 394.050 ;
        RECT 1024.950 393.600 1027.050 394.050 ;
        RECT 943.950 392.400 961.050 393.600 ;
        RECT 943.950 391.950 946.050 392.400 ;
        RECT 958.950 391.950 961.050 392.400 ;
        RECT 980.400 392.400 1027.050 393.600 ;
        RECT 727.950 389.400 765.600 390.600 ;
        RECT 811.950 390.600 814.050 391.050 ;
        RECT 817.950 390.600 820.050 391.050 ;
        RECT 811.950 389.400 820.050 390.600 ;
        RECT 727.950 388.950 730.050 389.400 ;
        RECT 811.950 388.950 814.050 389.400 ;
        RECT 817.950 388.950 820.050 389.400 ;
        RECT 880.950 390.600 883.050 391.050 ;
        RECT 907.950 390.600 910.050 391.050 ;
        RECT 880.950 389.400 910.050 390.600 ;
        RECT 880.950 388.950 883.050 389.400 ;
        RECT 907.950 388.950 910.050 389.400 ;
        RECT 922.950 390.600 925.050 391.050 ;
        RECT 980.400 390.600 981.600 392.400 ;
        RECT 1024.950 391.950 1027.050 392.400 ;
        RECT 922.950 389.400 981.600 390.600 ;
        RECT 922.950 388.950 925.050 389.400 ;
        RECT 103.950 387.600 106.050 388.050 ;
        RECT 148.950 387.600 151.050 388.050 ;
        RECT 103.950 386.400 151.050 387.600 ;
        RECT 103.950 385.950 106.050 386.400 ;
        RECT 148.950 385.950 151.050 386.400 ;
        RECT 439.950 387.600 442.050 388.050 ;
        RECT 547.950 387.600 550.050 388.050 ;
        RECT 439.950 386.400 550.050 387.600 ;
        RECT 439.950 385.950 442.050 386.400 ;
        RECT 547.950 385.950 550.050 386.400 ;
        RECT 565.950 387.600 568.050 388.050 ;
        RECT 571.950 387.600 574.050 388.050 ;
        RECT 565.950 386.400 574.050 387.600 ;
        RECT 565.950 385.950 568.050 386.400 ;
        RECT 571.950 385.950 574.050 386.400 ;
        RECT 583.950 387.600 586.050 388.050 ;
        RECT 592.950 387.600 595.050 388.050 ;
        RECT 583.950 386.400 595.050 387.600 ;
        RECT 583.950 385.950 586.050 386.400 ;
        RECT 592.950 385.950 595.050 386.400 ;
        RECT 661.950 387.600 664.050 388.050 ;
        RECT 781.950 387.600 784.050 388.050 ;
        RECT 661.950 386.400 784.050 387.600 ;
        RECT 661.950 385.950 664.050 386.400 ;
        RECT 781.950 385.950 784.050 386.400 ;
        RECT 805.950 387.600 808.050 388.050 ;
        RECT 859.950 387.600 862.050 388.050 ;
        RECT 805.950 386.400 862.050 387.600 ;
        RECT 805.950 385.950 808.050 386.400 ;
        RECT 859.950 385.950 862.050 386.400 ;
        RECT 910.950 387.600 913.050 388.050 ;
        RECT 988.950 387.600 991.050 388.050 ;
        RECT 910.950 386.400 991.050 387.600 ;
        RECT 910.950 385.950 913.050 386.400 ;
        RECT 988.950 385.950 991.050 386.400 ;
        RECT 142.950 384.600 145.050 385.050 ;
        RECT 187.950 384.600 190.050 385.050 ;
        RECT 142.950 383.400 190.050 384.600 ;
        RECT 142.950 382.950 145.050 383.400 ;
        RECT 187.950 382.950 190.050 383.400 ;
        RECT 358.950 384.600 361.050 385.050 ;
        RECT 421.950 384.600 424.050 385.050 ;
        RECT 358.950 383.400 424.050 384.600 ;
        RECT 358.950 382.950 361.050 383.400 ;
        RECT 421.950 382.950 424.050 383.400 ;
        RECT 574.950 384.600 577.050 385.050 ;
        RECT 622.950 384.600 625.050 385.050 ;
        RECT 574.950 383.400 625.050 384.600 ;
        RECT 574.950 382.950 577.050 383.400 ;
        RECT 622.950 382.950 625.050 383.400 ;
        RECT 694.950 384.600 697.050 385.050 ;
        RECT 703.950 384.600 706.050 385.050 ;
        RECT 694.950 383.400 706.050 384.600 ;
        RECT 694.950 382.950 697.050 383.400 ;
        RECT 703.950 382.950 706.050 383.400 ;
        RECT 862.950 384.600 865.050 385.050 ;
        RECT 880.950 384.600 883.050 385.050 ;
        RECT 862.950 383.400 883.050 384.600 ;
        RECT 862.950 382.950 865.050 383.400 ;
        RECT 880.950 382.950 883.050 383.400 ;
        RECT 931.950 384.600 934.050 385.050 ;
        RECT 955.950 384.600 958.050 385.050 ;
        RECT 931.950 383.400 958.050 384.600 ;
        RECT 931.950 382.950 934.050 383.400 ;
        RECT 955.950 382.950 958.050 383.400 ;
        RECT 970.950 384.600 973.050 385.050 ;
        RECT 1036.950 384.600 1039.050 385.050 ;
        RECT 970.950 383.400 1039.050 384.600 ;
        RECT 970.950 382.950 973.050 383.400 ;
        RECT 1036.950 382.950 1039.050 383.400 ;
        RECT 118.950 381.600 121.050 382.050 ;
        RECT 47.400 380.400 121.050 381.600 ;
        RECT 47.400 379.050 48.600 380.400 ;
        RECT 118.950 379.950 121.050 380.400 ;
        RECT 211.950 381.600 214.050 382.050 ;
        RECT 250.950 381.600 253.050 382.050 ;
        RECT 211.950 380.400 253.050 381.600 ;
        RECT 211.950 379.950 214.050 380.400 ;
        RECT 250.950 379.950 253.050 380.400 ;
        RECT 286.950 381.600 289.050 382.050 ;
        RECT 304.950 381.600 307.050 382.050 ;
        RECT 286.950 380.400 307.050 381.600 ;
        RECT 286.950 379.950 289.050 380.400 ;
        RECT 304.950 379.950 307.050 380.400 ;
        RECT 310.950 381.600 313.050 382.050 ;
        RECT 322.950 381.600 325.050 382.050 ;
        RECT 310.950 380.400 325.050 381.600 ;
        RECT 310.950 379.950 313.050 380.400 ;
        RECT 322.950 379.950 325.050 380.400 ;
        RECT 745.950 381.600 748.050 382.050 ;
        RECT 769.950 381.600 772.050 382.050 ;
        RECT 745.950 380.400 772.050 381.600 ;
        RECT 745.950 379.950 748.050 380.400 ;
        RECT 769.950 379.950 772.050 380.400 ;
        RECT 823.950 381.600 826.050 382.050 ;
        RECT 838.950 381.600 841.050 382.050 ;
        RECT 823.950 380.400 841.050 381.600 ;
        RECT 823.950 379.950 826.050 380.400 ;
        RECT 838.950 379.950 841.050 380.400 ;
        RECT 910.950 381.600 913.050 382.050 ;
        RECT 979.950 381.600 982.050 382.050 ;
        RECT 910.950 380.400 982.050 381.600 ;
        RECT 910.950 379.950 913.050 380.400 ;
        RECT 979.950 379.950 982.050 380.400 ;
        RECT 16.950 378.600 19.050 379.050 ;
        RECT 37.950 378.600 40.050 379.050 ;
        RECT 46.950 378.600 49.050 379.050 ;
        RECT 265.950 378.600 268.050 379.050 ;
        RECT 16.950 377.400 49.050 378.600 ;
        RECT 16.950 376.950 19.050 377.400 ;
        RECT 37.950 376.950 40.050 377.400 ;
        RECT 46.950 376.950 49.050 377.400 ;
        RECT 257.400 377.400 268.050 378.600 ;
        RECT 235.950 375.600 238.050 376.050 ;
        RECT 257.400 375.600 258.600 377.400 ;
        RECT 265.950 376.950 268.050 377.400 ;
        RECT 271.950 378.600 274.050 379.050 ;
        RECT 355.950 378.600 358.050 379.050 ;
        RECT 271.950 377.400 358.050 378.600 ;
        RECT 271.950 376.950 274.050 377.400 ;
        RECT 355.950 376.950 358.050 377.400 ;
        RECT 379.950 378.600 382.050 379.050 ;
        RECT 439.950 378.600 442.050 379.050 ;
        RECT 379.950 377.400 442.050 378.600 ;
        RECT 379.950 376.950 382.050 377.400 ;
        RECT 439.950 376.950 442.050 377.400 ;
        RECT 463.950 378.600 466.050 379.050 ;
        RECT 532.950 378.600 535.050 379.050 ;
        RECT 463.950 377.400 535.050 378.600 ;
        RECT 463.950 376.950 466.050 377.400 ;
        RECT 532.950 376.950 535.050 377.400 ;
        RECT 586.950 378.600 589.050 379.050 ;
        RECT 661.950 378.600 664.050 379.050 ;
        RECT 586.950 377.400 664.050 378.600 ;
        RECT 586.950 376.950 589.050 377.400 ;
        RECT 661.950 376.950 664.050 377.400 ;
        RECT 676.950 378.600 679.050 379.050 ;
        RECT 682.950 378.600 685.050 379.050 ;
        RECT 721.950 378.600 724.050 379.050 ;
        RECT 676.950 377.400 724.050 378.600 ;
        RECT 676.950 376.950 679.050 377.400 ;
        RECT 682.950 376.950 685.050 377.400 ;
        RECT 721.950 376.950 724.050 377.400 ;
        RECT 805.950 378.600 808.050 379.050 ;
        RECT 820.950 378.600 823.050 379.050 ;
        RECT 805.950 377.400 823.050 378.600 ;
        RECT 805.950 376.950 808.050 377.400 ;
        RECT 820.950 376.950 823.050 377.400 ;
        RECT 844.950 378.600 847.050 379.050 ;
        RECT 856.950 378.600 859.050 379.050 ;
        RECT 844.950 377.400 859.050 378.600 ;
        RECT 844.950 376.950 847.050 377.400 ;
        RECT 856.950 376.950 859.050 377.400 ;
        RECT 919.950 378.600 922.050 379.050 ;
        RECT 931.950 378.600 934.050 379.050 ;
        RECT 919.950 377.400 934.050 378.600 ;
        RECT 919.950 376.950 922.050 377.400 ;
        RECT 931.950 376.950 934.050 377.400 ;
        RECT 967.950 378.600 970.050 379.050 ;
        RECT 976.950 378.600 979.050 379.050 ;
        RECT 967.950 377.400 979.050 378.600 ;
        RECT 967.950 376.950 970.050 377.400 ;
        RECT 976.950 376.950 979.050 377.400 ;
        RECT 1012.950 378.600 1015.050 379.050 ;
        RECT 1024.950 378.600 1027.050 379.050 ;
        RECT 1012.950 377.400 1027.050 378.600 ;
        RECT 1012.950 376.950 1015.050 377.400 ;
        RECT 1024.950 376.950 1027.050 377.400 ;
        RECT 235.950 374.400 258.600 375.600 ;
        RECT 316.950 375.600 319.050 376.050 ;
        RECT 358.950 375.600 361.050 376.050 ;
        RECT 316.950 374.400 361.050 375.600 ;
        RECT 235.950 373.950 238.050 374.400 ;
        RECT 316.950 373.950 319.050 374.400 ;
        RECT 358.950 373.950 361.050 374.400 ;
        RECT 370.950 375.600 373.050 376.050 ;
        RECT 448.950 375.600 451.050 376.050 ;
        RECT 547.950 375.600 550.050 376.050 ;
        RECT 574.950 375.600 577.050 376.050 ;
        RECT 370.950 374.400 451.050 375.600 ;
        RECT 370.950 373.950 373.050 374.400 ;
        RECT 448.950 373.950 451.050 374.400 ;
        RECT 524.400 374.400 577.050 375.600 ;
        RECT 79.950 372.600 82.050 373.050 ;
        RECT 112.950 372.600 115.050 373.200 ;
        RECT 79.950 371.400 115.050 372.600 ;
        RECT 79.950 370.950 82.050 371.400 ;
        RECT 112.950 371.100 115.050 371.400 ;
        RECT 157.950 372.750 160.050 373.200 ;
        RECT 163.950 372.750 166.050 373.200 ;
        RECT 157.950 371.550 166.050 372.750 ;
        RECT 157.950 371.100 160.050 371.550 ;
        RECT 163.950 371.100 166.050 371.550 ;
        RECT 184.950 372.600 187.050 373.050 ;
        RECT 223.950 372.600 226.050 373.050 ;
        RECT 184.950 371.400 226.050 372.600 ;
        RECT 184.950 370.950 187.050 371.400 ;
        RECT 223.950 370.950 226.050 371.400 ;
        RECT 229.950 370.950 232.050 373.050 ;
        RECT 241.950 371.100 244.050 373.200 ;
        RECT 250.950 372.750 253.050 373.200 ;
        RECT 259.950 372.750 262.050 373.200 ;
        RECT 250.950 371.550 262.050 372.750 ;
        RECT 250.950 371.100 253.050 371.550 ;
        RECT 259.950 371.100 262.050 371.550 ;
        RECT 230.400 367.050 231.600 370.950 ;
        RECT 242.400 367.050 243.600 371.100 ;
        RECT 295.950 370.950 298.050 373.050 ;
        RECT 328.950 372.750 331.050 373.200 ;
        RECT 340.950 372.750 343.050 373.200 ;
        RECT 328.950 371.550 343.050 372.750 ;
        RECT 328.950 371.100 331.050 371.550 ;
        RECT 340.950 371.100 343.050 371.550 ;
        RECT 400.950 372.600 403.050 373.200 ;
        RECT 430.950 372.600 433.050 373.200 ;
        RECT 400.950 371.400 433.050 372.600 ;
        RECT 400.950 371.100 403.050 371.400 ;
        RECT 430.950 371.100 433.050 371.400 ;
        RECT 436.950 372.750 439.050 373.200 ;
        RECT 445.950 372.750 448.050 373.200 ;
        RECT 436.950 371.550 448.050 372.750 ;
        RECT 436.950 371.100 439.050 371.550 ;
        RECT 445.950 371.100 448.050 371.550 ;
        RECT 454.950 372.600 457.050 373.200 ;
        RECT 475.950 372.600 478.050 373.200 ;
        RECT 454.950 371.400 478.050 372.600 ;
        RECT 454.950 371.100 457.050 371.400 ;
        RECT 475.950 371.100 478.050 371.400 ;
        RECT 481.950 372.600 484.050 373.200 ;
        RECT 499.950 372.600 502.050 373.200 ;
        RECT 520.950 372.600 523.050 373.200 ;
        RECT 481.950 371.400 523.050 372.600 ;
        RECT 481.950 371.100 484.050 371.400 ;
        RECT 499.950 371.100 502.050 371.400 ;
        RECT 520.950 371.100 523.050 371.400 ;
        RECT 247.950 369.600 250.050 370.050 ;
        RECT 271.950 369.600 274.050 370.050 ;
        RECT 247.950 368.400 274.050 369.600 ;
        RECT 247.950 367.950 250.050 368.400 ;
        RECT 271.950 367.950 274.050 368.400 ;
        RECT 43.950 366.450 46.050 366.900 ;
        RECT 52.950 366.450 55.050 366.900 ;
        RECT 43.950 365.250 55.050 366.450 ;
        RECT 43.950 364.800 46.050 365.250 ;
        RECT 52.950 364.800 55.050 365.250 ;
        RECT 73.950 366.600 76.050 367.050 ;
        RECT 88.950 366.600 91.050 366.900 ;
        RECT 103.950 366.600 106.050 367.050 ;
        RECT 73.950 365.400 106.050 366.600 ;
        RECT 73.950 364.950 76.050 365.400 ;
        RECT 88.950 364.800 91.050 365.400 ;
        RECT 103.950 364.950 106.050 365.400 ;
        RECT 121.950 366.600 124.050 366.900 ;
        RECT 145.950 366.600 148.050 366.900 ;
        RECT 121.950 365.400 148.050 366.600 ;
        RECT 121.950 364.800 124.050 365.400 ;
        RECT 145.950 364.800 148.050 365.400 ;
        RECT 172.950 366.450 175.050 366.900 ;
        RECT 184.950 366.450 187.050 366.900 ;
        RECT 172.950 365.250 187.050 366.450 ;
        RECT 172.950 364.800 175.050 365.250 ;
        RECT 184.950 364.800 187.050 365.250 ;
        RECT 229.950 364.950 232.050 367.050 ;
        RECT 242.400 365.400 247.050 367.050 ;
        RECT 243.000 364.950 247.050 365.400 ;
        RECT 280.950 366.600 283.050 367.050 ;
        RECT 296.400 366.600 297.600 370.950 ;
        RECT 280.950 365.400 297.600 366.600 ;
        RECT 313.950 366.600 316.050 366.900 ;
        RECT 328.950 366.600 331.050 367.050 ;
        RECT 313.950 365.400 331.050 366.600 ;
        RECT 280.950 364.950 283.050 365.400 ;
        RECT 313.950 364.800 316.050 365.400 ;
        RECT 328.950 364.950 331.050 365.400 ;
        RECT 343.950 366.600 346.050 366.900 ;
        RECT 352.950 366.600 355.050 367.050 ;
        RECT 524.400 366.900 525.600 374.400 ;
        RECT 547.950 373.950 550.050 374.400 ;
        RECT 574.950 373.950 577.050 374.400 ;
        RECT 601.950 375.600 604.050 376.050 ;
        RECT 616.950 375.600 619.050 376.050 ;
        RECT 601.950 374.400 619.050 375.600 ;
        RECT 601.950 373.950 604.050 374.400 ;
        RECT 616.950 373.950 619.050 374.400 ;
        RECT 664.950 375.600 667.050 376.050 ;
        RECT 751.950 375.600 754.050 376.050 ;
        RECT 757.950 375.600 760.050 376.050 ;
        RECT 802.950 375.600 805.050 376.050 ;
        RECT 664.950 374.400 687.600 375.600 ;
        RECT 664.950 373.950 667.050 374.400 ;
        RECT 526.950 371.100 529.050 373.200 ;
        RECT 531.000 372.600 535.050 373.050 ;
        RECT 343.950 365.400 355.050 366.600 ;
        RECT 343.950 364.800 346.050 365.400 ;
        RECT 352.950 364.950 355.050 365.400 ;
        RECT 406.950 366.600 409.050 366.900 ;
        RECT 427.950 366.600 430.050 366.900 ;
        RECT 406.950 366.450 430.050 366.600 ;
        RECT 442.950 366.450 445.050 366.900 ;
        RECT 406.950 365.400 445.050 366.450 ;
        RECT 406.950 364.800 409.050 365.400 ;
        RECT 427.950 365.250 445.050 365.400 ;
        RECT 427.950 364.800 430.050 365.250 ;
        RECT 442.950 364.800 445.050 365.250 ;
        RECT 502.950 366.450 505.050 366.900 ;
        RECT 508.950 366.450 511.050 366.900 ;
        RECT 502.950 365.250 511.050 366.450 ;
        RECT 502.950 364.800 505.050 365.250 ;
        RECT 508.950 364.800 511.050 365.250 ;
        RECT 523.950 364.800 526.050 366.900 ;
        RECT 527.400 364.050 528.600 371.100 ;
        RECT 530.400 370.950 535.050 372.600 ;
        RECT 562.950 372.600 565.050 373.050 ;
        RECT 580.950 372.600 583.050 373.200 ;
        RECT 625.950 372.600 628.050 373.200 ;
        RECT 646.950 372.600 649.050 373.200 ;
        RECT 686.400 373.050 687.600 374.400 ;
        RECT 751.950 374.400 760.050 375.600 ;
        RECT 751.950 373.950 754.050 374.400 ;
        RECT 757.950 373.950 760.050 374.400 ;
        RECT 785.400 374.400 805.050 375.600 ;
        RECT 562.950 371.400 649.050 372.600 ;
        RECT 562.950 370.950 565.050 371.400 ;
        RECT 580.950 371.100 583.050 371.400 ;
        RECT 625.950 371.100 628.050 371.400 ;
        RECT 646.950 371.100 649.050 371.400 ;
        RECT 682.800 372.000 684.900 373.050 ;
        RECT 685.950 372.750 688.050 373.050 ;
        RECT 712.950 372.750 715.050 373.200 ;
        RECT 682.800 370.950 685.050 372.000 ;
        RECT 685.950 371.550 715.050 372.750 ;
        RECT 685.950 370.950 688.050 371.550 ;
        RECT 712.950 371.100 715.050 371.550 ;
        RECT 724.950 372.600 727.050 373.050 ;
        RECT 733.950 372.600 736.050 373.200 ;
        RECT 724.950 371.400 736.050 372.600 ;
        RECT 724.950 370.950 727.050 371.400 ;
        RECT 733.950 371.100 736.050 371.400 ;
        RECT 739.950 372.600 742.050 373.050 ;
        RECT 739.950 371.400 762.600 372.600 ;
        RECT 739.950 370.950 742.050 371.400 ;
        RECT 530.400 366.900 531.600 370.950 ;
        RECT 682.950 370.050 685.050 370.950 ;
        RECT 682.950 369.900 687.000 370.050 ;
        RECT 682.950 369.000 688.050 369.900 ;
        RECT 683.400 368.400 688.050 369.000 ;
        RECT 684.000 367.950 688.050 368.400 ;
        RECT 685.950 367.800 688.050 367.950 ;
        RECT 761.400 367.050 762.600 371.400 ;
        RECT 763.950 369.600 766.050 373.050 ;
        RECT 785.400 372.600 786.600 374.400 ;
        RECT 802.950 373.950 805.050 374.400 ;
        RECT 823.800 375.000 825.900 376.050 ;
        RECT 826.950 375.600 829.050 376.200 ;
        RECT 835.950 375.750 838.050 376.200 ;
        RECT 844.950 375.750 847.050 375.900 ;
        RECT 835.950 375.600 847.050 375.750 ;
        RECT 823.800 373.950 826.050 375.000 ;
        RECT 826.950 374.550 847.050 375.600 ;
        RECT 826.950 374.400 838.050 374.550 ;
        RECT 826.950 374.100 829.050 374.400 ;
        RECT 835.950 374.100 838.050 374.400 ;
        RECT 776.400 371.400 786.600 372.600 ;
        RECT 823.950 372.600 826.050 373.950 ;
        RECT 844.950 373.800 847.050 374.550 ;
        RECT 859.950 375.600 862.050 376.050 ;
        RECT 988.950 375.600 991.050 376.050 ;
        RECT 1000.950 375.600 1003.050 376.050 ;
        RECT 859.950 374.400 891.600 375.600 ;
        RECT 859.950 373.950 862.050 374.400 ;
        RECT 823.950 372.000 834.600 372.600 ;
        RECT 824.400 371.400 835.050 372.000 ;
        RECT 769.950 369.600 772.050 370.050 ;
        RECT 776.400 369.900 777.600 371.400 ;
        RECT 763.950 369.000 772.050 369.600 ;
        RECT 764.400 368.400 772.050 369.000 ;
        RECT 769.950 367.950 772.050 368.400 ;
        RECT 775.950 367.800 778.050 369.900 ;
        RECT 802.800 368.100 804.900 370.200 ;
        RECT 805.950 369.600 808.050 370.050 ;
        RECT 805.950 369.000 822.600 369.600 ;
        RECT 805.950 368.400 823.050 369.000 ;
        RECT 529.950 364.800 532.050 366.900 ;
        RECT 568.950 366.450 571.050 366.900 ;
        RECT 598.950 366.450 601.050 366.900 ;
        RECT 568.950 365.250 601.050 366.450 ;
        RECT 568.950 364.800 571.050 365.250 ;
        RECT 598.950 364.800 601.050 365.250 ;
        RECT 604.950 366.450 607.050 366.900 ;
        RECT 610.950 366.450 613.050 366.900 ;
        RECT 604.950 365.250 613.050 366.450 ;
        RECT 604.950 364.800 607.050 365.250 ;
        RECT 610.950 364.800 613.050 365.250 ;
        RECT 616.950 366.450 619.050 366.900 ;
        RECT 622.950 366.450 625.050 366.900 ;
        RECT 616.950 365.250 625.050 366.450 ;
        RECT 616.950 364.800 619.050 365.250 ;
        RECT 622.950 364.800 625.050 365.250 ;
        RECT 628.950 366.450 631.050 366.900 ;
        RECT 658.950 366.450 661.050 366.900 ;
        RECT 628.950 365.250 661.050 366.450 ;
        RECT 628.950 364.800 631.050 365.250 ;
        RECT 658.950 364.800 661.050 365.250 ;
        RECT 667.950 366.600 670.050 367.050 ;
        RECT 673.950 366.600 676.050 366.900 ;
        RECT 697.950 366.600 700.050 366.900 ;
        RECT 730.950 366.600 733.050 366.900 ;
        RECT 667.950 365.400 733.050 366.600 ;
        RECT 667.950 364.950 670.050 365.400 ;
        RECT 673.950 364.800 676.050 365.400 ;
        RECT 697.950 364.800 700.050 365.400 ;
        RECT 730.950 364.800 733.050 365.400 ;
        RECT 748.950 366.450 751.050 366.900 ;
        RECT 754.950 366.450 757.050 366.900 ;
        RECT 748.950 365.250 757.050 366.450 ;
        RECT 761.400 365.400 766.050 367.050 ;
        RECT 748.950 364.800 751.050 365.250 ;
        RECT 754.950 364.800 757.050 365.250 ;
        RECT 762.000 364.950 766.050 365.400 ;
        RECT 781.950 366.600 784.050 367.050 ;
        RECT 803.400 366.600 804.600 368.100 ;
        RECT 805.950 367.950 808.050 368.400 ;
        RECT 781.950 365.400 804.600 366.600 ;
        RECT 781.950 364.950 784.050 365.400 ;
        RECT 820.950 364.950 823.050 368.400 ;
        RECT 832.950 367.950 835.050 371.400 ;
        RECT 856.800 369.000 858.900 370.050 ;
        RECT 859.950 369.750 862.050 370.200 ;
        RECT 880.950 369.750 883.050 370.200 ;
        RECT 856.800 367.950 859.050 369.000 ;
        RECT 859.950 368.550 883.050 369.750 ;
        RECT 859.950 368.100 862.050 368.550 ;
        RECT 880.950 368.100 883.050 368.550 ;
        RECT 843.000 366.600 847.050 367.050 ;
        RECT 842.400 364.950 847.050 366.600 ;
        RECT 856.950 366.600 859.050 367.950 ;
        RECT 890.400 367.050 891.600 374.400 ;
        RECT 988.950 374.400 1003.050 375.600 ;
        RECT 988.950 373.950 991.050 374.400 ;
        RECT 1000.950 373.950 1003.050 374.400 ;
        RECT 1018.950 375.600 1021.050 376.050 ;
        RECT 1027.950 375.600 1030.050 376.050 ;
        RECT 1018.950 374.400 1030.050 375.600 ;
        RECT 1018.950 373.950 1021.050 374.400 ;
        RECT 1027.950 373.950 1030.050 374.400 ;
        RECT 901.950 372.600 904.050 373.050 ;
        RECT 916.950 372.750 919.050 373.200 ;
        RECT 922.950 372.750 925.050 373.200 ;
        RECT 916.950 372.600 925.050 372.750 ;
        RECT 901.950 371.550 925.050 372.600 ;
        RECT 901.950 371.400 919.050 371.550 ;
        RECT 901.950 370.950 904.050 371.400 ;
        RECT 916.950 371.100 919.050 371.400 ;
        RECT 922.950 371.100 925.050 371.550 ;
        RECT 928.950 372.600 931.050 373.050 ;
        RECT 937.950 372.600 940.050 373.200 ;
        RECT 949.950 372.600 952.050 373.050 ;
        RECT 928.950 371.400 940.050 372.600 ;
        RECT 928.950 370.950 931.050 371.400 ;
        RECT 937.950 371.100 940.050 371.400 ;
        RECT 941.400 371.400 952.050 372.600 ;
        RECT 941.400 369.600 942.600 371.400 ;
        RECT 949.950 370.950 952.050 371.400 ;
        RECT 976.950 372.600 979.050 373.050 ;
        RECT 985.950 372.750 988.050 373.200 ;
        RECT 991.950 372.750 994.050 373.200 ;
        RECT 976.950 371.400 984.600 372.600 ;
        RECT 976.950 370.950 979.050 371.400 ;
        RECT 926.400 368.400 942.600 369.600 ;
        RECT 983.400 369.600 984.600 371.400 ;
        RECT 985.950 371.550 994.050 372.750 ;
        RECT 985.950 371.100 988.050 371.550 ;
        RECT 991.950 371.100 994.050 371.550 ;
        RECT 1003.950 370.950 1006.050 373.050 ;
        RECT 983.400 368.400 993.600 369.600 ;
        RECT 856.950 366.000 888.600 366.600 ;
        RECT 857.400 365.400 888.600 366.000 ;
        RECT 115.950 363.600 118.050 364.050 ;
        RECT 130.950 363.600 133.050 364.050 ;
        RECT 115.950 362.400 133.050 363.600 ;
        RECT 115.950 361.950 118.050 362.400 ;
        RECT 130.950 361.950 133.050 362.400 ;
        RECT 142.950 363.600 145.050 364.050 ;
        RECT 151.950 363.600 154.050 364.050 ;
        RECT 142.950 362.400 154.050 363.600 ;
        RECT 142.950 361.950 145.050 362.400 ;
        RECT 151.950 361.950 154.050 362.400 ;
        RECT 232.950 363.600 235.050 364.050 ;
        RECT 250.950 363.600 253.050 364.050 ;
        RECT 265.950 363.600 268.050 364.050 ;
        RECT 232.950 362.400 268.050 363.600 ;
        RECT 232.950 361.950 235.050 362.400 ;
        RECT 250.950 361.950 253.050 362.400 ;
        RECT 265.950 361.950 268.050 362.400 ;
        RECT 274.950 363.600 277.050 364.050 ;
        RECT 289.950 363.600 292.050 364.050 ;
        RECT 274.950 362.400 292.050 363.600 ;
        RECT 274.950 361.950 277.050 362.400 ;
        RECT 289.950 361.950 292.050 362.400 ;
        RECT 526.950 361.950 529.050 364.050 ;
        RECT 574.950 363.600 577.050 364.050 ;
        RECT 592.950 363.600 595.050 364.050 ;
        RECT 574.950 362.400 595.050 363.600 ;
        RECT 574.950 361.950 577.050 362.400 ;
        RECT 592.950 361.950 595.050 362.400 ;
        RECT 640.950 363.600 643.050 364.050 ;
        RECT 661.950 363.600 664.050 364.050 ;
        RECT 640.950 362.400 664.050 363.600 ;
        RECT 640.950 361.950 643.050 362.400 ;
        RECT 661.950 361.950 664.050 362.400 ;
        RECT 679.950 363.600 682.050 364.050 ;
        RECT 685.950 363.600 688.050 364.050 ;
        RECT 679.950 362.400 688.050 363.600 ;
        RECT 679.950 361.950 682.050 362.400 ;
        RECT 685.950 361.950 688.050 362.400 ;
        RECT 826.950 363.600 829.050 364.050 ;
        RECT 842.400 363.600 843.600 364.950 ;
        RECT 826.950 362.400 843.600 363.600 ;
        RECT 887.400 363.600 888.600 365.400 ;
        RECT 889.950 364.950 892.050 367.050 ;
        RECT 919.950 366.600 922.050 366.900 ;
        RECT 926.400 366.600 927.600 368.400 ;
        RECT 919.950 365.400 927.600 366.600 ;
        RECT 940.950 366.600 943.050 366.900 ;
        RECT 964.950 366.600 967.050 366.900 ;
        RECT 940.950 365.400 967.050 366.600 ;
        RECT 919.950 364.800 922.050 365.400 ;
        RECT 940.950 364.800 943.050 365.400 ;
        RECT 964.950 364.800 967.050 365.400 ;
        RECT 970.950 366.600 973.050 366.900 ;
        RECT 979.950 366.600 982.050 367.050 ;
        RECT 970.950 365.400 982.050 366.600 ;
        RECT 992.400 366.600 993.600 368.400 ;
        RECT 1004.400 367.050 1005.600 370.950 ;
        RECT 994.950 366.600 997.050 366.900 ;
        RECT 992.400 365.400 997.050 366.600 ;
        RECT 970.950 364.800 973.050 365.400 ;
        RECT 979.950 364.950 982.050 365.400 ;
        RECT 994.950 364.800 997.050 365.400 ;
        RECT 1003.950 364.950 1006.050 367.050 ;
        RECT 1009.950 366.600 1012.050 367.050 ;
        RECT 1021.950 366.600 1024.050 366.900 ;
        RECT 1009.950 365.400 1024.050 366.600 ;
        RECT 1009.950 364.950 1012.050 365.400 ;
        RECT 1021.950 364.800 1024.050 365.400 ;
        RECT 1027.950 366.450 1030.050 366.900 ;
        RECT 1033.950 366.450 1036.050 366.900 ;
        RECT 1027.950 365.250 1036.050 366.450 ;
        RECT 1027.950 364.800 1030.050 365.250 ;
        RECT 1033.950 364.800 1036.050 365.250 ;
        RECT 943.950 363.600 946.050 364.050 ;
        RECT 958.950 363.600 961.050 364.050 ;
        RECT 887.400 362.400 918.600 363.600 ;
        RECT 826.950 361.950 829.050 362.400 ;
        RECT 19.950 360.600 22.050 361.050 ;
        RECT 25.950 360.600 28.050 361.050 ;
        RECT 64.950 360.600 67.050 361.050 ;
        RECT 79.950 360.600 82.050 361.050 ;
        RECT 19.950 359.400 82.050 360.600 ;
        RECT 19.950 358.950 22.050 359.400 ;
        RECT 25.950 358.950 28.050 359.400 ;
        RECT 64.950 358.950 67.050 359.400 ;
        RECT 79.950 358.950 82.050 359.400 ;
        RECT 139.950 360.600 142.050 361.050 ;
        RECT 166.950 360.600 169.050 361.050 ;
        RECT 139.950 359.400 169.050 360.600 ;
        RECT 139.950 358.950 142.050 359.400 ;
        RECT 166.950 358.950 169.050 359.400 ;
        RECT 172.950 360.600 175.050 361.050 ;
        RECT 178.950 360.600 181.050 361.050 ;
        RECT 172.950 359.400 181.050 360.600 ;
        RECT 172.950 358.950 175.050 359.400 ;
        RECT 178.950 358.950 181.050 359.400 ;
        RECT 313.950 360.600 316.050 361.050 ;
        RECT 322.950 360.600 325.050 361.050 ;
        RECT 313.950 359.400 325.050 360.600 ;
        RECT 313.950 358.950 316.050 359.400 ;
        RECT 322.950 358.950 325.050 359.400 ;
        RECT 550.950 360.600 553.050 361.050 ;
        RECT 562.950 360.600 565.050 361.050 ;
        RECT 550.950 359.400 565.050 360.600 ;
        RECT 550.950 358.950 553.050 359.400 ;
        RECT 562.950 358.950 565.050 359.400 ;
        RECT 598.950 360.600 601.050 361.050 ;
        RECT 607.950 360.600 610.050 361.050 ;
        RECT 598.950 359.400 610.050 360.600 ;
        RECT 598.950 358.950 601.050 359.400 ;
        RECT 607.950 358.950 610.050 359.400 ;
        RECT 652.950 360.600 655.050 361.050 ;
        RECT 658.950 360.600 661.050 361.050 ;
        RECT 703.950 360.600 706.050 361.050 ;
        RECT 652.950 359.400 706.050 360.600 ;
        RECT 652.950 358.950 655.050 359.400 ;
        RECT 658.950 358.950 661.050 359.400 ;
        RECT 703.950 358.950 706.050 359.400 ;
        RECT 724.950 360.600 727.050 361.050 ;
        RECT 760.950 360.600 763.050 361.050 ;
        RECT 724.950 359.400 763.050 360.600 ;
        RECT 724.950 358.950 727.050 359.400 ;
        RECT 760.950 358.950 763.050 359.400 ;
        RECT 775.950 360.600 778.050 361.050 ;
        RECT 781.950 360.600 784.050 361.050 ;
        RECT 775.950 359.400 784.050 360.600 ;
        RECT 775.950 358.950 778.050 359.400 ;
        RECT 781.950 358.950 784.050 359.400 ;
        RECT 844.950 360.600 847.050 361.050 ;
        RECT 886.950 360.600 889.050 361.050 ;
        RECT 900.000 360.900 903.000 361.050 ;
        RECT 844.950 359.400 889.050 360.600 ;
        RECT 844.950 358.950 847.050 359.400 ;
        RECT 886.950 358.950 889.050 359.400 ;
        RECT 898.950 360.600 903.000 360.900 ;
        RECT 917.400 360.600 918.600 362.400 ;
        RECT 943.950 362.400 961.050 363.600 ;
        RECT 943.950 361.950 946.050 362.400 ;
        RECT 958.950 361.950 961.050 362.400 ;
        RECT 967.950 363.600 970.050 364.050 ;
        RECT 982.950 363.600 985.050 364.050 ;
        RECT 967.950 362.400 985.050 363.600 ;
        RECT 967.950 361.950 970.050 362.400 ;
        RECT 982.950 361.950 985.050 362.400 ;
        RECT 949.950 360.600 952.050 361.050 ;
        RECT 898.950 358.950 903.600 360.600 ;
        RECT 917.400 359.400 952.050 360.600 ;
        RECT 949.950 358.950 952.050 359.400 ;
        RECT 1000.950 360.600 1003.050 361.050 ;
        RECT 1015.950 360.600 1018.050 361.050 ;
        RECT 1000.950 359.400 1018.050 360.600 ;
        RECT 1000.950 358.950 1003.050 359.400 ;
        RECT 1015.950 358.950 1018.050 359.400 ;
        RECT 898.950 358.800 901.050 358.950 ;
        RECT 223.950 357.600 226.050 358.050 ;
        RECT 232.950 357.600 235.050 358.050 ;
        RECT 223.950 356.400 235.050 357.600 ;
        RECT 223.950 355.950 226.050 356.400 ;
        RECT 232.950 355.950 235.050 356.400 ;
        RECT 445.950 357.600 448.050 358.050 ;
        RECT 475.950 357.600 478.050 358.050 ;
        RECT 445.950 356.400 478.050 357.600 ;
        RECT 445.950 355.950 448.050 356.400 ;
        RECT 475.950 355.950 478.050 356.400 ;
        RECT 727.950 357.600 730.050 358.050 ;
        RECT 736.950 357.600 739.050 358.050 ;
        RECT 895.950 357.600 898.050 358.050 ;
        RECT 727.950 356.400 739.050 357.600 ;
        RECT 854.400 357.000 898.050 357.600 ;
        RECT 727.950 355.950 730.050 356.400 ;
        RECT 736.950 355.950 739.050 356.400 ;
        RECT 853.950 356.400 898.050 357.000 ;
        RECT 902.400 357.600 903.600 358.950 ;
        RECT 919.950 357.600 922.050 358.050 ;
        RECT 902.400 356.400 922.050 357.600 ;
        RECT 115.950 354.600 118.050 355.050 ;
        RECT 247.950 354.600 250.050 355.050 ;
        RECT 115.950 353.400 250.050 354.600 ;
        RECT 115.950 352.950 118.050 353.400 ;
        RECT 247.950 352.950 250.050 353.400 ;
        RECT 373.950 354.600 376.050 355.050 ;
        RECT 514.950 354.600 517.050 355.050 ;
        RECT 373.950 353.400 517.050 354.600 ;
        RECT 373.950 352.950 376.050 353.400 ;
        RECT 514.950 352.950 517.050 353.400 ;
        RECT 520.950 354.600 523.050 355.050 ;
        RECT 565.950 354.600 568.050 355.050 ;
        RECT 520.950 353.400 568.050 354.600 ;
        RECT 520.950 352.950 523.050 353.400 ;
        RECT 565.950 352.950 568.050 353.400 ;
        RECT 631.950 354.600 634.050 355.050 ;
        RECT 649.950 354.600 652.050 355.050 ;
        RECT 631.950 353.400 652.050 354.600 ;
        RECT 631.950 352.950 634.050 353.400 ;
        RECT 649.950 352.950 652.050 353.400 ;
        RECT 697.950 354.600 700.050 355.050 ;
        RECT 739.950 354.600 742.050 355.050 ;
        RECT 697.950 353.400 742.050 354.600 ;
        RECT 697.950 352.950 700.050 353.400 ;
        RECT 739.950 352.950 742.050 353.400 ;
        RECT 745.950 354.600 748.050 355.050 ;
        RECT 751.950 354.600 754.050 355.050 ;
        RECT 775.950 354.600 778.050 355.050 ;
        RECT 745.950 353.400 754.050 354.600 ;
        RECT 745.950 352.950 748.050 353.400 ;
        RECT 751.950 352.950 754.050 353.400 ;
        RECT 755.400 353.400 778.050 354.600 ;
        RECT 7.950 351.600 10.050 352.050 ;
        RECT 28.950 351.600 31.050 352.050 ;
        RECT 7.950 350.400 31.050 351.600 ;
        RECT 7.950 349.950 10.050 350.400 ;
        RECT 28.950 349.950 31.050 350.400 ;
        RECT 37.950 349.950 40.050 352.050 ;
        RECT 70.950 351.600 73.050 352.050 ;
        RECT 127.950 351.600 130.050 352.050 ;
        RECT 70.950 350.400 130.050 351.600 ;
        RECT 70.950 349.950 73.050 350.400 ;
        RECT 127.950 349.950 130.050 350.400 ;
        RECT 286.950 351.600 289.050 352.050 ;
        RECT 298.950 351.600 301.050 352.050 ;
        RECT 286.950 350.400 301.050 351.600 ;
        RECT 286.950 349.950 289.050 350.400 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 358.950 351.600 361.050 352.050 ;
        RECT 376.800 351.600 378.900 352.050 ;
        RECT 358.950 350.400 378.900 351.600 ;
        RECT 358.950 349.950 361.050 350.400 ;
        RECT 376.800 349.950 378.900 350.400 ;
        RECT 379.950 351.600 382.050 352.050 ;
        RECT 391.950 351.600 394.050 352.050 ;
        RECT 379.950 350.400 394.050 351.600 ;
        RECT 379.950 349.950 382.050 350.400 ;
        RECT 391.950 349.950 394.050 350.400 ;
        RECT 412.950 351.600 415.050 352.050 ;
        RECT 445.950 351.600 448.050 352.050 ;
        RECT 676.950 351.600 679.050 352.050 ;
        RECT 412.950 350.400 448.050 351.600 ;
        RECT 412.950 349.950 415.050 350.400 ;
        RECT 445.950 349.950 448.050 350.400 ;
        RECT 587.400 350.400 679.050 351.600 ;
        RECT 38.400 345.600 39.600 349.950 ;
        RECT 587.400 349.050 588.600 350.400 ;
        RECT 676.950 349.950 679.050 350.400 ;
        RECT 733.950 351.600 736.050 352.050 ;
        RECT 755.400 351.600 756.600 353.400 ;
        RECT 775.950 352.950 778.050 353.400 ;
        RECT 781.950 354.600 784.050 355.050 ;
        RECT 781.950 353.400 822.600 354.600 ;
        RECT 781.950 352.950 784.050 353.400 ;
        RECT 733.950 350.400 756.600 351.600 ;
        RECT 821.400 351.600 822.600 353.400 ;
        RECT 853.950 352.950 856.050 356.400 ;
        RECT 895.950 355.950 898.050 356.400 ;
        RECT 919.950 355.950 922.050 356.400 ;
        RECT 967.950 357.600 970.050 358.050 ;
        RECT 1003.950 357.600 1006.050 358.050 ;
        RECT 967.950 356.400 1006.050 357.600 ;
        RECT 967.950 355.950 970.050 356.400 ;
        RECT 1003.950 355.950 1006.050 356.400 ;
        RECT 988.950 354.600 991.050 355.050 ;
        RECT 1012.950 354.600 1015.050 355.050 ;
        RECT 1018.950 354.600 1021.050 355.050 ;
        RECT 988.950 353.400 1021.050 354.600 ;
        RECT 988.950 352.950 991.050 353.400 ;
        RECT 1012.950 352.950 1015.050 353.400 ;
        RECT 1018.950 352.950 1021.050 353.400 ;
        RECT 844.950 351.600 847.050 352.050 ;
        RECT 821.400 350.400 847.050 351.600 ;
        RECT 733.950 349.950 736.050 350.400 ;
        RECT 844.950 349.950 847.050 350.400 ;
        RECT 856.950 351.600 859.050 352.050 ;
        RECT 898.950 351.600 901.050 352.050 ;
        RECT 856.950 350.400 901.050 351.600 ;
        RECT 856.950 349.950 859.050 350.400 ;
        RECT 898.950 349.950 901.050 350.400 ;
        RECT 940.950 351.600 943.050 352.050 ;
        RECT 952.950 351.600 955.050 352.050 ;
        RECT 940.950 350.400 955.050 351.600 ;
        RECT 940.950 349.950 943.050 350.400 ;
        RECT 952.950 349.950 955.050 350.400 ;
        RECT 991.950 351.600 994.050 352.050 ;
        RECT 1006.950 351.600 1009.050 352.050 ;
        RECT 991.950 350.400 1009.050 351.600 ;
        RECT 991.950 349.950 994.050 350.400 ;
        RECT 1006.950 349.950 1009.050 350.400 ;
        RECT 136.950 348.600 139.050 349.050 ;
        RECT 220.950 348.600 223.050 349.050 ;
        RECT 136.950 347.400 223.050 348.600 ;
        RECT 136.950 346.950 139.050 347.400 ;
        RECT 220.950 346.950 223.050 347.400 ;
        RECT 262.950 348.600 265.050 349.050 ;
        RECT 301.950 348.600 304.050 349.050 ;
        RECT 310.950 348.600 313.050 349.050 ;
        RECT 262.950 347.400 313.050 348.600 ;
        RECT 262.950 346.950 265.050 347.400 ;
        RECT 301.950 346.950 304.050 347.400 ;
        RECT 310.950 346.950 313.050 347.400 ;
        RECT 466.950 348.600 469.050 349.050 ;
        RECT 544.950 348.600 547.050 349.050 ;
        RECT 466.950 347.400 547.050 348.600 ;
        RECT 466.950 346.950 469.050 347.400 ;
        RECT 544.950 346.950 547.050 347.400 ;
        RECT 562.950 348.600 565.050 349.050 ;
        RECT 577.950 348.600 580.050 349.050 ;
        RECT 562.950 347.400 580.050 348.600 ;
        RECT 562.950 346.950 565.050 347.400 ;
        RECT 577.950 346.950 580.050 347.400 ;
        RECT 583.950 347.400 588.600 349.050 ;
        RECT 616.950 348.600 619.050 349.050 ;
        RECT 634.950 348.600 637.050 349.050 ;
        RECT 616.950 347.400 637.050 348.600 ;
        RECT 583.950 346.950 588.000 347.400 ;
        RECT 616.950 346.950 619.050 347.400 ;
        RECT 634.950 346.950 637.050 347.400 ;
        RECT 679.950 348.600 682.050 349.050 ;
        RECT 706.950 348.600 709.050 349.050 ;
        RECT 679.950 347.400 709.050 348.600 ;
        RECT 679.950 346.950 682.050 347.400 ;
        RECT 706.950 346.950 709.050 347.400 ;
        RECT 715.950 348.600 718.050 349.050 ;
        RECT 724.950 348.600 727.050 349.050 ;
        RECT 715.950 347.400 727.050 348.600 ;
        RECT 715.950 346.950 718.050 347.400 ;
        RECT 724.950 346.950 727.050 347.400 ;
        RECT 730.950 348.600 733.050 349.050 ;
        RECT 766.950 348.600 769.050 349.050 ;
        RECT 730.950 347.400 769.050 348.600 ;
        RECT 730.950 346.950 733.050 347.400 ;
        RECT 766.950 346.950 769.050 347.400 ;
        RECT 817.950 348.600 820.050 349.050 ;
        RECT 823.950 348.600 826.050 349.050 ;
        RECT 880.950 348.600 883.050 349.050 ;
        RECT 955.950 348.600 958.050 349.050 ;
        RECT 961.950 348.600 964.050 349.050 ;
        RECT 817.950 347.400 826.050 348.600 ;
        RECT 817.950 346.950 820.050 347.400 ;
        RECT 823.950 346.950 826.050 347.400 ;
        RECT 860.400 347.400 894.600 348.600 ;
        RECT 35.400 344.400 39.600 345.600 ;
        RECT 181.950 345.600 184.050 346.050 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 181.950 344.400 202.050 345.600 ;
        RECT 35.400 339.600 36.600 344.400 ;
        RECT 181.950 343.950 184.050 344.400 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 229.950 345.600 232.050 346.050 ;
        RECT 259.950 345.600 262.050 346.050 ;
        RECT 229.950 344.400 262.050 345.600 ;
        RECT 229.950 343.950 232.050 344.400 ;
        RECT 259.950 343.950 262.050 344.400 ;
        RECT 280.950 345.600 283.050 346.050 ;
        RECT 292.950 345.600 295.050 346.050 ;
        RECT 280.950 344.400 295.050 345.600 ;
        RECT 280.950 343.950 283.050 344.400 ;
        RECT 292.950 343.950 295.050 344.400 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 385.950 345.600 388.050 346.050 ;
        RECT 355.950 344.400 388.050 345.600 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 385.950 343.950 388.050 344.400 ;
        RECT 439.950 345.600 442.050 346.050 ;
        RECT 460.950 345.600 463.050 346.050 ;
        RECT 439.950 344.400 463.050 345.600 ;
        RECT 439.950 343.950 442.050 344.400 ;
        RECT 460.950 343.950 463.050 344.400 ;
        RECT 553.950 345.600 556.050 346.050 ;
        RECT 559.950 345.600 562.050 346.050 ;
        RECT 553.950 344.400 562.050 345.600 ;
        RECT 553.950 343.950 556.050 344.400 ;
        RECT 559.950 343.950 562.050 344.400 ;
        RECT 589.950 345.600 592.050 346.050 ;
        RECT 601.950 345.600 604.050 346.050 ;
        RECT 589.950 344.400 604.050 345.600 ;
        RECT 589.950 343.950 592.050 344.400 ;
        RECT 601.950 343.950 604.050 344.400 ;
        RECT 637.950 345.600 640.050 346.050 ;
        RECT 673.950 345.600 676.050 346.050 ;
        RECT 637.950 344.400 676.050 345.600 ;
        RECT 637.950 343.950 640.050 344.400 ;
        RECT 673.950 343.950 676.050 344.400 ;
        RECT 769.950 345.600 772.050 346.050 ;
        RECT 799.950 345.600 802.050 346.050 ;
        RECT 769.950 344.400 802.050 345.600 ;
        RECT 769.950 343.950 772.050 344.400 ;
        RECT 799.950 343.950 802.050 344.400 ;
        RECT 844.950 345.600 847.050 346.050 ;
        RECT 860.400 345.600 861.600 347.400 ;
        RECT 880.950 346.950 883.050 347.400 ;
        RECT 844.950 344.400 861.600 345.600 ;
        RECT 893.400 345.600 894.600 347.400 ;
        RECT 955.950 347.400 964.050 348.600 ;
        RECT 955.950 346.950 958.050 347.400 ;
        RECT 961.950 346.950 964.050 347.400 ;
        RECT 904.950 345.600 907.050 346.050 ;
        RECT 893.400 344.400 907.050 345.600 ;
        RECT 844.950 343.950 847.050 344.400 ;
        RECT 904.950 343.950 907.050 344.400 ;
        RECT 916.950 345.600 919.050 346.050 ;
        RECT 925.950 345.600 928.050 346.050 ;
        RECT 916.950 344.400 928.050 345.600 ;
        RECT 916.950 343.950 919.050 344.400 ;
        RECT 925.950 343.950 928.050 344.400 ;
        RECT 946.950 345.600 949.050 346.050 ;
        RECT 979.950 345.600 982.050 346.050 ;
        RECT 1012.950 345.600 1015.050 346.050 ;
        RECT 1036.950 345.600 1039.050 346.050 ;
        RECT 946.950 344.400 1002.600 345.600 ;
        RECT 946.950 343.950 949.050 344.400 ;
        RECT 979.950 343.950 982.050 344.400 ;
        RECT 55.950 342.600 58.050 343.050 ;
        RECT 109.950 342.600 112.050 343.050 ;
        RECT 55.950 341.400 112.050 342.600 ;
        RECT 55.950 340.950 58.050 341.400 ;
        RECT 109.950 340.950 112.050 341.400 ;
        RECT 32.400 338.400 36.600 339.600 ;
        RECT 139.950 339.750 142.050 340.200 ;
        RECT 148.950 339.750 151.050 340.200 ;
        RECT 139.950 338.550 151.050 339.750 ;
        RECT 7.950 334.950 10.050 337.050 ;
        RECT 4.950 330.600 7.050 330.900 ;
        RECT 8.400 330.600 9.600 334.950 ;
        RECT 32.400 334.050 33.600 338.400 ;
        RECT 139.950 338.100 142.050 338.550 ;
        RECT 148.950 338.100 151.050 338.550 ;
        RECT 163.950 339.600 166.050 340.050 ;
        RECT 172.950 339.600 175.050 340.200 ;
        RECT 163.950 338.400 175.050 339.600 ;
        RECT 163.950 337.950 166.050 338.400 ;
        RECT 172.950 338.100 175.050 338.400 ;
        RECT 187.950 339.750 190.050 340.200 ;
        RECT 193.950 339.750 196.050 340.200 ;
        RECT 187.950 338.550 196.050 339.750 ;
        RECT 226.950 339.600 229.050 343.050 ;
        RECT 274.950 342.600 277.050 343.050 ;
        RECT 304.950 342.600 307.050 343.050 ;
        RECT 274.950 341.400 309.600 342.600 ;
        RECT 274.950 340.950 277.050 341.400 ;
        RECT 304.950 340.950 307.050 341.400 ;
        RECT 232.950 339.600 235.050 340.050 ;
        RECT 226.950 339.000 235.050 339.600 ;
        RECT 187.950 338.100 190.050 338.550 ;
        RECT 193.950 338.100 196.050 338.550 ;
        RECT 227.400 338.400 235.050 339.000 ;
        RECT 232.950 337.950 235.050 338.400 ;
        RECT 241.950 338.100 244.050 340.200 ;
        RECT 268.950 339.750 271.050 340.200 ;
        RECT 277.950 339.750 280.050 340.050 ;
        RECT 283.950 339.750 286.050 340.200 ;
        RECT 308.400 340.050 309.600 341.400 ;
        RECT 349.950 340.950 352.050 343.050 ;
        RECT 484.950 342.600 487.050 343.050 ;
        RECT 514.950 342.600 517.050 343.050 ;
        RECT 484.950 341.400 517.050 342.600 ;
        RECT 484.950 340.950 487.050 341.400 ;
        RECT 514.950 340.950 517.050 341.400 ;
        RECT 526.950 342.600 529.050 343.050 ;
        RECT 538.950 342.600 541.050 343.050 ;
        RECT 583.950 342.600 586.050 343.050 ;
        RECT 526.950 341.400 586.050 342.600 ;
        RECT 526.950 340.950 529.050 341.400 ;
        RECT 538.950 340.950 541.050 341.400 ;
        RECT 583.950 340.950 586.050 341.400 ;
        RECT 676.950 342.600 679.050 343.050 ;
        RECT 718.950 342.600 721.050 343.050 ;
        RECT 676.950 341.400 721.050 342.600 ;
        RECT 676.950 340.950 679.050 341.400 ;
        RECT 718.950 340.950 721.050 341.400 ;
        RECT 727.950 342.600 730.050 343.050 ;
        RECT 736.950 342.600 739.050 343.050 ;
        RECT 748.950 342.600 751.050 343.050 ;
        RECT 727.950 341.400 739.050 342.600 ;
        RECT 727.950 340.950 730.050 341.400 ;
        RECT 736.950 340.950 739.050 341.400 ;
        RECT 740.400 341.400 751.050 342.600 ;
        RECT 268.950 338.550 286.050 339.750 ;
        RECT 268.950 338.100 271.050 338.550 ;
        RECT 242.400 334.050 243.600 338.100 ;
        RECT 277.950 337.950 280.050 338.550 ;
        RECT 283.950 338.100 286.050 338.550 ;
        RECT 307.950 339.600 310.050 340.050 ;
        RECT 322.950 339.600 325.050 340.200 ;
        RECT 307.950 338.400 325.050 339.600 ;
        RECT 307.950 337.950 310.050 338.400 ;
        RECT 322.950 338.100 325.050 338.400 ;
        RECT 334.950 339.600 337.050 340.050 ;
        RECT 346.950 339.600 349.050 340.200 ;
        RECT 334.950 338.400 349.050 339.600 ;
        RECT 334.950 337.950 337.050 338.400 ;
        RECT 346.950 338.100 349.050 338.400 ;
        RECT 350.400 336.600 351.600 340.950 ;
        RECT 358.950 339.750 361.050 340.200 ;
        RECT 364.950 339.750 367.050 340.200 ;
        RECT 358.950 338.550 367.050 339.750 ;
        RECT 358.950 338.100 361.050 338.550 ;
        RECT 364.950 338.100 367.050 338.550 ;
        RECT 433.950 339.750 436.050 340.200 ;
        RECT 454.950 339.750 457.050 340.200 ;
        RECT 433.950 338.550 457.050 339.750 ;
        RECT 433.950 338.100 436.050 338.550 ;
        RECT 454.950 338.100 457.050 338.550 ;
        RECT 478.950 339.750 481.050 340.200 ;
        RECT 484.950 339.750 487.050 340.200 ;
        RECT 478.950 338.550 487.050 339.750 ;
        RECT 478.950 338.100 481.050 338.550 ;
        RECT 484.950 338.100 487.050 338.550 ;
        RECT 490.950 339.600 493.050 340.200 ;
        RECT 505.950 339.600 508.050 340.050 ;
        RECT 490.950 338.400 508.050 339.600 ;
        RECT 490.950 338.100 493.050 338.400 ;
        RECT 505.950 337.950 508.050 338.400 ;
        RECT 568.950 339.600 571.050 340.200 ;
        RECT 580.950 339.600 583.050 340.050 ;
        RECT 568.950 338.400 583.050 339.600 ;
        RECT 568.950 338.100 571.050 338.400 ;
        RECT 580.950 337.950 583.050 338.400 ;
        RECT 595.950 339.750 598.050 340.200 ;
        RECT 604.950 339.750 607.050 340.200 ;
        RECT 595.950 339.600 607.050 339.750 ;
        RECT 622.950 339.600 625.050 340.200 ;
        RECT 595.950 338.550 625.050 339.600 ;
        RECT 595.950 338.100 598.050 338.550 ;
        RECT 604.950 338.400 625.050 338.550 ;
        RECT 604.950 338.100 607.050 338.400 ;
        RECT 622.950 338.100 625.050 338.400 ;
        RECT 667.950 339.750 670.050 340.200 ;
        RECT 673.950 339.750 676.050 340.200 ;
        RECT 667.950 338.550 676.050 339.750 ;
        RECT 667.950 338.100 670.050 338.550 ;
        RECT 673.950 338.100 676.050 338.550 ;
        RECT 679.950 339.600 682.050 340.200 ;
        RECT 740.400 339.600 741.600 341.400 ;
        RECT 748.950 340.950 751.050 341.400 ;
        RECT 811.950 342.600 814.050 343.050 ;
        RECT 820.950 342.600 823.050 343.050 ;
        RECT 811.950 341.400 823.050 342.600 ;
        RECT 811.950 340.950 814.050 341.400 ;
        RECT 820.950 340.950 823.050 341.400 ;
        RECT 889.950 342.600 892.050 343.050 ;
        RECT 907.950 342.600 910.050 343.050 ;
        RECT 889.950 341.400 910.050 342.600 ;
        RECT 889.950 340.950 892.050 341.400 ;
        RECT 907.950 340.950 910.050 341.400 ;
        RECT 928.950 342.600 931.050 343.050 ;
        RECT 937.950 342.600 940.050 343.050 ;
        RECT 928.950 341.400 940.050 342.600 ;
        RECT 928.950 340.950 931.050 341.400 ;
        RECT 937.950 340.950 940.050 341.400 ;
        RECT 949.950 342.600 952.050 343.050 ;
        RECT 964.950 342.600 967.050 343.050 ;
        RECT 949.950 341.400 967.050 342.600 ;
        RECT 949.950 340.950 952.050 341.400 ;
        RECT 964.950 340.950 967.050 341.400 ;
        RECT 679.950 338.400 687.600 339.600 ;
        RECT 679.950 338.100 682.050 338.400 ;
        RECT 28.950 332.400 33.600 334.050 ;
        RECT 130.950 333.600 133.050 333.900 ;
        RECT 139.950 333.600 142.050 334.050 ;
        RECT 130.950 332.400 142.050 333.600 ;
        RECT 28.950 331.950 33.000 332.400 ;
        RECT 130.950 331.800 133.050 332.400 ;
        RECT 139.950 331.950 142.050 332.400 ;
        RECT 151.950 333.600 154.050 333.900 ;
        RECT 160.950 333.600 163.050 334.050 ;
        RECT 151.950 332.400 163.050 333.600 ;
        RECT 151.950 331.800 154.050 332.400 ;
        RECT 160.950 331.950 163.050 332.400 ;
        RECT 166.950 333.600 169.050 334.050 ;
        RECT 175.950 333.600 178.050 333.900 ;
        RECT 214.950 333.600 217.050 334.050 ;
        RECT 166.950 332.400 217.050 333.600 ;
        RECT 166.950 331.950 169.050 332.400 ;
        RECT 175.950 331.800 178.050 332.400 ;
        RECT 214.950 331.950 217.050 332.400 ;
        RECT 238.950 332.400 243.600 334.050 ;
        RECT 245.400 335.400 351.600 336.600 ;
        RECT 245.400 333.900 246.600 335.400 ;
        RECT 350.400 333.900 351.600 335.400 ;
        RECT 238.950 331.950 243.000 332.400 ;
        RECT 244.950 331.800 247.050 333.900 ;
        RECT 250.950 333.450 253.050 333.900 ;
        RECT 283.950 333.450 286.050 333.900 ;
        RECT 250.950 332.250 286.050 333.450 ;
        RECT 250.950 331.800 253.050 332.250 ;
        RECT 283.950 331.800 286.050 332.250 ;
        RECT 295.950 333.450 298.050 333.900 ;
        RECT 307.800 333.450 309.900 333.900 ;
        RECT 295.950 332.250 309.900 333.450 ;
        RECT 295.950 331.800 298.050 332.250 ;
        RECT 307.800 331.800 309.900 332.250 ;
        RECT 310.950 333.450 313.050 333.900 ;
        RECT 319.950 333.450 322.050 333.900 ;
        RECT 310.950 332.250 322.050 333.450 ;
        RECT 310.950 331.800 313.050 332.250 ;
        RECT 319.950 331.800 322.050 332.250 ;
        RECT 325.950 333.450 328.050 333.900 ;
        RECT 334.950 333.450 337.050 333.900 ;
        RECT 325.950 332.250 337.050 333.450 ;
        RECT 325.950 331.800 328.050 332.250 ;
        RECT 334.950 331.800 337.050 332.250 ;
        RECT 349.950 331.800 352.050 333.900 ;
        RECT 367.950 333.600 370.050 333.900 ;
        RECT 376.950 333.600 379.050 337.050 ;
        RECT 601.950 336.600 604.050 337.050 ;
        RECT 658.950 336.600 661.050 337.050 ;
        RECT 601.950 335.400 661.050 336.600 ;
        RECT 601.950 334.950 604.050 335.400 ;
        RECT 658.950 334.950 661.050 335.400 ;
        RECT 367.950 333.000 379.050 333.600 ;
        RECT 409.950 333.600 412.050 334.050 ;
        RECT 439.950 333.600 442.050 334.050 ;
        RECT 367.950 332.400 378.600 333.000 ;
        RECT 409.950 332.400 442.050 333.600 ;
        RECT 367.950 331.800 370.050 332.400 ;
        RECT 409.950 331.950 412.050 332.400 ;
        RECT 439.950 331.950 442.050 332.400 ;
        RECT 445.950 333.450 448.050 333.900 ;
        RECT 457.950 333.450 460.050 333.900 ;
        RECT 445.950 332.250 460.050 333.450 ;
        RECT 445.950 331.800 448.050 332.250 ;
        RECT 457.950 331.800 460.050 332.250 ;
        RECT 475.950 333.450 478.050 333.900 ;
        RECT 493.950 333.450 496.050 333.900 ;
        RECT 475.950 332.250 496.050 333.450 ;
        RECT 475.950 331.800 478.050 332.250 ;
        RECT 493.950 331.800 496.050 332.250 ;
        RECT 505.950 333.450 508.050 333.900 ;
        RECT 517.950 333.450 520.050 333.900 ;
        RECT 505.950 332.250 520.050 333.450 ;
        RECT 505.950 331.800 508.050 332.250 ;
        RECT 517.950 331.800 520.050 332.250 ;
        RECT 580.950 333.450 583.050 333.900 ;
        RECT 586.950 333.450 589.050 333.900 ;
        RECT 580.950 332.250 589.050 333.450 ;
        RECT 580.950 331.800 583.050 332.250 ;
        RECT 586.950 331.800 589.050 332.250 ;
        RECT 607.950 333.450 610.050 333.900 ;
        RECT 619.950 333.450 622.050 333.900 ;
        RECT 607.950 332.250 622.050 333.450 ;
        RECT 607.950 331.800 610.050 332.250 ;
        RECT 619.950 331.800 622.050 332.250 ;
        RECT 634.950 333.450 637.050 333.900 ;
        RECT 640.950 333.450 643.050 333.900 ;
        RECT 634.950 332.250 643.050 333.450 ;
        RECT 659.400 333.600 660.600 334.950 ;
        RECT 686.400 334.050 687.600 338.400 ;
        RECT 737.400 338.400 741.600 339.600 ;
        RECT 754.950 339.600 757.050 340.050 ;
        RECT 763.950 339.600 766.050 340.200 ;
        RECT 754.950 338.400 766.050 339.600 ;
        RECT 670.950 333.600 673.050 334.050 ;
        RECT 676.950 333.600 679.050 333.900 ;
        RECT 659.400 332.400 679.050 333.600 ;
        RECT 634.950 331.800 637.050 332.250 ;
        RECT 640.950 331.800 643.050 332.250 ;
        RECT 670.950 331.950 673.050 332.400 ;
        RECT 676.950 331.800 679.050 332.400 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 737.400 333.900 738.600 338.400 ;
        RECT 754.950 337.950 757.050 338.400 ;
        RECT 763.950 338.100 766.050 338.400 ;
        RECT 778.950 339.750 781.050 340.200 ;
        RECT 787.950 339.750 790.050 340.200 ;
        RECT 778.950 338.550 790.050 339.750 ;
        RECT 778.950 338.100 781.050 338.550 ;
        RECT 787.950 338.100 790.050 338.550 ;
        RECT 793.950 339.600 796.050 340.200 ;
        RECT 805.950 339.600 808.050 340.050 ;
        RECT 793.950 338.400 808.050 339.600 ;
        RECT 793.950 338.100 796.050 338.400 ;
        RECT 805.950 337.950 808.050 338.400 ;
        RECT 847.950 339.600 850.050 340.200 ;
        RECT 859.950 339.600 862.050 340.050 ;
        RECT 847.950 338.400 862.050 339.600 ;
        RECT 847.950 338.100 850.050 338.400 ;
        RECT 859.950 337.950 862.050 338.400 ;
        RECT 865.950 338.100 868.050 340.200 ;
        RECT 871.950 339.600 874.050 340.200 ;
        RECT 886.950 339.600 889.050 340.050 ;
        RECT 871.950 338.400 889.050 339.600 ;
        RECT 871.950 338.100 874.050 338.400 ;
        RECT 866.400 334.050 867.600 338.100 ;
        RECT 886.950 337.950 889.050 338.400 ;
        RECT 898.950 338.100 901.050 340.200 ;
        RECT 904.950 339.600 907.050 340.050 ;
        RECT 913.950 339.600 916.050 340.050 ;
        RECT 919.950 339.600 922.050 340.200 ;
        RECT 904.950 338.400 912.600 339.600 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 757.950 333.600 760.050 334.050 ;
        RECT 781.950 333.600 784.050 333.900 ;
        RECT 757.950 333.450 784.050 333.600 ;
        RECT 790.950 333.450 793.050 333.900 ;
        RECT 757.950 332.400 793.050 333.450 ;
        RECT 757.950 331.950 760.050 332.400 ;
        RECT 781.950 332.250 793.050 332.400 ;
        RECT 781.950 331.800 784.050 332.250 ;
        RECT 790.950 331.800 793.050 332.250 ;
        RECT 796.950 333.450 799.050 333.900 ;
        RECT 802.950 333.450 805.050 333.900 ;
        RECT 796.950 332.250 805.050 333.450 ;
        RECT 796.950 331.800 799.050 332.250 ;
        RECT 802.950 331.800 805.050 332.250 ;
        RECT 814.950 333.600 817.050 333.900 ;
        RECT 826.950 333.600 829.050 334.050 ;
        RECT 814.950 332.400 829.050 333.600 ;
        RECT 814.950 331.800 817.050 332.400 ;
        RECT 826.950 331.950 829.050 332.400 ;
        RECT 862.950 332.400 867.600 334.050 ;
        RECT 877.950 333.600 880.050 334.050 ;
        RECT 899.400 333.600 900.600 338.100 ;
        RECT 904.950 337.950 907.050 338.400 ;
        RECT 911.400 336.600 912.600 338.400 ;
        RECT 913.950 338.400 922.050 339.600 ;
        RECT 913.950 337.950 916.050 338.400 ;
        RECT 919.950 338.100 922.050 338.400 ;
        RECT 925.950 338.100 928.050 340.200 ;
        RECT 926.400 336.600 927.600 338.100 ;
        RECT 943.950 336.600 946.050 340.050 ;
        RECT 973.950 339.600 976.050 340.200 ;
        RECT 997.950 339.600 1000.050 340.200 ;
        RECT 973.950 338.400 1000.050 339.600 ;
        RECT 973.950 338.100 976.050 338.400 ;
        RECT 997.950 338.100 1000.050 338.400 ;
        RECT 911.400 335.400 924.600 336.600 ;
        RECT 926.400 336.000 946.050 336.600 ;
        RECT 926.400 335.400 945.600 336.000 ;
        RECT 877.950 332.400 900.600 333.600 ;
        RECT 923.400 333.600 924.600 335.400 ;
        RECT 931.950 333.600 934.050 334.050 ;
        RECT 923.400 332.400 934.050 333.600 ;
        RECT 935.400 333.600 936.600 335.400 ;
        RECT 943.950 333.600 946.050 334.050 ;
        RECT 935.400 332.400 946.050 333.600 ;
        RECT 862.950 331.950 867.000 332.400 ;
        RECT 877.950 331.950 880.050 332.400 ;
        RECT 931.950 331.950 934.050 332.400 ;
        RECT 943.950 331.950 946.050 332.400 ;
        RECT 976.950 333.600 979.050 333.900 ;
        RECT 988.950 333.600 991.050 334.050 ;
        RECT 1001.400 333.900 1002.600 344.400 ;
        RECT 1012.950 344.400 1039.050 345.600 ;
        RECT 1012.950 343.950 1015.050 344.400 ;
        RECT 1036.950 343.950 1039.050 344.400 ;
        RECT 1003.950 339.600 1006.050 340.200 ;
        RECT 1012.950 339.600 1015.050 340.050 ;
        RECT 1003.950 338.400 1015.050 339.600 ;
        RECT 1003.950 338.100 1006.050 338.400 ;
        RECT 1012.950 337.950 1015.050 338.400 ;
        RECT 976.950 332.400 991.050 333.600 ;
        RECT 976.950 331.800 979.050 332.400 ;
        RECT 988.950 331.950 991.050 332.400 ;
        RECT 1000.950 331.800 1003.050 333.900 ;
        RECT 1027.950 333.600 1030.050 333.900 ;
        RECT 1033.950 333.600 1036.050 334.050 ;
        RECT 1039.950 333.600 1042.050 334.050 ;
        RECT 1027.950 332.400 1042.050 333.600 ;
        RECT 1027.950 331.800 1030.050 332.400 ;
        RECT 1033.950 331.950 1036.050 332.400 ;
        RECT 1039.950 331.950 1042.050 332.400 ;
        RECT 4.950 329.400 9.600 330.600 ;
        RECT 226.950 330.600 229.050 331.050 ;
        RECT 553.950 330.600 556.050 331.050 ;
        RECT 565.950 330.600 568.050 331.050 ;
        RECT 226.950 329.400 342.600 330.600 ;
        RECT 4.950 328.800 7.050 329.400 ;
        RECT 226.950 328.950 229.050 329.400 ;
        RECT 341.400 328.050 342.600 329.400 ;
        RECT 553.950 329.400 568.050 330.600 ;
        RECT 553.950 328.950 556.050 329.400 ;
        RECT 565.950 328.950 568.050 329.400 ;
        RECT 577.950 330.600 580.050 331.050 ;
        RECT 613.950 330.600 616.050 331.050 ;
        RECT 577.950 329.400 616.050 330.600 ;
        RECT 577.950 328.950 580.050 329.400 ;
        RECT 613.950 328.950 616.050 329.400 ;
        RECT 646.950 330.600 649.050 331.050 ;
        RECT 679.950 330.600 682.050 331.050 ;
        RECT 646.950 329.400 682.050 330.600 ;
        RECT 646.950 328.950 649.050 329.400 ;
        RECT 679.950 328.950 682.050 329.400 ;
        RECT 718.950 330.600 721.050 331.050 ;
        RECT 742.950 330.600 745.050 331.050 ;
        RECT 754.950 330.600 757.050 331.050 ;
        RECT 718.950 329.400 757.050 330.600 ;
        RECT 718.950 328.950 721.050 329.400 ;
        RECT 742.950 328.950 745.050 329.400 ;
        RECT 754.950 328.950 757.050 329.400 ;
        RECT 844.950 330.600 847.050 331.050 ;
        RECT 892.950 330.600 895.050 331.050 ;
        RECT 844.950 329.400 895.050 330.600 ;
        RECT 844.950 328.950 847.050 329.400 ;
        RECT 892.950 328.950 895.050 329.400 ;
        RECT 94.950 327.600 97.050 328.050 ;
        RECT 220.950 327.600 223.050 328.050 ;
        RECT 94.950 326.400 223.050 327.600 ;
        RECT 94.950 325.950 97.050 326.400 ;
        RECT 220.950 325.950 223.050 326.400 ;
        RECT 247.950 327.600 250.050 328.050 ;
        RECT 259.950 327.600 262.050 328.050 ;
        RECT 247.950 326.400 262.050 327.600 ;
        RECT 247.950 325.950 250.050 326.400 ;
        RECT 259.950 325.950 262.050 326.400 ;
        RECT 301.950 327.600 304.050 328.050 ;
        RECT 325.950 327.600 328.050 328.050 ;
        RECT 301.950 326.400 328.050 327.600 ;
        RECT 301.950 325.950 304.050 326.400 ;
        RECT 325.950 325.950 328.050 326.400 ;
        RECT 340.950 327.600 343.050 328.050 ;
        RECT 358.950 327.600 361.050 328.050 ;
        RECT 340.950 326.400 361.050 327.600 ;
        RECT 340.950 325.950 343.050 326.400 ;
        RECT 358.950 325.950 361.050 326.400 ;
        RECT 433.950 327.600 436.050 328.050 ;
        RECT 451.950 327.600 454.050 328.050 ;
        RECT 433.950 326.400 454.050 327.600 ;
        RECT 433.950 325.950 436.050 326.400 ;
        RECT 451.950 325.950 454.050 326.400 ;
        RECT 487.950 327.600 490.050 328.050 ;
        RECT 511.950 327.600 514.050 328.050 ;
        RECT 541.950 327.600 544.050 328.050 ;
        RECT 487.950 326.400 544.050 327.600 ;
        RECT 487.950 325.950 490.050 326.400 ;
        RECT 511.950 325.950 514.050 326.400 ;
        RECT 541.950 325.950 544.050 326.400 ;
        RECT 631.950 327.600 634.050 328.050 ;
        RECT 709.950 327.600 712.050 328.050 ;
        RECT 631.950 326.400 712.050 327.600 ;
        RECT 631.950 325.950 634.050 326.400 ;
        RECT 709.950 325.950 712.050 326.400 ;
        RECT 826.950 327.600 829.050 328.050 ;
        RECT 856.950 327.600 859.050 328.050 ;
        RECT 826.950 326.400 859.050 327.600 ;
        RECT 826.950 325.950 829.050 326.400 ;
        RECT 856.950 325.950 859.050 326.400 ;
        RECT 886.950 327.600 889.050 328.050 ;
        RECT 901.950 327.600 904.050 328.050 ;
        RECT 886.950 326.400 904.050 327.600 ;
        RECT 886.950 325.950 889.050 326.400 ;
        RECT 901.950 325.950 904.050 326.400 ;
        RECT 106.950 324.600 109.050 325.050 ;
        RECT 136.950 324.600 139.050 325.050 ;
        RECT 106.950 323.400 139.050 324.600 ;
        RECT 106.950 322.950 109.050 323.400 ;
        RECT 136.950 322.950 139.050 323.400 ;
        RECT 262.950 324.600 265.050 325.050 ;
        RECT 289.950 324.600 292.050 325.050 ;
        RECT 262.950 323.400 292.050 324.600 ;
        RECT 262.950 322.950 265.050 323.400 ;
        RECT 289.950 322.950 292.050 323.400 ;
        RECT 442.950 324.600 445.050 325.050 ;
        RECT 463.950 324.600 466.050 325.050 ;
        RECT 442.950 323.400 466.050 324.600 ;
        RECT 442.950 322.950 445.050 323.400 ;
        RECT 463.950 322.950 466.050 323.400 ;
        RECT 619.950 324.600 622.050 325.050 ;
        RECT 628.950 324.600 631.050 325.050 ;
        RECT 619.950 323.400 631.050 324.600 ;
        RECT 619.950 322.950 622.050 323.400 ;
        RECT 628.950 322.950 631.050 323.400 ;
        RECT 679.950 324.600 682.050 325.050 ;
        RECT 823.950 324.600 826.050 325.050 ;
        RECT 679.950 323.400 826.050 324.600 ;
        RECT 679.950 322.950 682.050 323.400 ;
        RECT 823.950 322.950 826.050 323.400 ;
        RECT 835.950 324.600 838.050 325.050 ;
        RECT 853.950 324.600 856.050 325.050 ;
        RECT 835.950 323.400 856.050 324.600 ;
        RECT 835.950 322.950 838.050 323.400 ;
        RECT 853.950 322.950 856.050 323.400 ;
        RECT 874.950 324.600 877.050 325.050 ;
        RECT 913.950 324.600 916.050 325.050 ;
        RECT 874.950 323.400 916.050 324.600 ;
        RECT 874.950 322.950 877.050 323.400 ;
        RECT 913.950 322.950 916.050 323.400 ;
        RECT 196.950 321.600 199.050 322.050 ;
        RECT 223.950 321.600 226.050 322.050 ;
        RECT 196.950 320.400 226.050 321.600 ;
        RECT 196.950 319.950 199.050 320.400 ;
        RECT 223.950 319.950 226.050 320.400 ;
        RECT 322.950 321.600 325.050 322.050 ;
        RECT 337.950 321.600 340.050 322.050 ;
        RECT 322.950 320.400 340.050 321.600 ;
        RECT 322.950 319.950 325.050 320.400 ;
        RECT 337.950 319.950 340.050 320.400 ;
        RECT 379.950 321.600 382.050 322.050 ;
        RECT 595.950 321.600 598.050 322.050 ;
        RECT 643.950 321.600 646.050 322.050 ;
        RECT 667.950 321.600 670.050 322.050 ;
        RECT 379.950 320.400 670.050 321.600 ;
        RECT 379.950 319.950 382.050 320.400 ;
        RECT 595.950 319.950 598.050 320.400 ;
        RECT 643.950 319.950 646.050 320.400 ;
        RECT 667.950 319.950 670.050 320.400 ;
        RECT 802.950 321.600 805.050 322.050 ;
        RECT 832.950 321.600 835.050 322.050 ;
        RECT 802.950 320.400 835.050 321.600 ;
        RECT 802.950 319.950 805.050 320.400 ;
        RECT 832.950 319.950 835.050 320.400 ;
        RECT 910.950 321.600 913.050 322.050 ;
        RECT 916.950 321.600 919.050 322.050 ;
        RECT 976.950 321.600 979.050 322.050 ;
        RECT 910.950 320.400 979.050 321.600 ;
        RECT 910.950 319.950 913.050 320.400 ;
        RECT 916.950 319.950 919.050 320.400 ;
        RECT 976.950 319.950 979.050 320.400 ;
        RECT 70.950 318.600 73.050 319.050 ;
        RECT 85.950 318.600 88.050 319.050 ;
        RECT 70.950 317.400 88.050 318.600 ;
        RECT 70.950 316.950 73.050 317.400 ;
        RECT 85.950 316.950 88.050 317.400 ;
        RECT 238.950 318.600 241.050 319.050 ;
        RECT 463.950 318.600 466.050 319.050 ;
        RECT 559.950 318.600 562.050 319.050 ;
        RECT 592.950 318.600 595.050 319.050 ;
        RECT 238.950 317.400 336.600 318.600 ;
        RECT 238.950 316.950 241.050 317.400 ;
        RECT 61.950 315.600 64.050 316.050 ;
        RECT 112.950 315.600 115.050 316.050 ;
        RECT 61.950 314.400 115.050 315.600 ;
        RECT 61.950 313.950 64.050 314.400 ;
        RECT 112.950 313.950 115.050 314.400 ;
        RECT 181.950 315.600 184.050 316.050 ;
        RECT 196.950 315.600 199.050 316.050 ;
        RECT 181.950 314.400 199.050 315.600 ;
        RECT 181.950 313.950 184.050 314.400 ;
        RECT 196.950 313.950 199.050 314.400 ;
        RECT 220.950 315.600 223.050 316.050 ;
        RECT 313.950 315.600 316.050 316.050 ;
        RECT 328.950 315.600 331.050 316.050 ;
        RECT 220.950 314.400 331.050 315.600 ;
        RECT 335.400 315.600 336.600 317.400 ;
        RECT 463.950 317.400 595.050 318.600 ;
        RECT 463.950 316.950 466.050 317.400 ;
        RECT 559.950 316.950 562.050 317.400 ;
        RECT 592.950 316.950 595.050 317.400 ;
        RECT 613.950 318.600 616.050 319.050 ;
        RECT 727.950 318.600 730.050 319.050 ;
        RECT 613.950 317.400 730.050 318.600 ;
        RECT 613.950 316.950 616.050 317.400 ;
        RECT 727.950 316.950 730.050 317.400 ;
        RECT 763.950 318.600 766.050 319.050 ;
        RECT 823.950 318.600 826.050 319.050 ;
        RECT 763.950 317.400 826.050 318.600 ;
        RECT 763.950 316.950 766.050 317.400 ;
        RECT 823.950 316.950 826.050 317.400 ;
        RECT 841.950 318.600 844.050 319.050 ;
        RECT 895.950 318.600 898.050 319.050 ;
        RECT 937.950 318.600 940.050 319.050 ;
        RECT 841.950 317.400 940.050 318.600 ;
        RECT 841.950 316.950 844.050 317.400 ;
        RECT 895.950 316.950 898.050 317.400 ;
        RECT 937.950 316.950 940.050 317.400 ;
        RECT 988.950 318.600 991.050 319.050 ;
        RECT 1036.950 318.600 1039.050 319.050 ;
        RECT 988.950 317.400 1039.050 318.600 ;
        RECT 988.950 316.950 991.050 317.400 ;
        RECT 1036.950 316.950 1039.050 317.400 ;
        RECT 343.950 315.600 346.050 316.050 ;
        RECT 335.400 314.400 346.050 315.600 ;
        RECT 220.950 313.950 223.050 314.400 ;
        RECT 313.950 313.950 316.050 314.400 ;
        RECT 328.950 313.950 331.050 314.400 ;
        RECT 343.950 313.950 346.050 314.400 ;
        RECT 472.950 315.600 475.050 316.050 ;
        RECT 514.950 315.600 517.050 316.050 ;
        RECT 472.950 314.400 517.050 315.600 ;
        RECT 472.950 313.950 475.050 314.400 ;
        RECT 514.950 313.950 517.050 314.400 ;
        RECT 628.950 315.600 631.050 316.050 ;
        RECT 679.950 315.600 682.050 316.050 ;
        RECT 628.950 314.400 682.050 315.600 ;
        RECT 628.950 313.950 631.050 314.400 ;
        RECT 679.950 313.950 682.050 314.400 ;
        RECT 760.950 315.600 763.050 316.050 ;
        RECT 826.800 315.600 828.900 316.050 ;
        RECT 760.950 314.400 828.900 315.600 ;
        RECT 760.950 313.950 763.050 314.400 ;
        RECT 826.800 313.950 828.900 314.400 ;
        RECT 871.950 315.600 874.050 316.050 ;
        RECT 880.950 315.600 883.050 316.050 ;
        RECT 871.950 314.400 883.050 315.600 ;
        RECT 871.950 313.950 874.050 314.400 ;
        RECT 880.950 313.950 883.050 314.400 ;
        RECT 919.950 315.600 922.050 316.050 ;
        RECT 934.950 315.600 937.050 316.050 ;
        RECT 919.950 314.400 937.050 315.600 ;
        RECT 919.950 313.950 922.050 314.400 ;
        RECT 934.950 313.950 937.050 314.400 ;
        RECT 970.950 315.600 973.050 316.050 ;
        RECT 1012.950 315.600 1015.050 316.050 ;
        RECT 970.950 314.400 1015.050 315.600 ;
        RECT 970.950 313.950 973.050 314.400 ;
        RECT 1012.950 313.950 1015.050 314.400 ;
        RECT 694.950 312.600 697.050 313.050 ;
        RECT 730.950 312.600 733.050 313.050 ;
        RECT 694.950 311.400 733.050 312.600 ;
        RECT 694.950 310.950 697.050 311.400 ;
        RECT 730.950 310.950 733.050 311.400 ;
        RECT 775.950 312.600 778.050 313.050 ;
        RECT 841.950 312.600 844.050 313.050 ;
        RECT 775.950 311.400 844.050 312.600 ;
        RECT 775.950 310.950 778.050 311.400 ;
        RECT 841.950 310.950 844.050 311.400 ;
        RECT 862.950 312.600 865.050 313.050 ;
        RECT 922.950 312.600 925.050 313.050 ;
        RECT 1009.950 312.600 1012.050 313.050 ;
        RECT 862.950 311.400 1012.050 312.600 ;
        RECT 862.950 310.950 865.050 311.400 ;
        RECT 922.950 310.950 925.050 311.400 ;
        RECT 1009.950 310.950 1012.050 311.400 ;
        RECT 118.950 309.600 121.050 310.050 ;
        RECT 226.950 309.600 229.050 310.050 ;
        RECT 118.950 308.400 229.050 309.600 ;
        RECT 118.950 307.950 121.050 308.400 ;
        RECT 226.950 307.950 229.050 308.400 ;
        RECT 244.950 309.600 247.050 310.050 ;
        RECT 277.950 309.600 280.050 310.050 ;
        RECT 244.950 308.400 280.050 309.600 ;
        RECT 244.950 307.950 247.050 308.400 ;
        RECT 277.950 307.950 280.050 308.400 ;
        RECT 505.950 309.600 508.050 310.050 ;
        RECT 601.950 309.600 604.050 310.050 ;
        RECT 505.950 308.400 604.050 309.600 ;
        RECT 505.950 307.950 508.050 308.400 ;
        RECT 601.950 307.950 604.050 308.400 ;
        RECT 607.950 309.600 610.050 310.050 ;
        RECT 646.950 309.600 649.050 310.050 ;
        RECT 607.950 308.400 649.050 309.600 ;
        RECT 607.950 307.950 610.050 308.400 ;
        RECT 646.950 307.950 649.050 308.400 ;
        RECT 838.950 309.600 841.050 310.050 ;
        RECT 919.950 309.600 922.050 310.050 ;
        RECT 838.950 308.400 922.050 309.600 ;
        RECT 838.950 307.950 841.050 308.400 ;
        RECT 919.950 307.950 922.050 308.400 ;
        RECT 937.950 309.600 940.050 310.050 ;
        RECT 943.950 309.600 946.050 310.050 ;
        RECT 937.950 308.400 946.050 309.600 ;
        RECT 937.950 307.950 940.050 308.400 ;
        RECT 943.950 307.950 946.050 308.400 ;
        RECT 964.950 309.600 967.050 310.050 ;
        RECT 979.950 309.600 982.050 310.050 ;
        RECT 964.950 308.400 982.050 309.600 ;
        RECT 964.950 307.950 967.050 308.400 ;
        RECT 979.950 307.950 982.050 308.400 ;
        RECT 64.950 306.600 67.050 307.050 ;
        RECT 73.950 306.600 76.050 307.050 ;
        RECT 64.950 305.400 76.050 306.600 ;
        RECT 64.950 304.950 67.050 305.400 ;
        RECT 73.950 304.950 76.050 305.400 ;
        RECT 379.950 306.600 382.050 307.050 ;
        RECT 427.950 306.600 430.050 307.050 ;
        RECT 379.950 305.400 430.050 306.600 ;
        RECT 379.950 304.950 382.050 305.400 ;
        RECT 427.950 304.950 430.050 305.400 ;
        RECT 583.950 306.600 586.050 307.050 ;
        RECT 628.950 306.600 631.050 307.050 ;
        RECT 583.950 305.400 631.050 306.600 ;
        RECT 583.950 304.950 586.050 305.400 ;
        RECT 628.950 304.950 631.050 305.400 ;
        RECT 682.950 306.600 685.050 307.050 ;
        RECT 754.950 306.600 757.050 307.050 ;
        RECT 763.950 306.600 766.050 307.050 ;
        RECT 682.950 305.400 766.050 306.600 ;
        RECT 682.950 304.950 685.050 305.400 ;
        RECT 754.950 304.950 757.050 305.400 ;
        RECT 763.950 304.950 766.050 305.400 ;
        RECT 808.950 306.600 811.050 307.050 ;
        RECT 839.400 306.600 840.600 307.950 ;
        RECT 808.950 305.400 840.600 306.600 ;
        RECT 928.950 306.600 931.050 307.050 ;
        RECT 946.950 306.600 949.050 307.050 ;
        RECT 991.950 306.600 994.050 307.050 ;
        RECT 928.950 305.400 994.050 306.600 ;
        RECT 808.950 304.950 811.050 305.400 ;
        RECT 928.950 304.950 931.050 305.400 ;
        RECT 946.950 304.950 949.050 305.400 ;
        RECT 991.950 304.950 994.050 305.400 ;
        RECT 1009.950 306.600 1012.050 307.050 ;
        RECT 1015.950 306.600 1018.050 307.050 ;
        RECT 1027.950 306.600 1030.050 307.050 ;
        RECT 1009.950 305.400 1030.050 306.600 ;
        RECT 1009.950 304.950 1012.050 305.400 ;
        RECT 1015.950 304.950 1018.050 305.400 ;
        RECT 1027.950 304.950 1030.050 305.400 ;
        RECT 154.950 303.600 157.050 304.050 ;
        RECT 253.950 303.600 256.050 304.050 ;
        RECT 154.950 302.400 256.050 303.600 ;
        RECT 154.950 301.950 157.050 302.400 ;
        RECT 253.950 301.950 256.050 302.400 ;
        RECT 661.950 303.600 664.050 304.050 ;
        RECT 760.950 303.600 763.050 304.050 ;
        RECT 661.950 302.400 763.050 303.600 ;
        RECT 661.950 301.950 664.050 302.400 ;
        RECT 760.950 301.950 763.050 302.400 ;
        RECT 889.950 303.600 892.050 304.050 ;
        RECT 916.950 303.600 919.050 304.050 ;
        RECT 889.950 302.400 919.050 303.600 ;
        RECT 889.950 301.950 892.050 302.400 ;
        RECT 916.950 301.950 919.050 302.400 ;
        RECT 76.950 300.600 79.050 301.050 ;
        RECT 100.950 300.600 103.050 301.050 ;
        RECT 76.950 299.400 103.050 300.600 ;
        RECT 76.950 298.950 79.050 299.400 ;
        RECT 100.950 298.950 103.050 299.400 ;
        RECT 220.950 300.600 223.050 301.050 ;
        RECT 232.950 300.600 235.050 301.050 ;
        RECT 220.950 299.400 235.050 300.600 ;
        RECT 220.950 298.950 223.050 299.400 ;
        RECT 232.950 298.950 235.050 299.400 ;
        RECT 256.950 300.600 259.050 301.050 ;
        RECT 292.950 300.600 295.050 301.050 ;
        RECT 256.950 299.400 295.050 300.600 ;
        RECT 256.950 298.950 259.050 299.400 ;
        RECT 292.950 298.950 295.050 299.400 ;
        RECT 361.950 300.600 364.050 301.050 ;
        RECT 409.950 300.600 412.050 301.050 ;
        RECT 361.950 299.400 412.050 300.600 ;
        RECT 361.950 298.950 364.050 299.400 ;
        RECT 409.950 298.950 412.050 299.400 ;
        RECT 424.950 300.600 427.050 301.050 ;
        RECT 442.950 300.600 445.050 301.050 ;
        RECT 424.950 299.400 445.050 300.600 ;
        RECT 424.950 298.950 427.050 299.400 ;
        RECT 442.950 298.950 445.050 299.400 ;
        RECT 544.950 300.600 547.050 301.050 ;
        RECT 586.950 300.600 589.050 301.050 ;
        RECT 544.950 299.400 589.050 300.600 ;
        RECT 544.950 298.950 547.050 299.400 ;
        RECT 586.950 298.950 589.050 299.400 ;
        RECT 676.950 300.600 679.050 301.050 ;
        RECT 691.950 300.600 694.050 301.050 ;
        RECT 676.950 299.400 694.050 300.600 ;
        RECT 676.950 298.950 679.050 299.400 ;
        RECT 691.950 298.950 694.050 299.400 ;
        RECT 772.950 300.600 775.050 301.050 ;
        RECT 805.950 300.600 808.050 301.050 ;
        RECT 772.950 299.400 808.050 300.600 ;
        RECT 772.950 298.950 775.050 299.400 ;
        RECT 805.950 298.950 808.050 299.400 ;
        RECT 922.950 300.600 925.050 301.050 ;
        RECT 967.950 300.600 970.050 300.900 ;
        RECT 922.950 299.400 970.050 300.600 ;
        RECT 922.950 298.950 925.050 299.400 ;
        RECT 967.950 298.800 970.050 299.400 ;
        RECT 979.950 300.600 982.050 301.050 ;
        RECT 1015.950 300.600 1018.050 301.050 ;
        RECT 979.950 299.400 1018.050 300.600 ;
        RECT 979.950 298.950 982.050 299.400 ;
        RECT 1015.950 298.950 1018.050 299.400 ;
        RECT 235.950 297.600 238.050 298.050 ;
        RECT 241.950 297.600 244.050 298.050 ;
        RECT 235.950 296.400 244.050 297.600 ;
        RECT 235.950 295.950 238.050 296.400 ;
        RECT 241.950 295.950 244.050 296.400 ;
        RECT 271.950 297.600 274.050 297.900 ;
        RECT 307.950 297.600 310.050 298.050 ;
        RECT 271.950 296.400 310.050 297.600 ;
        RECT 271.950 295.800 274.050 296.400 ;
        RECT 307.950 295.950 310.050 296.400 ;
        RECT 451.950 297.750 454.050 298.200 ;
        RECT 460.950 297.750 463.050 298.200 ;
        RECT 451.950 297.600 463.050 297.750 ;
        RECT 520.950 297.600 523.050 298.200 ;
        RECT 451.950 296.550 501.600 297.600 ;
        RECT 451.950 296.100 454.050 296.550 ;
        RECT 460.950 296.400 501.600 296.550 ;
        RECT 460.950 296.100 463.050 296.400 ;
        RECT 16.950 293.100 19.050 295.200 ;
        RECT 22.950 293.100 25.050 295.200 ;
        RECT 37.950 294.750 40.050 295.200 ;
        RECT 43.950 294.750 46.050 295.200 ;
        RECT 37.950 293.550 46.050 294.750 ;
        RECT 37.950 293.100 40.050 293.550 ;
        RECT 43.950 293.100 46.050 293.550 ;
        RECT 49.950 293.100 52.050 295.200 ;
        RECT 70.950 293.100 73.050 295.200 ;
        RECT 88.950 294.750 91.050 295.200 ;
        RECT 94.950 294.750 97.050 295.200 ;
        RECT 88.950 293.550 97.050 294.750 ;
        RECT 88.950 293.100 91.050 293.550 ;
        RECT 94.950 293.100 97.050 293.550 ;
        RECT 112.950 294.750 115.050 295.200 ;
        RECT 124.950 294.750 127.050 295.200 ;
        RECT 112.950 293.550 127.050 294.750 ;
        RECT 112.950 293.100 115.050 293.550 ;
        RECT 124.950 293.100 127.050 293.550 ;
        RECT 130.950 293.100 133.050 295.200 ;
        RECT 178.950 293.100 181.050 295.200 ;
        RECT 184.950 294.600 187.050 295.200 ;
        RECT 205.950 294.600 208.050 295.200 ;
        RECT 211.950 294.600 214.050 295.050 ;
        RECT 184.950 293.400 214.050 294.600 ;
        RECT 184.950 293.100 187.050 293.400 ;
        RECT 205.950 293.100 208.050 293.400 ;
        RECT 17.400 289.050 18.600 293.100 ;
        RECT 13.950 287.400 18.600 289.050 ;
        RECT 13.950 286.950 18.000 287.400 ;
        RECT 23.400 286.050 24.600 293.100 ;
        RECT 25.950 288.600 28.050 288.900 ;
        RECT 37.950 288.600 40.050 289.050 ;
        RECT 25.950 287.400 40.050 288.600 ;
        RECT 25.950 286.800 28.050 287.400 ;
        RECT 37.950 286.950 40.050 287.400 ;
        RECT 22.950 283.950 25.050 286.050 ;
        RECT 43.950 285.600 46.050 286.050 ;
        RECT 50.400 285.600 51.600 293.100 ;
        RECT 71.400 291.600 72.600 293.100 ;
        RECT 56.400 290.400 72.600 291.600 ;
        RECT 131.400 291.600 132.600 293.100 ;
        RECT 131.400 290.400 138.600 291.600 ;
        RECT 52.950 288.600 55.050 288.900 ;
        RECT 56.400 288.600 57.600 290.400 ;
        RECT 52.950 287.400 57.600 288.600 ;
        RECT 58.950 288.600 61.050 289.050 ;
        RECT 73.950 288.600 76.050 288.900 ;
        RECT 58.950 287.400 76.050 288.600 ;
        RECT 52.950 286.800 55.050 287.400 ;
        RECT 58.950 286.950 61.050 287.400 ;
        RECT 73.950 286.800 76.050 287.400 ;
        RECT 103.950 288.450 106.050 288.900 ;
        RECT 118.950 288.450 121.050 288.900 ;
        RECT 103.950 287.250 121.050 288.450 ;
        RECT 137.400 288.600 138.600 290.400 ;
        RECT 175.950 288.600 178.050 288.900 ;
        RECT 137.400 287.400 178.050 288.600 ;
        RECT 103.950 286.800 106.050 287.250 ;
        RECT 118.950 286.800 121.050 287.250 ;
        RECT 175.950 286.800 178.050 287.400 ;
        RECT 43.950 284.400 51.600 285.600 ;
        RECT 133.950 285.600 136.050 286.050 ;
        RECT 157.950 285.600 160.050 286.050 ;
        RECT 133.950 284.400 160.050 285.600 ;
        RECT 43.950 283.950 46.050 284.400 ;
        RECT 133.950 283.950 136.050 284.400 ;
        RECT 157.950 283.950 160.050 284.400 ;
        RECT 179.400 283.050 180.600 293.100 ;
        RECT 211.950 292.950 214.050 293.400 ;
        RECT 232.950 294.750 235.050 295.200 ;
        RECT 265.950 294.750 268.050 295.200 ;
        RECT 232.950 293.550 268.050 294.750 ;
        RECT 232.950 293.100 235.050 293.550 ;
        RECT 265.950 293.100 268.050 293.550 ;
        RECT 301.950 294.750 304.050 295.200 ;
        RECT 316.950 294.750 319.050 295.200 ;
        RECT 301.950 293.550 319.050 294.750 ;
        RECT 301.950 293.100 304.050 293.550 ;
        RECT 316.950 293.100 319.050 293.550 ;
        RECT 334.950 294.600 337.050 295.200 ;
        RECT 346.950 294.600 349.050 295.050 ;
        RECT 352.950 294.600 355.050 295.200 ;
        RECT 334.950 293.400 355.050 294.600 ;
        RECT 334.950 293.100 337.050 293.400 ;
        RECT 346.950 292.950 349.050 293.400 ;
        RECT 352.950 293.100 355.050 293.400 ;
        RECT 367.950 294.600 370.050 295.050 ;
        RECT 376.950 294.600 379.050 295.200 ;
        RECT 367.950 293.400 379.050 294.600 ;
        RECT 500.400 294.600 501.600 296.400 ;
        RECT 515.400 296.400 523.050 297.600 ;
        RECT 515.400 294.600 516.600 296.400 ;
        RECT 520.950 296.100 523.050 296.400 ;
        RECT 565.950 297.600 568.050 298.050 ;
        RECT 607.950 297.600 610.050 298.050 ;
        RECT 565.950 296.400 610.050 297.600 ;
        RECT 565.950 295.950 568.050 296.400 ;
        RECT 607.950 295.950 610.050 296.400 ;
        RECT 637.950 297.600 640.050 298.050 ;
        RECT 646.950 297.600 649.050 298.050 ;
        RECT 703.950 297.600 706.050 298.050 ;
        RECT 637.950 296.400 649.050 297.600 ;
        RECT 637.950 295.950 640.050 296.400 ;
        RECT 646.950 295.950 649.050 296.400 ;
        RECT 659.400 296.400 706.050 297.600 ;
        RECT 610.950 294.600 613.050 295.200 ;
        RECT 500.400 293.400 516.600 294.600 ;
        RECT 581.400 293.400 613.050 294.600 ;
        RECT 367.950 292.950 370.050 293.400 ;
        RECT 376.950 293.100 379.050 293.400 ;
        RECT 394.950 291.600 397.050 292.050 ;
        RECT 424.950 291.600 427.050 292.050 ;
        RECT 394.950 290.400 427.050 291.600 ;
        RECT 394.950 289.950 397.050 290.400 ;
        RECT 424.950 289.950 427.050 290.400 ;
        RECT 475.950 291.750 478.050 292.200 ;
        RECT 517.950 291.750 520.050 292.200 ;
        RECT 581.400 291.900 582.600 293.400 ;
        RECT 610.950 293.100 613.050 293.400 ;
        RECT 622.950 294.750 625.050 295.200 ;
        RECT 628.950 294.750 631.050 295.200 ;
        RECT 622.950 293.550 631.050 294.750 ;
        RECT 622.950 293.100 625.050 293.550 ;
        RECT 628.950 293.100 631.050 293.550 ;
        RECT 634.950 294.750 637.050 295.200 ;
        RECT 649.950 294.750 652.050 295.200 ;
        RECT 634.950 294.600 652.050 294.750 ;
        RECT 659.400 294.600 660.600 296.400 ;
        RECT 634.950 293.550 660.600 294.600 ;
        RECT 634.950 293.100 637.050 293.550 ;
        RECT 649.950 293.400 660.600 293.550 ;
        RECT 664.950 294.600 667.050 295.200 ;
        RECT 689.400 295.050 690.600 296.400 ;
        RECT 703.950 295.950 706.050 296.400 ;
        RECT 709.950 297.600 712.050 298.050 ;
        RECT 715.950 297.600 718.050 298.050 ;
        RECT 709.950 296.400 718.050 297.600 ;
        RECT 709.950 295.950 712.050 296.400 ;
        RECT 715.950 295.950 718.050 296.400 ;
        RECT 766.950 297.600 769.050 298.050 ;
        RECT 775.950 297.600 778.050 298.050 ;
        RECT 766.950 296.400 778.050 297.600 ;
        RECT 766.950 295.950 769.050 296.400 ;
        RECT 775.950 295.950 778.050 296.400 ;
        RECT 808.950 295.950 811.050 298.050 ;
        RECT 817.950 297.750 820.050 298.200 ;
        RECT 865.950 297.750 868.050 298.200 ;
        RECT 817.950 296.550 868.050 297.750 ;
        RECT 817.950 296.100 820.050 296.550 ;
        RECT 865.950 296.100 868.050 296.550 ;
        RECT 892.950 297.600 895.050 298.050 ;
        RECT 907.950 297.600 910.050 297.900 ;
        RECT 892.950 296.400 910.050 297.600 ;
        RECT 892.950 295.950 895.050 296.400 ;
        RECT 673.950 294.600 676.050 295.050 ;
        RECT 664.950 293.400 676.050 294.600 ;
        RECT 649.950 293.100 652.050 293.400 ;
        RECT 664.950 293.100 667.050 293.400 ;
        RECT 673.950 292.950 676.050 293.400 ;
        RECT 688.950 292.950 691.050 295.050 ;
        RECT 757.800 292.950 759.900 295.050 ;
        RECT 760.950 294.600 763.050 295.200 ;
        RECT 781.950 294.600 784.050 295.050 ;
        RECT 760.950 293.400 784.050 294.600 ;
        RECT 760.950 293.100 763.050 293.400 ;
        RECT 781.950 292.950 784.050 293.400 ;
        RECT 799.950 293.100 802.050 295.200 ;
        RECT 475.950 290.550 520.050 291.750 ;
        RECT 475.950 290.100 478.050 290.550 ;
        RECT 517.950 290.100 520.050 290.550 ;
        RECT 580.950 289.800 583.050 291.900 ;
        RECT 699.000 291.600 703.050 292.050 ;
        RECT 698.400 289.950 703.050 291.600 ;
        RECT 223.950 288.600 226.050 289.050 ;
        RECT 250.950 288.600 253.050 289.050 ;
        RECT 223.950 287.400 253.050 288.600 ;
        RECT 223.950 286.950 226.050 287.400 ;
        RECT 250.950 286.950 253.050 287.400 ;
        RECT 256.950 288.600 259.050 288.900 ;
        RECT 271.950 288.600 274.050 289.050 ;
        RECT 256.950 287.400 274.050 288.600 ;
        RECT 256.950 286.800 259.050 287.400 ;
        RECT 271.950 286.950 274.050 287.400 ;
        RECT 316.950 288.600 319.050 289.050 ;
        RECT 331.950 288.600 334.050 288.900 ;
        RECT 316.950 287.400 334.050 288.600 ;
        RECT 316.950 286.950 319.050 287.400 ;
        RECT 331.950 286.800 334.050 287.400 ;
        RECT 595.950 288.450 598.050 288.900 ;
        RECT 601.950 288.450 604.050 288.900 ;
        RECT 595.950 287.250 604.050 288.450 ;
        RECT 595.950 286.800 598.050 287.250 ;
        RECT 601.950 286.800 604.050 287.250 ;
        RECT 607.950 288.600 610.050 288.900 ;
        RECT 622.950 288.600 625.050 289.050 ;
        RECT 607.950 287.400 625.050 288.600 ;
        RECT 607.950 286.800 610.050 287.400 ;
        RECT 622.950 286.950 625.050 287.400 ;
        RECT 637.950 288.450 640.050 288.900 ;
        RECT 646.950 288.450 649.050 288.900 ;
        RECT 637.950 287.250 649.050 288.450 ;
        RECT 637.950 286.800 640.050 287.250 ;
        RECT 646.950 286.800 649.050 287.250 ;
        RECT 661.950 288.600 664.050 288.900 ;
        RECT 698.400 288.600 699.600 289.950 ;
        RECT 661.950 287.400 699.600 288.600 ;
        RECT 727.950 288.450 730.050 288.900 ;
        RECT 736.950 288.450 739.050 288.900 ;
        RECT 661.950 286.800 664.050 287.400 ;
        RECT 727.950 287.250 739.050 288.450 ;
        RECT 758.250 288.600 759.450 292.950 ;
        RECT 775.950 291.600 778.050 292.050 ;
        RECT 800.400 291.600 801.600 293.100 ;
        RECT 775.950 290.400 801.600 291.600 ;
        RECT 805.950 291.600 808.050 291.900 ;
        RECT 809.400 291.600 810.600 295.950 ;
        RECT 907.950 295.800 910.050 296.400 ;
        RECT 841.950 294.600 844.050 295.050 ;
        RECT 856.950 294.600 859.050 295.050 ;
        RECT 841.950 293.400 859.050 294.600 ;
        RECT 841.950 292.950 844.050 293.400 ;
        RECT 856.950 292.950 859.050 293.400 ;
        RECT 898.950 294.600 901.050 295.050 ;
        RECT 910.950 294.600 913.050 295.050 ;
        RECT 940.950 294.750 943.050 295.200 ;
        RECT 970.950 294.750 973.050 295.200 ;
        RECT 940.950 294.600 973.050 294.750 ;
        RECT 898.950 293.400 906.600 294.600 ;
        RECT 898.950 292.950 901.050 293.400 ;
        RECT 805.950 290.400 810.600 291.600 ;
        RECT 905.400 291.600 906.600 293.400 ;
        RECT 910.950 293.550 973.050 294.600 ;
        RECT 910.950 293.400 943.050 293.550 ;
        RECT 910.950 292.950 913.050 293.400 ;
        RECT 940.950 293.100 943.050 293.400 ;
        RECT 970.950 293.100 973.050 293.550 ;
        RECT 1021.950 294.750 1024.050 295.200 ;
        RECT 1033.950 294.750 1036.050 295.200 ;
        RECT 1021.950 293.550 1036.050 294.750 ;
        RECT 1021.950 293.100 1024.050 293.550 ;
        RECT 1033.950 293.100 1036.050 293.550 ;
        RECT 905.400 290.400 915.600 291.600 ;
        RECT 775.950 289.950 778.050 290.400 ;
        RECT 805.950 289.800 808.050 290.400 ;
        RECT 914.400 288.900 915.600 290.400 ;
        RECT 763.950 288.600 766.050 288.900 ;
        RECT 758.250 287.400 766.050 288.600 ;
        RECT 727.950 286.800 730.050 287.250 ;
        RECT 736.950 286.800 739.050 287.250 ;
        RECT 763.950 286.800 766.050 287.400 ;
        RECT 913.950 286.800 916.050 288.900 ;
        RECT 934.950 288.450 937.050 288.900 ;
        RECT 955.950 288.600 958.050 288.900 ;
        RECT 961.950 288.600 964.050 289.050 ;
        RECT 955.950 288.450 964.050 288.600 ;
        RECT 934.950 287.400 964.050 288.450 ;
        RECT 934.950 287.250 958.050 287.400 ;
        RECT 934.950 286.800 937.050 287.250 ;
        RECT 955.950 286.800 958.050 287.250 ;
        RECT 961.950 286.950 964.050 287.400 ;
        RECT 1006.950 288.450 1009.050 288.900 ;
        RECT 1024.950 288.450 1027.050 288.900 ;
        RECT 1006.950 287.250 1027.050 288.450 ;
        RECT 1006.950 286.800 1009.050 287.250 ;
        RECT 1024.950 286.800 1027.050 287.250 ;
        RECT 235.950 285.600 238.050 286.050 ;
        RECT 283.950 285.600 286.050 286.050 ;
        RECT 235.950 284.400 286.050 285.600 ;
        RECT 235.950 283.950 238.050 284.400 ;
        RECT 283.950 283.950 286.050 284.400 ;
        RECT 310.950 285.600 313.050 286.050 ;
        RECT 322.950 285.600 325.050 286.050 ;
        RECT 310.950 284.400 325.050 285.600 ;
        RECT 310.950 283.950 313.050 284.400 ;
        RECT 322.950 283.950 325.050 284.400 ;
        RECT 346.950 285.600 349.050 286.050 ;
        RECT 373.950 285.600 376.050 286.050 ;
        RECT 346.950 284.400 376.050 285.600 ;
        RECT 346.950 283.950 349.050 284.400 ;
        RECT 373.950 283.950 376.050 284.400 ;
        RECT 514.950 285.600 517.050 286.050 ;
        RECT 568.950 285.600 571.050 286.050 ;
        RECT 514.950 284.400 571.050 285.600 ;
        RECT 514.950 283.950 517.050 284.400 ;
        RECT 568.950 283.950 571.050 284.400 ;
        RECT 766.950 285.600 769.050 286.050 ;
        RECT 775.950 285.600 778.050 286.050 ;
        RECT 766.950 284.400 778.050 285.600 ;
        RECT 766.950 283.950 769.050 284.400 ;
        RECT 775.950 283.950 778.050 284.400 ;
        RECT 868.950 285.600 871.050 286.050 ;
        RECT 877.950 285.600 880.050 286.050 ;
        RECT 868.950 284.400 880.050 285.600 ;
        RECT 868.950 283.950 871.050 284.400 ;
        RECT 877.950 283.950 880.050 284.400 ;
        RECT 886.950 285.600 889.050 286.050 ;
        RECT 925.950 285.600 928.050 286.050 ;
        RECT 886.950 284.400 928.050 285.600 ;
        RECT 886.950 283.950 889.050 284.400 ;
        RECT 925.950 283.950 928.050 284.400 ;
        RECT 967.950 285.600 970.050 286.050 ;
        RECT 973.950 285.600 976.050 286.050 ;
        RECT 967.950 284.400 976.050 285.600 ;
        RECT 967.950 283.950 970.050 284.400 ;
        RECT 973.950 283.950 976.050 284.400 ;
        RECT 982.950 285.600 985.050 286.050 ;
        RECT 997.950 285.600 1000.050 286.050 ;
        RECT 982.950 284.400 1000.050 285.600 ;
        RECT 982.950 283.950 985.050 284.400 ;
        RECT 997.950 283.950 1000.050 284.400 ;
        RECT 103.950 282.600 106.050 283.050 ;
        RECT 115.950 282.600 118.050 283.050 ;
        RECT 103.950 281.400 118.050 282.600 ;
        RECT 103.950 280.950 106.050 281.400 ;
        RECT 115.950 280.950 118.050 281.400 ;
        RECT 175.950 281.400 180.600 283.050 ;
        RECT 199.950 282.600 202.050 283.050 ;
        RECT 223.950 282.600 226.050 283.050 ;
        RECT 199.950 281.400 226.050 282.600 ;
        RECT 175.950 280.950 180.000 281.400 ;
        RECT 199.950 280.950 202.050 281.400 ;
        RECT 223.950 280.950 226.050 281.400 ;
        RECT 247.950 282.600 250.050 283.050 ;
        RECT 256.950 282.600 259.050 283.050 ;
        RECT 247.950 281.400 259.050 282.600 ;
        RECT 247.950 280.950 250.050 281.400 ;
        RECT 256.950 280.950 259.050 281.400 ;
        RECT 445.950 282.600 448.050 283.050 ;
        RECT 505.950 282.600 508.050 283.050 ;
        RECT 445.950 281.400 508.050 282.600 ;
        RECT 445.950 280.950 448.050 281.400 ;
        RECT 505.950 280.950 508.050 281.400 ;
        RECT 517.950 282.600 520.050 283.050 ;
        RECT 586.950 282.600 589.050 283.050 ;
        RECT 631.950 282.600 634.050 283.050 ;
        RECT 685.950 282.600 688.050 283.050 ;
        RECT 517.950 281.400 570.600 282.600 ;
        RECT 517.950 280.950 520.050 281.400 ;
        RECT 37.950 279.600 40.050 280.050 ;
        RECT 88.950 279.600 91.050 280.050 ;
        RECT 37.950 278.400 91.050 279.600 ;
        RECT 37.950 277.950 40.050 278.400 ;
        RECT 88.950 277.950 91.050 278.400 ;
        RECT 97.950 279.600 100.050 280.050 ;
        RECT 136.950 279.600 139.050 280.050 ;
        RECT 97.950 278.400 139.050 279.600 ;
        RECT 97.950 277.950 100.050 278.400 ;
        RECT 136.950 277.950 139.050 278.400 ;
        RECT 181.950 279.600 184.050 280.050 ;
        RECT 211.950 279.600 214.050 280.050 ;
        RECT 181.950 278.400 214.050 279.600 ;
        RECT 181.950 277.950 184.050 278.400 ;
        RECT 211.950 277.950 214.050 278.400 ;
        RECT 325.950 279.600 328.050 280.050 ;
        RECT 355.950 279.600 358.050 280.050 ;
        RECT 361.950 279.600 364.050 280.050 ;
        RECT 325.950 278.400 364.050 279.600 ;
        RECT 325.950 277.950 328.050 278.400 ;
        RECT 355.950 277.950 358.050 278.400 ;
        RECT 361.950 277.950 364.050 278.400 ;
        RECT 367.950 279.600 370.050 280.050 ;
        RECT 382.950 279.600 385.050 280.050 ;
        RECT 367.950 278.400 385.050 279.600 ;
        RECT 367.950 277.950 370.050 278.400 ;
        RECT 382.950 277.950 385.050 278.400 ;
        RECT 517.950 279.600 520.050 279.900 ;
        RECT 565.950 279.600 568.050 280.050 ;
        RECT 517.950 278.400 568.050 279.600 ;
        RECT 569.400 279.600 570.600 281.400 ;
        RECT 586.950 281.400 634.050 282.600 ;
        RECT 586.950 280.950 589.050 281.400 ;
        RECT 631.950 280.950 634.050 281.400 ;
        RECT 635.400 281.400 688.050 282.600 ;
        RECT 635.400 279.600 636.600 281.400 ;
        RECT 685.950 280.950 688.050 281.400 ;
        RECT 703.950 282.600 706.050 283.050 ;
        RECT 718.950 282.600 721.050 283.050 ;
        RECT 703.950 281.400 721.050 282.600 ;
        RECT 703.950 280.950 706.050 281.400 ;
        RECT 718.950 280.950 721.050 281.400 ;
        RECT 730.950 282.600 733.050 283.050 ;
        RECT 742.950 282.600 745.050 283.050 ;
        RECT 790.950 282.600 793.050 283.050 ;
        RECT 730.950 281.400 745.050 282.600 ;
        RECT 730.950 280.950 733.050 281.400 ;
        RECT 742.950 280.950 745.050 281.400 ;
        RECT 746.400 281.400 793.050 282.600 ;
        RECT 569.400 278.400 636.600 279.600 ;
        RECT 691.950 279.600 694.050 280.050 ;
        RECT 746.400 279.600 747.600 281.400 ;
        RECT 790.950 280.950 793.050 281.400 ;
        RECT 937.950 282.600 940.050 283.050 ;
        RECT 943.950 282.600 946.050 283.050 ;
        RECT 937.950 281.400 946.050 282.600 ;
        RECT 937.950 280.950 940.050 281.400 ;
        RECT 943.950 280.950 946.050 281.400 ;
        RECT 979.950 282.600 982.050 283.050 ;
        RECT 1030.950 282.600 1033.050 283.050 ;
        RECT 979.950 281.400 1033.050 282.600 ;
        RECT 979.950 280.950 982.050 281.400 ;
        RECT 1030.950 280.950 1033.050 281.400 ;
        RECT 691.950 278.400 747.600 279.600 ;
        RECT 856.950 279.600 859.050 280.050 ;
        RECT 892.950 279.600 895.050 280.050 ;
        RECT 856.950 278.400 895.050 279.600 ;
        RECT 517.950 277.800 520.050 278.400 ;
        RECT 565.950 277.950 568.050 278.400 ;
        RECT 691.950 277.950 694.050 278.400 ;
        RECT 856.950 277.950 859.050 278.400 ;
        RECT 892.950 277.950 895.050 278.400 ;
        RECT 949.950 279.600 952.050 280.050 ;
        RECT 961.950 279.600 964.050 279.900 ;
        RECT 949.950 278.400 964.050 279.600 ;
        RECT 949.950 277.950 952.050 278.400 ;
        RECT 961.950 277.800 964.050 278.400 ;
        RECT 151.950 276.600 154.050 277.050 ;
        RECT 229.950 276.600 232.050 277.050 ;
        RECT 151.950 275.400 232.050 276.600 ;
        RECT 151.950 274.950 154.050 275.400 ;
        RECT 229.950 274.950 232.050 275.400 ;
        RECT 292.950 276.600 295.050 277.050 ;
        RECT 307.950 276.600 310.050 277.050 ;
        RECT 292.950 275.400 310.050 276.600 ;
        RECT 292.950 274.950 295.050 275.400 ;
        RECT 307.950 274.950 310.050 275.400 ;
        RECT 331.950 276.600 334.050 277.050 ;
        RECT 343.950 276.600 346.050 277.050 ;
        RECT 331.950 275.400 346.050 276.600 ;
        RECT 331.950 274.950 334.050 275.400 ;
        RECT 343.950 274.950 346.050 275.400 ;
        RECT 421.950 276.600 424.050 277.050 ;
        RECT 502.950 276.600 505.050 277.050 ;
        RECT 514.950 276.600 517.050 277.050 ;
        RECT 571.950 276.600 574.050 277.050 ;
        RECT 577.950 276.600 580.050 277.050 ;
        RECT 685.950 276.600 688.050 277.050 ;
        RECT 778.950 276.600 781.050 277.050 ;
        RECT 814.950 276.600 817.050 277.050 ;
        RECT 421.950 275.400 817.050 276.600 ;
        RECT 421.950 274.950 424.050 275.400 ;
        RECT 502.950 274.950 505.050 275.400 ;
        RECT 514.950 274.950 517.050 275.400 ;
        RECT 571.950 274.950 574.050 275.400 ;
        RECT 577.950 274.950 580.050 275.400 ;
        RECT 685.950 274.950 688.050 275.400 ;
        RECT 778.950 274.950 781.050 275.400 ;
        RECT 814.950 274.950 817.050 275.400 ;
        RECT 949.950 276.600 952.050 276.900 ;
        RECT 958.950 276.600 961.050 277.050 ;
        RECT 949.950 275.400 961.050 276.600 ;
        RECT 949.950 274.800 952.050 275.400 ;
        RECT 958.950 274.950 961.050 275.400 ;
        RECT 970.950 276.600 973.050 277.050 ;
        RECT 994.950 276.600 997.050 277.050 ;
        RECT 970.950 275.400 997.050 276.600 ;
        RECT 970.950 274.950 973.050 275.400 ;
        RECT 994.950 274.950 997.050 275.400 ;
        RECT 127.950 273.600 130.050 274.050 ;
        RECT 304.950 273.600 307.050 274.050 ;
        RECT 127.950 272.400 307.050 273.600 ;
        RECT 127.950 271.950 130.050 272.400 ;
        RECT 304.950 271.950 307.050 272.400 ;
        RECT 496.950 273.600 499.050 274.050 ;
        RECT 508.950 273.600 511.050 274.050 ;
        RECT 496.950 272.400 511.050 273.600 ;
        RECT 496.950 271.950 499.050 272.400 ;
        RECT 508.950 271.950 511.050 272.400 ;
        RECT 592.950 273.600 595.050 274.050 ;
        RECT 604.950 273.600 607.050 274.050 ;
        RECT 592.950 272.400 607.050 273.600 ;
        RECT 592.950 271.950 595.050 272.400 ;
        RECT 604.950 271.950 607.050 272.400 ;
        RECT 643.950 273.600 646.050 274.050 ;
        RECT 655.950 273.600 658.050 274.050 ;
        RECT 643.950 272.400 658.050 273.600 ;
        RECT 643.950 271.950 646.050 272.400 ;
        RECT 655.950 271.950 658.050 272.400 ;
        RECT 691.950 273.600 694.050 274.050 ;
        RECT 697.950 273.600 700.050 274.050 ;
        RECT 691.950 272.400 700.050 273.600 ;
        RECT 691.950 271.950 694.050 272.400 ;
        RECT 697.950 271.950 700.050 272.400 ;
        RECT 712.950 271.950 715.050 274.050 ;
        RECT 724.950 273.600 727.050 274.050 ;
        RECT 745.950 273.600 748.050 274.050 ;
        RECT 724.950 272.400 748.050 273.600 ;
        RECT 724.950 271.950 727.050 272.400 ;
        RECT 745.950 271.950 748.050 272.400 ;
        RECT 757.950 273.600 760.050 274.050 ;
        RECT 775.950 273.600 778.050 274.050 ;
        RECT 757.950 272.400 778.050 273.600 ;
        RECT 757.950 271.950 760.050 272.400 ;
        RECT 775.950 271.950 778.050 272.400 ;
        RECT 925.950 273.600 928.050 274.050 ;
        RECT 964.950 273.600 967.050 274.050 ;
        RECT 925.950 272.400 967.050 273.600 ;
        RECT 925.950 271.950 928.050 272.400 ;
        RECT 964.950 271.950 967.050 272.400 ;
        RECT 973.950 273.600 976.050 274.050 ;
        RECT 982.950 273.600 985.050 274.050 ;
        RECT 973.950 272.400 985.050 273.600 ;
        RECT 973.950 271.950 976.050 272.400 ;
        RECT 982.950 271.950 985.050 272.400 ;
        RECT 46.950 270.600 49.050 271.050 ;
        RECT 58.950 270.600 61.050 271.050 ;
        RECT 46.950 269.400 61.050 270.600 ;
        RECT 46.950 268.950 49.050 269.400 ;
        RECT 58.950 268.950 61.050 269.400 ;
        RECT 208.950 270.600 211.050 271.050 ;
        RECT 217.950 270.600 220.050 271.050 ;
        RECT 226.950 270.600 229.050 271.050 ;
        RECT 208.950 269.400 229.050 270.600 ;
        RECT 208.950 268.950 211.050 269.400 ;
        RECT 217.950 268.950 220.050 269.400 ;
        RECT 226.950 268.950 229.050 269.400 ;
        RECT 547.950 270.600 550.050 271.050 ;
        RECT 619.950 270.600 622.050 271.050 ;
        RECT 547.950 269.400 622.050 270.600 ;
        RECT 547.950 268.950 550.050 269.400 ;
        RECT 619.950 268.950 622.050 269.400 ;
        RECT 13.950 267.600 16.050 268.050 ;
        RECT 73.950 267.600 76.050 268.050 ;
        RECT 13.950 266.400 76.050 267.600 ;
        RECT 13.950 265.950 16.050 266.400 ;
        RECT 73.950 265.950 76.050 266.400 ;
        RECT 289.950 267.600 292.050 268.050 ;
        RECT 304.950 267.600 307.050 268.050 ;
        RECT 289.950 266.400 307.050 267.600 ;
        RECT 289.950 265.950 292.050 266.400 ;
        RECT 304.950 265.950 307.050 266.400 ;
        RECT 409.950 267.600 412.050 268.050 ;
        RECT 622.950 267.600 625.050 268.050 ;
        RECT 409.950 266.400 625.050 267.600 ;
        RECT 409.950 265.950 412.050 266.400 ;
        RECT 622.950 265.950 625.050 266.400 ;
        RECT 655.950 267.600 658.050 268.050 ;
        RECT 670.950 267.600 673.050 268.050 ;
        RECT 655.950 266.400 673.050 267.600 ;
        RECT 655.950 265.950 658.050 266.400 ;
        RECT 670.950 265.950 673.050 266.400 ;
        RECT 676.950 267.600 679.050 268.050 ;
        RECT 682.950 267.600 685.050 268.050 ;
        RECT 676.950 266.400 685.050 267.600 ;
        RECT 676.950 265.950 679.050 266.400 ;
        RECT 682.950 265.950 685.050 266.400 ;
        RECT 115.950 264.600 118.050 265.050 ;
        RECT 148.950 264.600 151.050 265.050 ;
        RECT 115.950 263.400 151.050 264.600 ;
        RECT 115.950 262.950 118.050 263.400 ;
        RECT 148.950 262.950 151.050 263.400 ;
        RECT 190.950 264.600 193.050 265.050 ;
        RECT 238.950 264.600 241.050 265.050 ;
        RECT 190.950 263.400 241.050 264.600 ;
        RECT 190.950 262.950 193.050 263.400 ;
        RECT 238.950 262.950 241.050 263.400 ;
        RECT 16.950 261.600 19.050 262.200 ;
        RECT 52.950 261.750 55.050 262.200 ;
        RECT 61.950 261.750 64.050 262.200 ;
        RECT 52.950 261.600 64.050 261.750 ;
        RECT 16.950 260.550 64.050 261.600 ;
        RECT 16.950 260.400 55.050 260.550 ;
        RECT 16.950 260.100 19.050 260.400 ;
        RECT 52.950 260.100 55.050 260.400 ;
        RECT 61.950 260.100 64.050 260.550 ;
        RECT 97.950 261.750 100.050 262.200 ;
        RECT 109.950 261.750 112.050 262.200 ;
        RECT 97.950 260.550 112.050 261.750 ;
        RECT 97.950 260.100 100.050 260.550 ;
        RECT 109.950 260.100 112.050 260.550 ;
        RECT 118.950 261.750 121.050 262.200 ;
        RECT 127.950 261.750 130.050 262.200 ;
        RECT 118.950 260.550 130.050 261.750 ;
        RECT 118.950 260.100 121.050 260.550 ;
        RECT 127.950 260.100 130.050 260.550 ;
        RECT 154.950 261.750 157.050 262.200 ;
        RECT 163.950 261.750 166.050 262.200 ;
        RECT 154.950 260.550 166.050 261.750 ;
        RECT 154.950 260.100 157.050 260.550 ;
        RECT 163.950 260.100 166.050 260.550 ;
        RECT 181.950 261.750 184.050 262.200 ;
        RECT 187.950 261.750 190.050 262.200 ;
        RECT 181.950 260.550 190.050 261.750 ;
        RECT 181.950 260.100 184.050 260.550 ;
        RECT 187.950 260.100 190.050 260.550 ;
        RECT 193.950 261.600 196.050 262.050 ;
        RECT 202.950 261.600 205.050 262.200 ;
        RECT 193.950 260.400 205.050 261.600 ;
        RECT 193.950 259.950 196.050 260.400 ;
        RECT 202.950 260.100 205.050 260.400 ;
        RECT 211.950 261.600 214.050 262.050 ;
        RECT 232.950 261.600 235.050 262.050 ;
        RECT 211.950 260.400 235.050 261.600 ;
        RECT 211.950 259.950 214.050 260.400 ;
        RECT 232.950 259.950 235.050 260.400 ;
        RECT 250.950 261.600 253.050 262.200 ;
        RECT 268.950 261.600 271.050 262.200 ;
        RECT 250.950 260.400 271.050 261.600 ;
        RECT 250.950 260.100 253.050 260.400 ;
        RECT 268.950 260.100 271.050 260.400 ;
        RECT 283.950 261.750 286.050 262.200 ;
        RECT 295.950 261.750 298.050 262.200 ;
        RECT 283.950 260.550 298.050 261.750 ;
        RECT 283.950 260.100 286.050 260.550 ;
        RECT 295.950 260.100 298.050 260.550 ;
        RECT 301.950 261.600 304.050 262.050 ;
        RECT 316.950 261.600 319.050 262.200 ;
        RECT 301.950 260.400 319.050 261.600 ;
        RECT 301.950 259.950 304.050 260.400 ;
        RECT 316.950 260.100 319.050 260.400 ;
        RECT 334.950 261.600 337.050 262.050 ;
        RECT 403.950 261.600 406.050 262.050 ;
        RECT 409.950 261.600 412.050 262.050 ;
        RECT 589.950 261.600 592.050 262.200 ;
        RECT 334.950 260.400 412.050 261.600 ;
        RECT 334.950 259.950 337.050 260.400 ;
        RECT 403.950 259.950 406.050 260.400 ;
        RECT 409.950 259.950 412.050 260.400 ;
        RECT 581.400 260.400 592.050 261.600 ;
        RECT 325.950 257.100 328.050 259.200 ;
        RECT 361.950 258.450 364.050 258.900 ;
        RECT 382.950 258.450 385.050 258.900 ;
        RECT 361.950 257.250 385.050 258.450 ;
        RECT 326.400 256.050 327.600 257.100 ;
        RECT 361.950 256.800 364.050 257.250 ;
        RECT 382.950 256.800 385.050 257.250 ;
        RECT 394.950 258.750 397.050 259.200 ;
        RECT 400.950 258.750 403.050 259.200 ;
        RECT 394.950 257.550 403.050 258.750 ;
        RECT 394.950 257.100 397.050 257.550 ;
        RECT 400.950 257.100 403.050 257.550 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 487.950 258.450 490.050 258.900 ;
        RECT 517.950 258.450 520.050 258.900 ;
        RECT 581.400 258.600 582.600 260.400 ;
        RECT 589.950 260.100 592.050 260.400 ;
        RECT 598.950 261.600 601.050 262.050 ;
        RECT 613.950 261.600 616.050 262.200 ;
        RECT 598.950 260.400 616.050 261.600 ;
        RECT 598.950 259.950 601.050 260.400 ;
        RECT 613.950 260.100 616.050 260.400 ;
        RECT 628.950 261.600 631.050 262.050 ;
        RECT 637.950 261.600 640.050 262.200 ;
        RECT 628.950 260.400 640.050 261.600 ;
        RECT 628.950 259.950 631.050 260.400 ;
        RECT 637.950 260.100 640.050 260.400 ;
        RECT 643.950 261.600 646.050 262.200 ;
        RECT 661.950 261.600 664.050 262.200 ;
        RECT 643.950 260.400 664.050 261.600 ;
        RECT 643.950 260.100 646.050 260.400 ;
        RECT 661.950 260.100 664.050 260.400 ;
        RECT 667.950 261.600 670.050 262.200 ;
        RECT 667.950 260.400 675.600 261.600 ;
        RECT 667.950 260.100 670.050 260.400 ;
        RECT 487.950 257.250 520.050 258.450 ;
        RECT 31.950 255.450 34.050 255.900 ;
        RECT 40.950 255.450 43.050 255.900 ;
        RECT 31.950 254.250 43.050 255.450 ;
        RECT 31.950 253.800 34.050 254.250 ;
        RECT 40.950 253.800 43.050 254.250 ;
        RECT 64.950 255.450 67.050 255.900 ;
        RECT 70.950 255.450 73.050 255.900 ;
        RECT 64.950 254.250 73.050 255.450 ;
        RECT 64.950 253.800 67.050 254.250 ;
        RECT 70.950 253.800 73.050 254.250 ;
        RECT 106.950 255.600 109.050 256.050 ;
        RECT 112.950 255.600 115.050 256.050 ;
        RECT 106.950 254.400 115.050 255.600 ;
        RECT 106.950 253.950 109.050 254.400 ;
        RECT 112.950 253.950 115.050 254.400 ;
        RECT 142.950 255.600 145.050 256.050 ;
        RECT 151.950 255.600 154.050 255.900 ;
        RECT 142.950 254.400 154.050 255.600 ;
        RECT 142.950 253.950 145.050 254.400 ;
        RECT 151.950 253.800 154.050 254.400 ;
        RECT 178.950 255.450 181.050 255.900 ;
        RECT 193.950 255.450 196.050 255.900 ;
        RECT 178.950 254.250 196.050 255.450 ;
        RECT 178.950 253.800 181.050 254.250 ;
        RECT 193.950 253.800 196.050 254.250 ;
        RECT 229.950 255.450 232.050 255.900 ;
        RECT 253.950 255.450 256.050 255.900 ;
        RECT 229.950 254.250 256.050 255.450 ;
        RECT 229.950 253.800 232.050 254.250 ;
        RECT 253.950 253.800 256.050 254.250 ;
        RECT 271.950 255.600 274.050 255.900 ;
        RECT 286.950 255.600 289.050 256.050 ;
        RECT 271.950 254.400 289.050 255.600 ;
        RECT 271.950 253.800 274.050 254.400 ;
        RECT 286.950 253.950 289.050 254.400 ;
        RECT 307.950 255.450 310.050 255.900 ;
        RECT 313.950 255.450 316.050 255.900 ;
        RECT 307.950 254.250 316.050 255.450 ;
        RECT 307.950 253.800 310.050 254.250 ;
        RECT 313.950 253.800 316.050 254.250 ;
        RECT 322.950 254.400 327.600 256.050 ;
        RECT 322.950 253.950 327.000 254.400 ;
        RECT 175.950 252.600 178.050 253.050 ;
        RECT 199.950 252.600 202.050 253.050 ;
        RECT 175.950 251.400 202.050 252.600 ;
        RECT 175.950 250.950 178.050 251.400 ;
        RECT 199.950 250.950 202.050 251.400 ;
        RECT 280.950 252.600 283.050 253.050 ;
        RECT 292.950 252.600 295.050 253.050 ;
        RECT 280.950 251.400 295.050 252.600 ;
        RECT 280.950 250.950 283.050 251.400 ;
        RECT 292.950 250.950 295.050 251.400 ;
        RECT 382.950 252.600 385.050 253.050 ;
        RECT 409.950 252.600 412.050 253.050 ;
        RECT 382.950 251.400 412.050 252.600 ;
        RECT 382.950 250.950 385.050 251.400 ;
        RECT 409.950 250.950 412.050 251.400 ;
        RECT 454.950 252.600 457.050 252.900 ;
        RECT 461.400 252.600 462.600 256.950 ;
        RECT 487.950 256.800 490.050 257.250 ;
        RECT 517.950 256.800 520.050 257.250 ;
        RECT 548.400 257.400 582.600 258.600 ;
        RECT 526.950 255.600 529.050 256.050 ;
        RECT 544.950 255.600 547.050 255.900 ;
        RECT 548.400 255.600 549.600 257.400 ;
        RECT 674.400 256.050 675.600 260.400 ;
        RECT 713.400 258.900 714.600 271.950 ;
        RECT 772.950 270.600 775.050 271.050 ;
        RECT 799.950 270.600 802.050 271.050 ;
        RECT 772.950 269.400 802.050 270.600 ;
        RECT 772.950 268.950 775.050 269.400 ;
        RECT 799.950 268.950 802.050 269.400 ;
        RECT 805.950 270.600 808.050 271.050 ;
        RECT 820.950 270.600 823.050 271.050 ;
        RECT 805.950 269.400 823.050 270.600 ;
        RECT 805.950 268.950 808.050 269.400 ;
        RECT 820.950 268.950 823.050 269.400 ;
        RECT 934.950 270.600 937.050 271.050 ;
        RECT 970.950 270.600 973.050 271.050 ;
        RECT 934.950 269.400 973.050 270.600 ;
        RECT 934.950 268.950 937.050 269.400 ;
        RECT 970.950 268.950 973.050 269.400 ;
        RECT 976.950 270.600 979.050 271.050 ;
        RECT 988.950 270.600 991.050 271.050 ;
        RECT 976.950 269.400 991.050 270.600 ;
        RECT 976.950 268.950 979.050 269.400 ;
        RECT 988.950 268.950 991.050 269.400 ;
        RECT 811.950 267.600 814.050 268.050 ;
        RECT 817.950 267.600 820.050 268.050 ;
        RECT 811.950 266.400 820.050 267.600 ;
        RECT 811.950 265.950 814.050 266.400 ;
        RECT 817.950 265.950 820.050 266.400 ;
        RECT 892.950 267.600 895.050 268.050 ;
        RECT 907.950 267.600 910.050 268.050 ;
        RECT 892.950 266.400 910.050 267.600 ;
        RECT 971.400 267.600 972.600 268.950 ;
        RECT 997.950 267.600 1000.050 268.050 ;
        RECT 971.400 266.400 1000.050 267.600 ;
        RECT 892.950 265.950 895.050 266.400 ;
        RECT 907.950 265.950 910.050 266.400 ;
        RECT 997.950 265.950 1000.050 266.400 ;
        RECT 1012.950 265.050 1015.050 265.200 ;
        RECT 919.950 264.600 922.050 265.050 ;
        RECT 848.400 263.400 922.050 264.600 ;
        RECT 772.950 261.600 775.050 262.200 ;
        RECT 784.950 261.600 787.050 262.050 ;
        RECT 790.950 261.600 793.050 262.200 ;
        RECT 772.950 260.400 793.050 261.600 ;
        RECT 772.950 260.100 775.050 260.400 ;
        RECT 784.950 259.950 787.050 260.400 ;
        RECT 790.950 260.100 793.050 260.400 ;
        RECT 811.950 260.100 814.050 262.200 ;
        RECT 817.950 261.600 820.050 262.200 ;
        RECT 817.950 260.400 828.600 261.600 ;
        RECT 817.950 260.100 820.050 260.400 ;
        RECT 712.950 256.800 715.050 258.900 ;
        RECT 812.400 258.600 813.600 260.100 ;
        RECT 809.400 258.000 813.600 258.600 ;
        RECT 808.950 257.400 813.600 258.000 ;
        RECT 526.950 254.400 549.600 255.600 ;
        RECT 550.950 255.450 553.050 255.900 ;
        RECT 556.950 255.450 559.050 255.900 ;
        RECT 526.950 253.950 529.050 254.400 ;
        RECT 544.950 253.800 547.050 254.400 ;
        RECT 550.950 254.250 559.050 255.450 ;
        RECT 550.950 253.800 553.050 254.250 ;
        RECT 556.950 253.800 559.050 254.250 ;
        RECT 640.950 255.600 643.050 255.900 ;
        RECT 655.950 255.600 658.050 255.900 ;
        RECT 640.950 255.450 658.050 255.600 ;
        RECT 664.950 255.450 667.050 255.900 ;
        RECT 640.950 254.400 667.050 255.450 ;
        RECT 640.950 253.800 643.050 254.400 ;
        RECT 655.950 254.250 667.050 254.400 ;
        RECT 655.950 253.800 658.050 254.250 ;
        RECT 664.950 253.800 667.050 254.250 ;
        RECT 673.950 253.950 676.050 256.050 ;
        RECT 781.950 255.600 784.050 256.050 ;
        RECT 793.950 255.600 796.050 255.900 ;
        RECT 781.950 254.400 796.050 255.600 ;
        RECT 781.950 253.950 784.050 254.400 ;
        RECT 793.950 253.800 796.050 254.400 ;
        RECT 808.950 253.950 811.050 257.400 ;
        RECT 827.400 253.050 828.600 260.400 ;
        RECT 848.400 258.900 849.600 263.400 ;
        RECT 919.950 262.950 922.050 263.400 ;
        RECT 946.950 264.600 949.050 265.050 ;
        RECT 955.950 264.600 958.050 265.050 ;
        RECT 946.950 263.400 958.050 264.600 ;
        RECT 946.950 262.950 949.050 263.400 ;
        RECT 955.950 262.950 958.050 263.400 ;
        RECT 964.950 264.600 967.050 265.050 ;
        RECT 979.950 264.600 982.050 265.050 ;
        RECT 1011.000 264.600 1015.050 265.050 ;
        RECT 964.950 263.400 982.050 264.600 ;
        RECT 964.950 262.950 967.050 263.400 ;
        RECT 979.950 262.950 982.050 263.400 ;
        RECT 1010.400 263.100 1015.050 264.600 ;
        RECT 1021.950 264.600 1024.050 265.050 ;
        RECT 1033.950 264.600 1036.050 265.050 ;
        RECT 1021.950 263.400 1036.050 264.600 ;
        RECT 1010.400 262.950 1014.000 263.100 ;
        RECT 1021.950 262.950 1024.050 263.400 ;
        RECT 1033.950 262.950 1036.050 263.400 ;
        RECT 910.950 261.750 913.050 262.200 ;
        RECT 922.950 261.750 925.050 262.200 ;
        RECT 910.950 260.550 925.050 261.750 ;
        RECT 961.950 261.600 964.050 262.200 ;
        RECT 910.950 260.100 913.050 260.550 ;
        RECT 922.950 260.100 925.050 260.550 ;
        RECT 953.400 260.400 964.050 261.600 ;
        RECT 847.950 256.800 850.050 258.900 ;
        RECT 871.950 258.750 874.050 259.200 ;
        RECT 883.950 258.750 886.050 259.200 ;
        RECT 871.950 258.600 886.050 258.750 ;
        RECT 898.950 258.600 901.050 259.050 ;
        RECT 871.950 257.550 901.050 258.600 ;
        RECT 871.950 257.100 874.050 257.550 ;
        RECT 883.950 257.400 901.050 257.550 ;
        RECT 883.950 257.100 886.050 257.400 ;
        RECT 898.950 256.950 901.050 257.400 ;
        RECT 953.400 256.050 954.600 260.400 ;
        RECT 961.950 260.100 964.050 260.400 ;
        RECT 1000.950 261.600 1003.050 262.050 ;
        RECT 1006.950 261.600 1009.050 262.200 ;
        RECT 1000.950 260.400 1009.050 261.600 ;
        RECT 1000.950 259.950 1003.050 260.400 ;
        RECT 1006.950 260.100 1009.050 260.400 ;
        RECT 907.950 255.450 910.050 255.900 ;
        RECT 946.950 255.450 949.050 255.900 ;
        RECT 907.950 254.250 949.050 255.450 ;
        RECT 907.950 253.800 910.050 254.250 ;
        RECT 946.950 253.800 949.050 254.250 ;
        RECT 952.950 253.950 955.050 256.050 ;
        RECT 1010.400 255.900 1011.600 262.950 ;
        RECT 1012.950 261.600 1015.050 262.050 ;
        RECT 1024.950 261.600 1027.050 262.050 ;
        RECT 1012.950 260.400 1027.050 261.600 ;
        RECT 1012.950 259.950 1015.050 260.400 ;
        RECT 1024.950 259.950 1027.050 260.400 ;
        RECT 1039.800 260.100 1041.900 262.200 ;
        RECT 1042.950 261.600 1047.000 262.050 ;
        RECT 1040.400 256.050 1041.600 260.100 ;
        RECT 1042.950 259.950 1047.600 261.600 ;
        RECT 964.950 255.450 967.050 255.900 ;
        RECT 970.950 255.450 973.050 255.900 ;
        RECT 964.950 254.250 973.050 255.450 ;
        RECT 964.950 253.800 967.050 254.250 ;
        RECT 970.950 253.800 973.050 254.250 ;
        RECT 997.950 255.450 1000.050 255.900 ;
        RECT 1003.950 255.450 1006.050 255.900 ;
        RECT 997.950 254.250 1006.050 255.450 ;
        RECT 997.950 253.800 1000.050 254.250 ;
        RECT 1003.950 253.800 1006.050 254.250 ;
        RECT 1009.950 253.800 1012.050 255.900 ;
        RECT 1018.950 255.450 1021.050 255.900 ;
        RECT 1036.950 255.450 1039.050 255.900 ;
        RECT 1018.950 254.250 1039.050 255.450 ;
        RECT 1040.400 254.400 1045.050 256.050 ;
        RECT 1018.950 253.800 1021.050 254.250 ;
        RECT 1036.950 253.800 1039.050 254.250 ;
        RECT 1041.000 253.950 1045.050 254.400 ;
        RECT 463.950 252.600 466.050 252.900 ;
        RECT 454.950 252.450 466.050 252.600 ;
        RECT 487.950 252.450 490.050 252.900 ;
        RECT 454.950 251.400 490.050 252.450 ;
        RECT 454.950 250.800 457.050 251.400 ;
        RECT 463.950 251.250 490.050 251.400 ;
        RECT 463.950 250.800 466.050 251.250 ;
        RECT 487.950 250.800 490.050 251.250 ;
        RECT 826.950 250.950 829.050 253.050 ;
        RECT 847.950 252.600 850.050 253.050 ;
        RECT 877.950 252.600 880.050 253.050 ;
        RECT 913.950 252.600 916.050 253.050 ;
        RECT 847.950 251.400 916.050 252.600 ;
        RECT 847.950 250.950 850.050 251.400 ;
        RECT 877.950 250.950 880.050 251.400 ;
        RECT 913.950 250.950 916.050 251.400 ;
        RECT 1024.950 252.600 1027.050 253.050 ;
        RECT 1030.950 252.600 1033.050 253.050 ;
        RECT 1024.950 251.400 1033.050 252.600 ;
        RECT 1024.950 250.950 1027.050 251.400 ;
        RECT 1030.950 250.950 1033.050 251.400 ;
        RECT 1039.950 252.600 1042.050 253.050 ;
        RECT 1046.400 252.600 1047.600 259.950 ;
        RECT 1039.950 251.400 1047.600 252.600 ;
        RECT 1039.950 250.950 1042.050 251.400 ;
        RECT 247.950 249.600 250.050 250.050 ;
        RECT 262.950 249.600 265.050 250.050 ;
        RECT 247.950 248.400 265.050 249.600 ;
        RECT 247.950 247.950 250.050 248.400 ;
        RECT 262.950 247.950 265.050 248.400 ;
        RECT 322.950 249.600 325.050 250.050 ;
        RECT 334.950 249.600 337.050 250.050 ;
        RECT 322.950 248.400 337.050 249.600 ;
        RECT 322.950 247.950 325.050 248.400 ;
        RECT 334.950 247.950 337.050 248.400 ;
        RECT 592.950 249.600 595.050 250.050 ;
        RECT 610.950 249.600 613.050 250.050 ;
        RECT 727.950 249.600 730.050 250.050 ;
        RECT 592.950 248.400 730.050 249.600 ;
        RECT 592.950 247.950 595.050 248.400 ;
        RECT 610.950 247.950 613.050 248.400 ;
        RECT 727.950 247.950 730.050 248.400 ;
        RECT 736.950 249.600 739.050 250.050 ;
        RECT 805.950 249.600 808.050 250.050 ;
        RECT 823.950 249.600 826.050 250.050 ;
        RECT 736.950 248.400 826.050 249.600 ;
        RECT 736.950 247.950 739.050 248.400 ;
        RECT 805.950 247.950 808.050 248.400 ;
        RECT 823.950 247.950 826.050 248.400 ;
        RECT 898.950 249.600 901.050 250.050 ;
        RECT 931.950 249.600 934.050 250.050 ;
        RECT 898.950 248.400 934.050 249.600 ;
        RECT 898.950 247.950 901.050 248.400 ;
        RECT 931.950 247.950 934.050 248.400 ;
        RECT 43.950 246.600 46.050 247.050 ;
        RECT 52.950 246.600 55.050 247.050 ;
        RECT 43.950 245.400 55.050 246.600 ;
        RECT 43.950 244.950 46.050 245.400 ;
        RECT 52.950 244.950 55.050 245.400 ;
        RECT 127.950 246.600 130.050 247.050 ;
        RECT 133.950 246.600 136.050 247.050 ;
        RECT 127.950 245.400 136.050 246.600 ;
        RECT 127.950 244.950 130.050 245.400 ;
        RECT 133.950 244.950 136.050 245.400 ;
        RECT 187.950 246.600 190.050 247.050 ;
        RECT 223.950 246.600 226.050 247.050 ;
        RECT 301.950 246.600 304.050 247.050 ;
        RECT 310.950 246.600 313.050 247.050 ;
        RECT 187.950 245.400 313.050 246.600 ;
        RECT 187.950 244.950 190.050 245.400 ;
        RECT 223.950 244.950 226.050 245.400 ;
        RECT 301.950 244.950 304.050 245.400 ;
        RECT 310.950 244.950 313.050 245.400 ;
        RECT 511.950 246.600 514.050 247.050 ;
        RECT 550.950 246.600 553.050 247.050 ;
        RECT 511.950 245.400 553.050 246.600 ;
        RECT 511.950 244.950 514.050 245.400 ;
        RECT 550.950 244.950 553.050 245.400 ;
        RECT 979.950 246.600 982.050 247.050 ;
        RECT 991.950 246.600 994.050 247.050 ;
        RECT 979.950 245.400 994.050 246.600 ;
        RECT 979.950 244.950 982.050 245.400 ;
        RECT 991.950 244.950 994.050 245.400 ;
        RECT 100.950 243.600 103.050 244.050 ;
        RECT 130.950 243.600 133.050 244.050 ;
        RECT 100.950 242.400 133.050 243.600 ;
        RECT 100.950 241.950 103.050 242.400 ;
        RECT 130.950 241.950 133.050 242.400 ;
        RECT 319.950 243.600 322.050 244.050 ;
        RECT 400.950 243.600 403.050 244.050 ;
        RECT 319.950 242.400 403.050 243.600 ;
        RECT 319.950 241.950 322.050 242.400 ;
        RECT 400.950 241.950 403.050 242.400 ;
        RECT 517.950 243.600 520.050 244.050 ;
        RECT 598.950 243.600 601.050 244.050 ;
        RECT 517.950 242.400 601.050 243.600 ;
        RECT 517.950 241.950 520.050 242.400 ;
        RECT 598.950 241.950 601.050 242.400 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 808.950 243.600 811.050 244.050 ;
        RECT 649.950 242.400 811.050 243.600 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 808.950 241.950 811.050 242.400 ;
        RECT 40.950 240.600 43.050 241.050 ;
        RECT 109.950 240.600 112.050 241.050 ;
        RECT 256.950 240.600 259.050 241.050 ;
        RECT 484.950 240.600 487.050 241.050 ;
        RECT 40.950 239.400 123.600 240.600 ;
        RECT 40.950 238.950 43.050 239.400 ;
        RECT 109.950 238.950 112.050 239.400 ;
        RECT 122.400 237.600 123.600 239.400 ;
        RECT 256.950 239.400 487.050 240.600 ;
        RECT 256.950 238.950 259.050 239.400 ;
        RECT 484.950 238.950 487.050 239.400 ;
        RECT 814.950 240.600 817.050 241.050 ;
        RECT 847.950 240.600 850.050 241.050 ;
        RECT 814.950 239.400 850.050 240.600 ;
        RECT 814.950 238.950 817.050 239.400 ;
        RECT 847.950 238.950 850.050 239.400 ;
        RECT 1003.950 240.600 1006.050 241.050 ;
        RECT 1021.950 240.600 1024.050 241.050 ;
        RECT 1003.950 239.400 1024.050 240.600 ;
        RECT 1003.950 238.950 1006.050 239.400 ;
        RECT 1021.950 238.950 1024.050 239.400 ;
        RECT 133.950 237.600 136.050 238.050 ;
        RECT 122.400 236.400 136.050 237.600 ;
        RECT 133.950 235.950 136.050 236.400 ;
        RECT 196.950 237.600 199.050 238.050 ;
        RECT 232.950 237.600 235.050 238.050 ;
        RECT 196.950 236.400 235.050 237.600 ;
        RECT 196.950 235.950 199.050 236.400 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 340.950 237.600 343.050 238.050 ;
        RECT 352.950 237.600 355.050 238.050 ;
        RECT 340.950 236.400 355.050 237.600 ;
        RECT 340.950 235.950 343.050 236.400 ;
        RECT 352.950 235.950 355.050 236.400 ;
        RECT 430.950 237.600 433.050 238.050 ;
        RECT 439.950 237.600 442.050 238.050 ;
        RECT 430.950 236.400 442.050 237.600 ;
        RECT 430.950 235.950 433.050 236.400 ;
        RECT 439.950 235.950 442.050 236.400 ;
        RECT 616.950 237.600 619.050 238.050 ;
        RECT 724.950 237.600 727.050 238.050 ;
        RECT 616.950 236.400 727.050 237.600 ;
        RECT 616.950 235.950 619.050 236.400 ;
        RECT 724.950 235.950 727.050 236.400 ;
        RECT 799.950 237.600 802.050 238.050 ;
        RECT 808.950 237.600 811.050 238.050 ;
        RECT 799.950 236.400 811.050 237.600 ;
        RECT 799.950 235.950 802.050 236.400 ;
        RECT 808.950 235.950 811.050 236.400 ;
        RECT 892.950 237.600 895.050 238.050 ;
        RECT 985.950 237.600 988.050 238.050 ;
        RECT 892.950 236.400 988.050 237.600 ;
        RECT 892.950 235.950 895.050 236.400 ;
        RECT 985.950 235.950 988.050 236.400 ;
        RECT 997.950 237.600 1000.050 238.050 ;
        RECT 1033.950 237.600 1036.050 238.050 ;
        RECT 997.950 236.400 1036.050 237.600 ;
        RECT 997.950 235.950 1000.050 236.400 ;
        RECT 1033.950 235.950 1036.050 236.400 ;
        RECT 28.950 234.600 31.050 235.050 ;
        RECT 64.950 234.600 67.050 235.050 ;
        RECT 28.950 233.400 67.050 234.600 ;
        RECT 28.950 232.950 31.050 233.400 ;
        RECT 64.950 232.950 67.050 233.400 ;
        RECT 118.950 234.600 121.050 235.050 ;
        RECT 160.950 234.600 163.050 235.050 ;
        RECT 187.950 234.600 190.050 235.050 ;
        RECT 256.950 234.600 259.050 235.050 ;
        RECT 118.950 233.400 150.600 234.600 ;
        RECT 118.950 232.950 121.050 233.400 ;
        RECT 149.400 232.050 150.600 233.400 ;
        RECT 160.950 233.400 259.050 234.600 ;
        RECT 160.950 232.950 163.050 233.400 ;
        RECT 187.950 232.950 190.050 233.400 ;
        RECT 256.950 232.950 259.050 233.400 ;
        RECT 571.950 234.600 574.050 235.050 ;
        RECT 580.950 234.600 583.050 235.050 ;
        RECT 598.950 234.600 601.050 235.050 ;
        RECT 571.950 233.400 601.050 234.600 ;
        RECT 571.950 232.950 574.050 233.400 ;
        RECT 580.950 232.950 583.050 233.400 ;
        RECT 598.950 232.950 601.050 233.400 ;
        RECT 922.950 234.600 925.050 235.050 ;
        RECT 1006.950 234.600 1009.050 235.050 ;
        RECT 922.950 233.400 1009.050 234.600 ;
        RECT 922.950 232.950 925.050 233.400 ;
        RECT 1006.950 232.950 1009.050 233.400 ;
        RECT 76.950 231.600 79.050 232.050 ;
        RECT 115.950 231.600 118.050 232.050 ;
        RECT 76.950 230.400 118.050 231.600 ;
        RECT 76.950 229.950 79.050 230.400 ;
        RECT 115.950 229.950 118.050 230.400 ;
        RECT 148.950 231.600 151.050 232.050 ;
        RECT 211.950 231.600 214.050 232.050 ;
        RECT 148.950 230.400 214.050 231.600 ;
        RECT 148.950 229.950 151.050 230.400 ;
        RECT 211.950 229.950 214.050 230.400 ;
        RECT 412.950 231.600 415.050 232.050 ;
        RECT 445.950 231.600 448.050 231.900 ;
        RECT 412.950 230.400 448.050 231.600 ;
        RECT 412.950 229.950 415.050 230.400 ;
        RECT 445.950 229.800 448.050 230.400 ;
        RECT 460.950 231.600 463.050 232.050 ;
        RECT 478.950 231.600 481.050 232.050 ;
        RECT 514.950 231.600 517.050 232.050 ;
        RECT 460.950 230.400 481.050 231.600 ;
        RECT 460.950 229.950 463.050 230.400 ;
        RECT 478.950 229.950 481.050 230.400 ;
        RECT 485.400 230.400 517.050 231.600 ;
        RECT 22.950 228.600 25.050 229.050 ;
        RECT 64.950 228.600 67.050 229.050 ;
        RECT 94.950 228.600 97.050 229.050 ;
        RECT 22.950 227.400 97.050 228.600 ;
        RECT 22.950 226.950 25.050 227.400 ;
        RECT 64.950 226.950 67.050 227.400 ;
        RECT 94.950 226.950 97.050 227.400 ;
        RECT 121.950 228.600 124.050 229.050 ;
        RECT 130.950 228.600 133.050 229.050 ;
        RECT 121.950 227.400 133.050 228.600 ;
        RECT 121.950 226.950 124.050 227.400 ;
        RECT 130.950 226.950 133.050 227.400 ;
        RECT 166.950 228.600 169.050 229.050 ;
        RECT 196.950 228.600 199.050 229.050 ;
        RECT 166.950 227.400 199.050 228.600 ;
        RECT 166.950 226.950 169.050 227.400 ;
        RECT 196.950 226.950 199.050 227.400 ;
        RECT 295.950 228.600 298.050 229.050 ;
        RECT 304.950 228.600 307.050 229.050 ;
        RECT 322.950 228.600 325.050 229.050 ;
        RECT 295.950 227.400 325.050 228.600 ;
        RECT 295.950 226.950 298.050 227.400 ;
        RECT 304.950 226.950 307.050 227.400 ;
        RECT 322.950 226.950 325.050 227.400 ;
        RECT 328.950 228.600 331.050 229.050 ;
        RECT 364.950 228.600 367.050 229.050 ;
        RECT 328.950 227.400 367.050 228.600 ;
        RECT 328.950 226.950 331.050 227.400 ;
        RECT 364.950 226.950 367.050 227.400 ;
        RECT 376.950 228.600 379.050 229.050 ;
        RECT 485.400 228.600 486.600 230.400 ;
        RECT 514.950 229.950 517.050 230.400 ;
        RECT 520.950 231.600 523.050 232.050 ;
        RECT 655.950 231.600 658.050 232.050 ;
        RECT 679.950 231.600 682.050 232.050 ;
        RECT 520.950 230.400 682.050 231.600 ;
        RECT 520.950 229.950 523.050 230.400 ;
        RECT 655.950 229.950 658.050 230.400 ;
        RECT 679.950 229.950 682.050 230.400 ;
        RECT 766.950 231.600 769.050 232.050 ;
        RECT 802.950 231.600 805.050 232.050 ;
        RECT 766.950 230.400 805.050 231.600 ;
        RECT 766.950 229.950 769.050 230.400 ;
        RECT 802.950 229.950 805.050 230.400 ;
        RECT 844.950 231.600 847.050 232.050 ;
        RECT 892.950 231.600 895.050 232.050 ;
        RECT 844.950 230.400 895.050 231.600 ;
        RECT 844.950 229.950 847.050 230.400 ;
        RECT 892.950 229.950 895.050 230.400 ;
        RECT 376.950 227.400 486.600 228.600 ;
        RECT 487.950 228.600 490.050 229.050 ;
        RECT 517.950 228.600 520.050 229.050 ;
        RECT 487.950 227.400 520.050 228.600 ;
        RECT 376.950 226.950 379.050 227.400 ;
        RECT 487.950 226.950 490.050 227.400 ;
        RECT 517.950 226.950 520.050 227.400 ;
        RECT 568.950 228.600 571.050 229.050 ;
        RECT 583.950 228.600 586.050 229.050 ;
        RECT 568.950 227.400 586.050 228.600 ;
        RECT 568.950 226.950 571.050 227.400 ;
        RECT 583.950 226.950 586.050 227.400 ;
        RECT 604.950 228.600 607.050 229.050 ;
        RECT 646.950 228.600 649.050 229.050 ;
        RECT 604.950 227.400 649.050 228.600 ;
        RECT 604.950 226.950 607.050 227.400 ;
        RECT 646.950 226.950 649.050 227.400 ;
        RECT 691.950 228.600 694.050 229.050 ;
        RECT 712.950 228.600 715.050 229.050 ;
        RECT 691.950 227.400 715.050 228.600 ;
        RECT 691.950 226.950 694.050 227.400 ;
        RECT 712.950 226.950 715.050 227.400 ;
        RECT 70.950 225.600 73.050 226.050 ;
        RECT 76.950 225.600 79.050 226.050 ;
        RECT 70.950 224.400 79.050 225.600 ;
        RECT 70.950 223.950 73.050 224.400 ;
        RECT 76.950 223.950 79.050 224.400 ;
        RECT 241.950 225.600 244.050 226.050 ;
        RECT 265.950 225.600 268.050 226.050 ;
        RECT 241.950 224.400 268.050 225.600 ;
        RECT 241.950 223.950 244.050 224.400 ;
        RECT 265.950 223.950 268.050 224.400 ;
        RECT 283.950 225.600 286.050 226.050 ;
        RECT 586.950 225.600 589.050 226.050 ;
        RECT 634.950 225.600 637.050 226.050 ;
        RECT 727.950 225.600 730.050 226.050 ;
        RECT 283.950 224.400 730.050 225.600 ;
        RECT 283.950 223.950 286.050 224.400 ;
        RECT 586.950 223.950 589.050 224.400 ;
        RECT 634.950 223.950 637.050 224.400 ;
        RECT 727.950 223.950 730.050 224.400 ;
        RECT 856.950 225.600 859.050 226.050 ;
        RECT 937.950 225.600 940.050 226.050 ;
        RECT 943.950 225.600 946.050 226.050 ;
        RECT 856.950 224.400 946.050 225.600 ;
        RECT 856.950 223.950 859.050 224.400 ;
        RECT 937.950 223.950 940.050 224.400 ;
        RECT 943.950 223.950 946.050 224.400 ;
        RECT 34.950 222.600 37.050 223.050 ;
        RECT 49.950 222.600 52.050 223.050 ;
        RECT 34.950 221.400 52.050 222.600 ;
        RECT 34.950 220.950 37.050 221.400 ;
        RECT 49.950 220.950 52.050 221.400 ;
        RECT 91.950 222.600 94.050 223.050 ;
        RECT 124.950 222.600 127.050 223.050 ;
        RECT 157.950 222.600 160.050 223.050 ;
        RECT 91.950 221.400 160.050 222.600 ;
        RECT 91.950 220.950 94.050 221.400 ;
        RECT 124.950 220.950 127.050 221.400 ;
        RECT 157.950 220.950 160.050 221.400 ;
        RECT 217.950 222.600 220.050 223.050 ;
        RECT 226.950 222.600 229.050 223.050 ;
        RECT 217.950 221.400 229.050 222.600 ;
        RECT 217.950 220.950 220.050 221.400 ;
        RECT 226.950 220.950 229.050 221.400 ;
        RECT 292.950 222.600 295.050 223.050 ;
        RECT 304.950 222.600 307.050 223.050 ;
        RECT 316.950 222.600 319.050 223.050 ;
        RECT 358.950 222.600 361.050 223.050 ;
        RECT 292.950 221.400 361.050 222.600 ;
        RECT 292.950 220.950 295.050 221.400 ;
        RECT 304.950 220.950 307.050 221.400 ;
        RECT 316.950 220.950 319.050 221.400 ;
        RECT 358.950 220.950 361.050 221.400 ;
        RECT 370.950 222.600 373.050 223.050 ;
        RECT 376.950 222.600 379.050 223.050 ;
        RECT 370.950 221.400 379.050 222.600 ;
        RECT 370.950 220.950 373.050 221.400 ;
        RECT 376.950 220.950 379.050 221.400 ;
        RECT 385.950 222.600 388.050 223.050 ;
        RECT 439.950 222.600 442.050 223.050 ;
        RECT 472.950 222.600 475.050 223.050 ;
        RECT 385.950 221.400 429.600 222.600 ;
        RECT 385.950 220.950 388.050 221.400 ;
        RECT 428.400 220.200 429.600 221.400 ;
        RECT 439.950 221.400 475.050 222.600 ;
        RECT 439.950 220.950 442.050 221.400 ;
        RECT 472.950 220.950 475.050 221.400 ;
        RECT 484.950 222.600 487.050 223.050 ;
        RECT 505.950 222.600 508.050 223.050 ;
        RECT 484.950 221.400 508.050 222.600 ;
        RECT 484.950 220.950 487.050 221.400 ;
        RECT 505.950 220.950 508.050 221.400 ;
        RECT 619.950 222.600 622.050 223.050 ;
        RECT 670.950 222.600 673.050 223.050 ;
        RECT 619.950 221.400 673.050 222.600 ;
        RECT 619.950 220.950 622.050 221.400 ;
        RECT 670.950 220.950 673.050 221.400 ;
        RECT 730.950 222.600 733.050 223.050 ;
        RECT 745.950 222.600 748.050 223.050 ;
        RECT 730.950 221.400 748.050 222.600 ;
        RECT 730.950 220.950 733.050 221.400 ;
        RECT 745.950 220.950 748.050 221.400 ;
        RECT 826.950 222.600 829.050 223.050 ;
        RECT 838.950 222.600 841.050 223.050 ;
        RECT 826.950 221.400 841.050 222.600 ;
        RECT 826.950 220.950 829.050 221.400 ;
        RECT 838.950 220.950 841.050 221.400 ;
        RECT 919.950 222.600 922.050 223.050 ;
        RECT 931.950 222.600 934.050 223.050 ;
        RECT 919.950 221.400 934.050 222.600 ;
        RECT 919.950 220.950 922.050 221.400 ;
        RECT 931.950 220.950 934.050 221.400 ;
        RECT 973.950 222.600 976.050 223.050 ;
        RECT 1015.950 222.600 1018.050 223.050 ;
        RECT 973.950 221.400 1018.050 222.600 ;
        RECT 973.950 220.950 976.050 221.400 ;
        RECT 1015.950 220.950 1018.050 221.400 ;
        RECT 145.950 219.600 148.050 220.050 ;
        RECT 166.950 219.600 169.050 220.050 ;
        RECT 145.950 218.400 169.050 219.600 ;
        RECT 145.950 217.950 148.050 218.400 ;
        RECT 166.950 217.950 169.050 218.400 ;
        RECT 199.950 219.600 202.050 220.050 ;
        RECT 214.950 219.600 217.050 220.050 ;
        RECT 199.950 218.400 217.050 219.600 ;
        RECT 199.950 217.950 202.050 218.400 ;
        RECT 214.950 217.950 217.050 218.400 ;
        RECT 244.950 219.600 247.050 220.050 ;
        RECT 244.950 218.400 285.600 219.600 ;
        RECT 244.950 217.950 247.050 218.400 ;
        RECT 284.400 217.200 285.600 218.400 ;
        RECT 319.950 217.950 322.050 220.050 ;
        RECT 427.950 219.750 430.050 220.200 ;
        RECT 436.950 219.750 439.050 220.200 ;
        RECT 427.950 218.550 439.050 219.750 ;
        RECT 427.950 218.100 430.050 218.550 ;
        RECT 436.950 218.100 439.050 218.550 ;
        RECT 478.950 219.600 481.050 220.050 ;
        RECT 487.950 219.600 490.050 220.050 ;
        RECT 511.950 219.600 514.050 220.050 ;
        RECT 478.950 218.400 514.050 219.600 ;
        RECT 478.950 217.950 481.050 218.400 ;
        RECT 487.950 217.950 490.050 218.400 ;
        RECT 511.950 217.950 514.050 218.400 ;
        RECT 517.950 219.750 520.050 220.200 ;
        RECT 523.950 219.750 526.050 220.200 ;
        RECT 517.950 218.550 526.050 219.750 ;
        RECT 517.950 218.100 520.050 218.550 ;
        RECT 523.950 218.100 526.050 218.550 ;
        RECT 682.950 219.600 685.050 220.050 ;
        RECT 691.950 219.600 694.050 220.050 ;
        RECT 775.950 219.600 778.050 220.050 ;
        RECT 682.950 218.400 694.050 219.600 ;
        RECT 682.950 217.950 685.050 218.400 ;
        RECT 691.950 217.950 694.050 218.400 ;
        RECT 770.400 218.400 778.050 219.600 ;
        RECT 16.950 216.750 19.050 217.200 ;
        RECT 31.950 216.750 34.050 217.200 ;
        RECT 16.950 215.550 34.050 216.750 ;
        RECT 16.950 215.100 19.050 215.550 ;
        RECT 31.950 215.100 34.050 215.550 ;
        RECT 85.950 216.600 88.050 217.050 ;
        RECT 103.950 216.750 106.050 217.200 ;
        RECT 112.950 216.750 115.050 217.200 ;
        RECT 103.950 216.600 115.050 216.750 ;
        RECT 85.950 215.550 115.050 216.600 ;
        RECT 85.950 215.400 106.050 215.550 ;
        RECT 85.950 214.950 88.050 215.400 ;
        RECT 103.950 215.100 106.050 215.400 ;
        RECT 112.950 215.100 115.050 215.550 ;
        RECT 133.950 216.600 136.050 217.050 ;
        RECT 139.950 216.750 142.050 217.200 ;
        RECT 151.950 216.750 154.050 217.200 ;
        RECT 139.950 216.600 154.050 216.750 ;
        RECT 133.950 215.550 154.050 216.600 ;
        RECT 133.950 215.400 142.050 215.550 ;
        RECT 133.950 214.950 136.050 215.400 ;
        RECT 139.950 215.100 142.050 215.400 ;
        RECT 151.950 215.100 154.050 215.550 ;
        RECT 160.950 213.600 163.050 217.050 ;
        RECT 178.950 216.750 181.050 217.200 ;
        RECT 193.950 216.750 196.050 217.200 ;
        RECT 178.950 215.550 196.050 216.750 ;
        RECT 178.950 215.100 181.050 215.550 ;
        RECT 193.950 215.100 196.050 215.550 ;
        RECT 271.950 216.750 274.050 217.200 ;
        RECT 277.950 216.750 280.050 217.200 ;
        RECT 271.950 215.550 280.050 216.750 ;
        RECT 271.950 215.100 274.050 215.550 ;
        RECT 277.950 215.100 280.050 215.550 ;
        RECT 283.950 216.750 286.050 217.200 ;
        RECT 289.950 216.750 292.050 217.200 ;
        RECT 283.950 215.550 292.050 216.750 ;
        RECT 283.950 215.100 286.050 215.550 ;
        RECT 289.950 215.100 292.050 215.550 ;
        RECT 155.400 213.000 163.050 213.600 ;
        RECT 155.400 212.400 162.600 213.000 ;
        RECT 10.950 210.600 13.050 211.050 ;
        RECT 19.950 210.600 22.050 210.900 ;
        RECT 10.950 209.400 22.050 210.600 ;
        RECT 10.950 208.950 13.050 209.400 ;
        RECT 19.950 208.800 22.050 209.400 ;
        RECT 58.950 210.600 61.050 211.050 ;
        RECT 88.950 210.600 91.050 210.900 ;
        RECT 58.950 209.400 91.050 210.600 ;
        RECT 58.950 208.950 61.050 209.400 ;
        RECT 88.950 208.800 91.050 209.400 ;
        RECT 115.950 210.600 118.050 210.900 ;
        RECT 124.950 210.600 127.050 211.050 ;
        RECT 115.950 209.400 127.050 210.600 ;
        RECT 115.950 208.800 118.050 209.400 ;
        RECT 124.950 208.950 127.050 209.400 ;
        RECT 136.950 210.600 139.050 210.900 ;
        RECT 155.400 210.600 156.600 212.400 ;
        RECT 136.950 209.400 156.600 210.600 ;
        RECT 157.950 210.450 160.050 210.900 ;
        RECT 163.950 210.450 166.050 210.900 ;
        RECT 136.950 208.800 139.050 209.400 ;
        RECT 157.950 209.250 166.050 210.450 ;
        RECT 157.950 208.800 160.050 209.250 ;
        RECT 163.950 208.800 166.050 209.250 ;
        RECT 175.950 210.600 178.050 211.050 ;
        RECT 190.950 210.600 193.050 210.900 ;
        RECT 175.950 209.400 193.050 210.600 ;
        RECT 175.950 208.950 178.050 209.400 ;
        RECT 190.950 208.800 193.050 209.400 ;
        RECT 241.950 210.600 244.050 210.900 ;
        RECT 253.950 210.600 256.050 211.050 ;
        RECT 268.950 210.600 271.050 210.900 ;
        RECT 241.950 209.400 271.050 210.600 ;
        RECT 241.950 208.800 244.050 209.400 ;
        RECT 253.950 208.950 256.050 209.400 ;
        RECT 268.950 208.800 271.050 209.400 ;
        RECT 298.950 210.450 301.050 210.900 ;
        RECT 304.950 210.450 307.050 210.900 ;
        RECT 298.950 209.250 307.050 210.450 ;
        RECT 320.400 210.600 321.600 217.950 ;
        RECT 322.950 215.100 325.050 217.200 ;
        RECT 340.950 216.750 343.050 217.200 ;
        RECT 355.950 216.750 358.050 217.200 ;
        RECT 340.950 215.550 358.050 216.750 ;
        RECT 340.950 215.100 343.050 215.550 ;
        RECT 355.950 215.100 358.050 215.550 ;
        RECT 466.950 216.750 469.050 217.200 ;
        RECT 475.950 216.750 478.050 217.200 ;
        RECT 466.950 215.550 478.050 216.750 ;
        RECT 466.950 215.100 469.050 215.550 ;
        RECT 475.950 215.100 478.050 215.550 ;
        RECT 493.950 216.750 496.050 217.200 ;
        RECT 499.950 216.750 502.050 217.200 ;
        RECT 493.950 215.550 502.050 216.750 ;
        RECT 493.950 215.100 496.050 215.550 ;
        RECT 499.950 215.100 502.050 215.550 ;
        RECT 589.950 216.600 592.050 217.050 ;
        RECT 607.950 216.600 610.050 217.200 ;
        RECT 589.950 215.400 610.050 216.600 ;
        RECT 323.400 213.600 324.600 215.100 ;
        RECT 589.950 214.950 592.050 215.400 ;
        RECT 607.950 215.100 610.050 215.400 ;
        RECT 634.950 216.750 637.050 217.200 ;
        RECT 643.950 216.750 646.050 217.200 ;
        RECT 634.950 215.550 646.050 216.750 ;
        RECT 634.950 215.100 637.050 215.550 ;
        RECT 643.950 215.100 646.050 215.550 ;
        RECT 661.950 216.750 664.050 217.200 ;
        RECT 667.950 216.750 670.050 217.200 ;
        RECT 661.950 215.550 670.050 216.750 ;
        RECT 661.950 215.100 664.050 215.550 ;
        RECT 667.950 215.100 670.050 215.550 ;
        RECT 685.950 216.600 688.050 217.200 ;
        RECT 697.950 216.600 700.050 217.050 ;
        RECT 685.950 215.400 700.050 216.600 ;
        RECT 685.950 215.100 688.050 215.400 ;
        RECT 697.950 214.950 700.050 215.400 ;
        RECT 703.950 216.750 706.050 217.200 ;
        RECT 718.950 216.750 721.050 217.200 ;
        RECT 703.950 216.600 721.050 216.750 ;
        RECT 724.950 216.600 727.050 217.050 ;
        RECT 736.950 216.600 739.050 217.200 ;
        RECT 703.950 215.550 723.600 216.600 ;
        RECT 703.950 215.100 706.050 215.550 ;
        RECT 718.950 215.400 723.600 215.550 ;
        RECT 718.950 215.100 721.050 215.400 ;
        RECT 547.950 213.600 550.050 214.200 ;
        RECT 722.400 213.600 723.600 215.400 ;
        RECT 724.950 215.400 739.050 216.600 ;
        RECT 724.950 214.950 727.050 215.400 ;
        RECT 736.950 215.100 739.050 215.400 ;
        RECT 745.950 216.600 748.050 217.050 ;
        RECT 751.950 216.750 754.050 217.050 ;
        RECT 760.950 216.750 763.050 217.200 ;
        RECT 751.950 216.600 763.050 216.750 ;
        RECT 745.950 215.550 763.050 216.600 ;
        RECT 745.950 215.400 754.050 215.550 ;
        RECT 745.950 214.950 748.050 215.400 ;
        RECT 751.950 214.950 754.050 215.400 ;
        RECT 760.950 215.100 763.050 215.550 ;
        RECT 751.950 213.600 754.050 213.900 ;
        RECT 323.400 213.000 339.600 213.600 ;
        RECT 323.400 212.400 340.050 213.000 ;
        RECT 320.400 209.400 324.600 210.600 ;
        RECT 298.950 208.800 301.050 209.250 ;
        RECT 304.950 208.800 307.050 209.250 ;
        RECT 323.400 207.600 324.600 209.400 ;
        RECT 337.950 208.950 340.050 212.400 ;
        RECT 547.950 212.400 609.600 213.600 ;
        RECT 722.400 212.400 754.050 213.600 ;
        RECT 547.950 212.100 550.050 212.400 ;
        RECT 343.950 210.600 346.050 210.900 ;
        RECT 352.950 210.600 355.050 211.050 ;
        RECT 343.950 209.400 355.050 210.600 ;
        RECT 343.950 208.800 346.050 209.400 ;
        RECT 352.950 208.950 355.050 209.400 ;
        RECT 361.950 210.600 364.050 211.050 ;
        RECT 367.950 210.600 370.050 210.900 ;
        RECT 361.950 209.400 370.050 210.600 ;
        RECT 361.950 208.950 364.050 209.400 ;
        RECT 367.950 208.800 370.050 209.400 ;
        RECT 445.950 210.600 448.050 211.050 ;
        RECT 463.950 210.600 466.050 210.900 ;
        RECT 445.950 209.400 466.050 210.600 ;
        RECT 445.950 208.950 448.050 209.400 ;
        RECT 463.950 208.800 466.050 209.400 ;
        RECT 472.950 210.600 475.050 211.050 ;
        RECT 490.950 210.600 493.050 210.900 ;
        RECT 472.950 209.400 493.050 210.600 ;
        RECT 472.950 208.950 475.050 209.400 ;
        RECT 490.950 208.800 493.050 209.400 ;
        RECT 598.950 210.450 601.050 210.900 ;
        RECT 604.950 210.450 607.050 210.900 ;
        RECT 598.950 209.250 607.050 210.450 ;
        RECT 608.400 210.600 609.600 212.400 ;
        RECT 751.950 211.800 754.050 212.400 ;
        RECT 631.950 210.600 634.050 210.900 ;
        RECT 608.400 209.400 634.050 210.600 ;
        RECT 598.950 208.800 601.050 209.250 ;
        RECT 604.950 208.800 607.050 209.250 ;
        RECT 631.950 208.800 634.050 209.400 ;
        RECT 658.950 210.600 661.050 210.900 ;
        RECT 703.950 210.600 706.050 211.050 ;
        RECT 658.950 209.400 706.050 210.600 ;
        RECT 658.950 208.800 661.050 209.400 ;
        RECT 703.950 208.950 706.050 209.400 ;
        RECT 715.950 210.450 718.050 210.900 ;
        RECT 724.950 210.450 727.050 210.900 ;
        RECT 715.950 209.250 727.050 210.450 ;
        RECT 715.950 208.800 718.050 209.250 ;
        RECT 724.950 208.800 727.050 209.250 ;
        RECT 739.950 210.450 742.050 210.900 ;
        RECT 745.950 210.450 748.050 210.900 ;
        RECT 739.950 209.250 748.050 210.450 ;
        RECT 770.400 210.600 771.600 218.400 ;
        RECT 775.950 217.950 778.050 218.400 ;
        RECT 823.950 219.750 826.050 220.200 ;
        RECT 862.950 219.750 865.050 220.200 ;
        RECT 823.950 218.550 865.050 219.750 ;
        RECT 823.950 218.100 826.050 218.550 ;
        RECT 862.950 218.100 865.050 218.550 ;
        RECT 952.950 219.600 955.050 220.050 ;
        RECT 964.950 219.600 967.050 220.050 ;
        RECT 952.950 218.400 967.050 219.600 ;
        RECT 952.950 217.950 955.050 218.400 ;
        RECT 964.950 217.950 967.050 218.400 ;
        RECT 886.950 216.600 889.050 217.200 ;
        RECT 949.950 216.600 952.050 217.050 ;
        RECT 961.950 216.600 964.050 217.050 ;
        RECT 976.950 216.600 979.050 217.050 ;
        RECT 886.950 215.400 921.600 216.600 ;
        RECT 886.950 215.100 889.050 215.400 ;
        RECT 772.950 213.450 775.050 213.900 ;
        RECT 787.950 213.450 790.050 213.900 ;
        RECT 772.950 212.250 790.050 213.450 ;
        RECT 772.950 211.800 775.050 212.250 ;
        RECT 787.950 211.800 790.050 212.250 ;
        RECT 886.950 213.600 889.050 214.050 ;
        RECT 910.950 213.600 913.050 214.050 ;
        RECT 886.950 212.400 913.050 213.600 ;
        RECT 920.400 213.600 921.600 215.400 ;
        RECT 949.950 215.400 979.050 216.600 ;
        RECT 949.950 214.950 952.050 215.400 ;
        RECT 961.950 214.950 964.050 215.400 ;
        RECT 976.950 214.950 979.050 215.400 ;
        RECT 982.950 216.600 985.050 217.050 ;
        RECT 994.950 216.600 997.050 217.200 ;
        RECT 982.950 215.400 997.050 216.600 ;
        RECT 982.950 214.950 985.050 215.400 ;
        RECT 994.950 215.100 997.050 215.400 ;
        RECT 1000.950 216.750 1003.050 217.200 ;
        RECT 1021.950 216.750 1024.050 217.200 ;
        RECT 1000.950 215.550 1024.050 216.750 ;
        RECT 1000.950 215.100 1003.050 215.550 ;
        RECT 1021.950 215.100 1024.050 215.550 ;
        RECT 922.950 213.600 925.050 213.900 ;
        RECT 920.400 212.400 925.050 213.600 ;
        RECT 886.950 211.950 889.050 212.400 ;
        RECT 910.950 211.950 913.050 212.400 ;
        RECT 922.950 211.800 925.050 212.400 ;
        RECT 784.950 210.600 787.050 211.050 ;
        RECT 770.400 209.400 787.050 210.600 ;
        RECT 739.950 208.800 742.050 209.250 ;
        RECT 745.950 208.800 748.050 209.250 ;
        RECT 784.950 208.950 787.050 209.400 ;
        RECT 913.950 210.600 916.050 211.050 ;
        RECT 919.950 210.600 922.050 211.050 ;
        RECT 913.950 209.400 922.050 210.600 ;
        RECT 913.950 208.950 916.050 209.400 ;
        RECT 919.950 208.950 922.050 209.400 ;
        RECT 964.950 210.450 967.050 210.900 ;
        RECT 970.950 210.450 973.050 210.900 ;
        RECT 964.950 209.250 973.050 210.450 ;
        RECT 964.950 208.800 967.050 209.250 ;
        RECT 970.950 208.800 973.050 209.250 ;
        RECT 985.950 210.450 988.050 210.900 ;
        RECT 997.950 210.450 1000.050 210.900 ;
        RECT 985.950 209.250 1000.050 210.450 ;
        RECT 985.950 208.800 988.050 209.250 ;
        RECT 997.950 208.800 1000.050 209.250 ;
        RECT 1006.950 210.600 1009.050 211.050 ;
        RECT 1018.950 210.600 1021.050 210.900 ;
        RECT 1006.950 209.400 1021.050 210.600 ;
        RECT 1006.950 208.950 1009.050 209.400 ;
        RECT 1018.950 208.800 1021.050 209.400 ;
        RECT 328.950 207.600 331.050 208.050 ;
        RECT 323.400 206.400 331.050 207.600 ;
        RECT 328.950 205.950 331.050 206.400 ;
        RECT 334.950 207.600 337.050 208.050 ;
        RECT 340.950 207.600 343.050 208.050 ;
        RECT 334.950 206.400 343.050 207.600 ;
        RECT 334.950 205.950 337.050 206.400 ;
        RECT 340.950 205.950 343.050 206.400 ;
        RECT 508.950 207.600 511.050 208.050 ;
        RECT 574.950 207.600 577.050 208.050 ;
        RECT 508.950 206.400 577.050 207.600 ;
        RECT 508.950 205.950 511.050 206.400 ;
        RECT 574.950 205.950 577.050 206.400 ;
        RECT 688.950 207.600 691.050 208.050 ;
        RECT 730.950 207.600 733.050 208.050 ;
        RECT 688.950 206.400 733.050 207.600 ;
        RECT 688.950 205.950 691.050 206.400 ;
        RECT 730.950 205.950 733.050 206.400 ;
        RECT 751.950 207.600 754.050 208.050 ;
        RECT 763.950 207.600 766.050 208.050 ;
        RECT 751.950 206.400 766.050 207.600 ;
        RECT 751.950 205.950 754.050 206.400 ;
        RECT 763.950 205.950 766.050 206.400 ;
        RECT 115.950 204.600 118.050 205.050 ;
        RECT 121.950 204.600 124.050 205.050 ;
        RECT 115.950 203.400 124.050 204.600 ;
        RECT 115.950 202.950 118.050 203.400 ;
        RECT 121.950 202.950 124.050 203.400 ;
        RECT 130.950 204.600 133.050 205.050 ;
        RECT 142.950 204.600 145.050 205.050 ;
        RECT 130.950 203.400 145.050 204.600 ;
        RECT 130.950 202.950 133.050 203.400 ;
        RECT 142.950 202.950 145.050 203.400 ;
        RECT 205.950 204.600 208.050 205.050 ;
        RECT 241.950 204.600 244.050 205.050 ;
        RECT 205.950 203.400 244.050 204.600 ;
        RECT 205.950 202.950 208.050 203.400 ;
        RECT 241.950 202.950 244.050 203.400 ;
        RECT 277.950 204.600 280.050 205.050 ;
        RECT 319.950 204.600 322.050 205.050 ;
        RECT 277.950 203.400 322.050 204.600 ;
        RECT 277.950 202.950 280.050 203.400 ;
        RECT 319.950 202.950 322.050 203.400 ;
        RECT 430.950 204.600 433.050 205.050 ;
        RECT 745.950 204.600 748.050 205.050 ;
        RECT 760.950 204.600 763.050 205.050 ;
        RECT 430.950 203.400 603.600 204.600 ;
        RECT 430.950 202.950 433.050 203.400 ;
        RECT 223.950 201.600 226.050 202.050 ;
        RECT 292.950 201.600 295.050 202.050 ;
        RECT 223.950 200.400 295.050 201.600 ;
        RECT 223.950 199.950 226.050 200.400 ;
        RECT 292.950 199.950 295.050 200.400 ;
        RECT 337.950 201.600 340.050 202.050 ;
        RECT 382.950 201.600 385.050 202.050 ;
        RECT 337.950 200.400 385.050 201.600 ;
        RECT 337.950 199.950 340.050 200.400 ;
        RECT 382.950 199.950 385.050 200.400 ;
        RECT 475.950 201.600 478.050 202.050 ;
        RECT 583.950 201.600 586.050 202.050 ;
        RECT 475.950 200.400 586.050 201.600 ;
        RECT 602.400 201.600 603.600 203.400 ;
        RECT 745.950 203.400 763.050 204.600 ;
        RECT 745.950 202.950 748.050 203.400 ;
        RECT 760.950 202.950 763.050 203.400 ;
        RECT 952.950 204.600 955.050 205.050 ;
        RECT 958.950 204.600 961.050 205.050 ;
        RECT 952.950 203.400 961.050 204.600 ;
        RECT 952.950 202.950 955.050 203.400 ;
        RECT 958.950 202.950 961.050 203.400 ;
        RECT 667.950 201.600 670.050 202.050 ;
        RECT 682.950 201.600 685.050 202.050 ;
        RECT 602.400 200.400 685.050 201.600 ;
        RECT 475.950 199.950 478.050 200.400 ;
        RECT 583.950 199.950 586.050 200.400 ;
        RECT 667.950 199.950 670.050 200.400 ;
        RECT 682.950 199.950 685.050 200.400 ;
        RECT 997.950 201.600 1000.050 202.050 ;
        RECT 1039.950 201.600 1042.050 202.050 ;
        RECT 997.950 200.400 1042.050 201.600 ;
        RECT 997.950 199.950 1000.050 200.400 ;
        RECT 1039.950 199.950 1042.050 200.400 ;
        RECT 103.950 198.600 106.050 199.050 ;
        RECT 139.950 198.600 142.050 199.050 ;
        RECT 103.950 197.400 142.050 198.600 ;
        RECT 103.950 196.950 106.050 197.400 ;
        RECT 139.950 196.950 142.050 197.400 ;
        RECT 169.950 198.600 172.050 199.050 ;
        RECT 211.950 198.600 214.050 199.050 ;
        RECT 169.950 197.400 214.050 198.600 ;
        RECT 169.950 196.950 172.050 197.400 ;
        RECT 211.950 196.950 214.050 197.400 ;
        RECT 313.950 198.600 316.050 199.050 ;
        RECT 325.950 198.600 328.050 199.050 ;
        RECT 313.950 197.400 328.050 198.600 ;
        RECT 313.950 196.950 316.050 197.400 ;
        RECT 325.950 196.950 328.050 197.400 ;
        RECT 358.950 198.600 361.050 199.050 ;
        RECT 394.950 198.600 397.050 199.050 ;
        RECT 358.950 197.400 397.050 198.600 ;
        RECT 358.950 196.950 361.050 197.400 ;
        RECT 394.950 196.950 397.050 197.400 ;
        RECT 427.950 198.600 430.050 199.050 ;
        RECT 433.950 198.600 436.050 199.050 ;
        RECT 427.950 197.400 436.050 198.600 ;
        RECT 427.950 196.950 430.050 197.400 ;
        RECT 433.950 196.950 436.050 197.400 ;
        RECT 442.950 198.600 445.050 199.050 ;
        RECT 454.950 198.600 457.050 199.050 ;
        RECT 484.950 198.600 487.050 199.050 ;
        RECT 442.950 197.400 487.050 198.600 ;
        RECT 442.950 196.950 445.050 197.400 ;
        RECT 454.950 196.950 457.050 197.400 ;
        RECT 484.950 196.950 487.050 197.400 ;
        RECT 526.950 198.600 529.050 199.050 ;
        RECT 619.950 198.600 622.050 199.050 ;
        RECT 526.950 197.400 622.050 198.600 ;
        RECT 526.950 196.950 529.050 197.400 ;
        RECT 619.950 196.950 622.050 197.400 ;
        RECT 751.950 198.600 754.050 199.050 ;
        RECT 757.950 198.600 760.050 199.050 ;
        RECT 751.950 197.400 760.050 198.600 ;
        RECT 751.950 196.950 754.050 197.400 ;
        RECT 757.950 196.950 760.050 197.400 ;
        RECT 991.950 198.600 994.050 199.050 ;
        RECT 1027.950 198.600 1030.050 199.050 ;
        RECT 991.950 197.400 1030.050 198.600 ;
        RECT 991.950 196.950 994.050 197.400 ;
        RECT 1027.950 196.950 1030.050 197.400 ;
        RECT 67.950 195.600 70.050 196.050 ;
        RECT 73.950 195.600 76.050 196.050 ;
        RECT 82.950 195.600 85.050 196.050 ;
        RECT 67.950 194.400 85.050 195.600 ;
        RECT 67.950 193.950 70.050 194.400 ;
        RECT 73.950 193.950 76.050 194.400 ;
        RECT 82.950 193.950 85.050 194.400 ;
        RECT 367.950 195.600 370.050 196.050 ;
        RECT 373.950 195.600 376.050 196.050 ;
        RECT 367.950 194.400 376.050 195.600 ;
        RECT 367.950 193.950 370.050 194.400 ;
        RECT 373.950 193.950 376.050 194.400 ;
        RECT 499.950 195.600 502.050 196.050 ;
        RECT 634.800 195.600 636.900 196.050 ;
        RECT 499.950 194.400 636.900 195.600 ;
        RECT 499.950 193.950 502.050 194.400 ;
        RECT 634.800 193.950 636.900 194.400 ;
        RECT 637.950 195.600 640.050 196.050 ;
        RECT 649.950 195.600 652.050 196.050 ;
        RECT 664.950 195.600 667.050 196.050 ;
        RECT 703.950 195.600 706.050 196.050 ;
        RECT 637.950 194.400 706.050 195.600 ;
        RECT 637.950 193.950 640.050 194.400 ;
        RECT 649.950 193.950 652.050 194.400 ;
        RECT 664.950 193.950 667.050 194.400 ;
        RECT 703.950 193.950 706.050 194.400 ;
        RECT 712.950 195.600 715.050 196.050 ;
        RECT 739.950 195.600 742.050 196.050 ;
        RECT 712.950 194.400 742.050 195.600 ;
        RECT 712.950 193.950 715.050 194.400 ;
        RECT 739.950 193.950 742.050 194.400 ;
        RECT 817.950 195.600 820.050 196.050 ;
        RECT 838.950 195.600 841.050 196.050 ;
        RECT 817.950 194.400 841.050 195.600 ;
        RECT 817.950 193.950 820.050 194.400 ;
        RECT 838.950 193.950 841.050 194.400 ;
        RECT 871.950 195.600 874.050 196.050 ;
        RECT 892.950 195.600 895.050 196.050 ;
        RECT 871.950 194.400 895.050 195.600 ;
        RECT 871.950 193.950 874.050 194.400 ;
        RECT 892.950 193.950 895.050 194.400 ;
        RECT 907.950 195.600 910.050 196.050 ;
        RECT 992.400 195.600 993.600 196.950 ;
        RECT 907.950 194.400 993.600 195.600 ;
        RECT 907.950 193.950 910.050 194.400 ;
        RECT 19.950 192.600 22.050 193.050 ;
        RECT 31.950 192.600 34.050 193.050 ;
        RECT 58.950 192.600 61.050 193.050 ;
        RECT 88.950 192.600 91.050 193.050 ;
        RECT 19.950 191.400 91.050 192.600 ;
        RECT 19.950 190.950 22.050 191.400 ;
        RECT 31.950 190.950 34.050 191.400 ;
        RECT 58.950 190.950 61.050 191.400 ;
        RECT 88.950 190.950 91.050 191.400 ;
        RECT 94.950 192.600 97.050 193.050 ;
        RECT 172.950 192.600 175.050 193.050 ;
        RECT 94.950 191.400 175.050 192.600 ;
        RECT 94.950 190.950 97.050 191.400 ;
        RECT 172.950 190.950 175.050 191.400 ;
        RECT 253.950 192.600 256.050 193.050 ;
        RECT 316.950 192.600 319.050 193.050 ;
        RECT 253.950 191.400 319.050 192.600 ;
        RECT 253.950 190.950 256.050 191.400 ;
        RECT 316.950 190.950 319.050 191.400 ;
        RECT 328.950 192.600 331.050 193.050 ;
        RECT 355.950 192.600 358.050 193.050 ;
        RECT 328.950 191.400 358.050 192.600 ;
        RECT 328.950 190.950 331.050 191.400 ;
        RECT 355.950 190.950 358.050 191.400 ;
        RECT 376.950 192.600 379.050 193.050 ;
        RECT 526.950 192.600 529.050 193.050 ;
        RECT 376.950 191.400 529.050 192.600 ;
        RECT 376.950 190.950 379.050 191.400 ;
        RECT 526.950 190.950 529.050 191.400 ;
        RECT 913.950 192.600 916.050 193.050 ;
        RECT 940.950 192.600 943.050 193.050 ;
        RECT 913.950 191.400 943.050 192.600 ;
        RECT 913.950 190.950 916.050 191.400 ;
        RECT 940.950 190.950 943.050 191.400 ;
        RECT 37.950 189.600 40.050 190.050 ;
        RECT 43.950 189.600 46.050 190.050 ;
        RECT 37.950 188.400 46.050 189.600 ;
        RECT 37.950 187.950 40.050 188.400 ;
        RECT 43.950 187.950 46.050 188.400 ;
        RECT 256.950 189.600 259.050 190.050 ;
        RECT 298.950 189.600 301.050 190.050 ;
        RECT 256.950 188.400 301.050 189.600 ;
        RECT 256.950 187.950 259.050 188.400 ;
        RECT 298.950 187.950 301.050 188.400 ;
        RECT 319.950 189.600 322.050 190.050 ;
        RECT 334.950 189.600 337.050 190.050 ;
        RECT 319.950 188.400 337.050 189.600 ;
        RECT 319.950 187.950 322.050 188.400 ;
        RECT 334.950 187.950 337.050 188.400 ;
        RECT 448.950 189.600 451.050 190.050 ;
        RECT 457.950 189.600 460.050 190.050 ;
        RECT 448.950 188.400 460.050 189.600 ;
        RECT 448.950 187.950 451.050 188.400 ;
        RECT 457.950 187.950 460.050 188.400 ;
        RECT 577.950 189.600 580.050 190.050 ;
        RECT 610.950 189.600 613.050 190.050 ;
        RECT 577.950 188.400 613.050 189.600 ;
        RECT 577.950 187.950 580.050 188.400 ;
        RECT 610.950 187.950 613.050 188.400 ;
        RECT 643.950 189.600 646.050 190.050 ;
        RECT 682.950 189.600 685.050 190.050 ;
        RECT 643.950 188.400 685.050 189.600 ;
        RECT 643.950 187.950 646.050 188.400 ;
        RECT 682.950 187.950 685.050 188.400 ;
        RECT 709.950 189.600 712.050 190.050 ;
        RECT 718.950 189.600 721.050 190.050 ;
        RECT 709.950 188.400 721.050 189.600 ;
        RECT 709.950 187.950 712.050 188.400 ;
        RECT 718.950 187.950 721.050 188.400 ;
        RECT 769.950 189.600 772.050 190.050 ;
        RECT 838.950 189.600 841.050 190.050 ;
        RECT 769.950 188.400 841.050 189.600 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 838.950 187.950 841.050 188.400 ;
        RECT 916.950 189.600 919.050 190.050 ;
        RECT 922.950 189.600 925.050 190.050 ;
        RECT 916.950 188.400 925.050 189.600 ;
        RECT 916.950 187.950 919.050 188.400 ;
        RECT 922.950 187.950 925.050 188.400 ;
        RECT 946.950 189.600 949.050 190.050 ;
        RECT 958.950 189.600 961.050 190.050 ;
        RECT 946.950 188.400 961.050 189.600 ;
        RECT 946.950 187.950 949.050 188.400 ;
        RECT 958.950 187.950 961.050 188.400 ;
        RECT 967.950 189.600 970.050 190.050 ;
        RECT 982.950 189.600 985.050 190.050 ;
        RECT 1000.950 189.600 1003.050 190.050 ;
        RECT 967.950 188.400 1003.050 189.600 ;
        RECT 967.950 187.950 970.050 188.400 ;
        RECT 982.950 187.950 985.050 188.400 ;
        RECT 1000.950 187.950 1003.050 188.400 ;
        RECT 79.950 186.600 82.050 187.050 ;
        RECT 163.950 186.600 166.050 187.050 ;
        RECT 175.950 186.600 178.050 187.050 ;
        RECT 79.950 185.400 178.050 186.600 ;
        RECT 79.950 184.950 82.050 185.400 ;
        RECT 163.950 184.950 166.050 185.400 ;
        RECT 175.950 184.950 178.050 185.400 ;
        RECT 214.950 184.950 217.050 187.050 ;
        RECT 262.950 184.950 265.050 187.050 ;
        RECT 271.950 186.600 274.050 187.050 ;
        RECT 280.950 186.600 283.050 187.050 ;
        RECT 271.950 185.400 283.050 186.600 ;
        RECT 271.950 184.950 274.050 185.400 ;
        RECT 280.950 184.950 283.050 185.400 ;
        RECT 316.950 186.600 319.050 187.050 ;
        RECT 331.950 186.600 334.050 187.050 ;
        RECT 376.950 186.600 379.050 187.050 ;
        RECT 997.950 186.600 1000.050 187.050 ;
        RECT 316.950 185.400 379.050 186.600 ;
        RECT 316.950 184.950 319.050 185.400 ;
        RECT 331.950 184.950 334.050 185.400 ;
        RECT 376.950 184.950 379.050 185.400 ;
        RECT 935.400 185.400 1000.050 186.600 ;
        RECT 25.950 183.600 28.050 184.050 ;
        RECT 34.950 183.600 37.050 184.050 ;
        RECT 25.950 182.400 37.050 183.600 ;
        RECT 25.950 181.950 28.050 182.400 ;
        RECT 34.950 181.950 37.050 182.400 ;
        RECT 52.950 183.600 55.050 184.050 ;
        RECT 67.950 183.600 70.050 184.200 ;
        RECT 52.950 182.400 70.050 183.600 ;
        RECT 52.950 181.950 55.050 182.400 ;
        RECT 67.950 182.100 70.050 182.400 ;
        RECT 94.950 183.750 97.050 184.200 ;
        RECT 100.950 183.750 103.050 184.200 ;
        RECT 94.950 182.550 103.050 183.750 ;
        RECT 94.950 182.100 97.050 182.550 ;
        RECT 100.950 182.100 103.050 182.550 ;
        RECT 181.950 183.600 184.050 184.050 ;
        RECT 190.950 183.600 193.050 184.200 ;
        RECT 181.950 182.400 193.050 183.600 ;
        RECT 181.950 181.950 184.050 182.400 ;
        RECT 190.950 182.100 193.050 182.400 ;
        RECT 215.400 180.600 216.600 184.950 ;
        RECT 217.950 183.750 220.050 184.200 ;
        RECT 253.950 183.750 256.050 184.200 ;
        RECT 217.950 182.550 256.050 183.750 ;
        RECT 217.950 182.100 220.050 182.550 ;
        RECT 253.950 182.100 256.050 182.550 ;
        RECT 179.400 179.400 195.600 180.600 ;
        RECT 215.400 179.400 219.600 180.600 ;
        RECT 46.950 177.450 49.050 177.900 ;
        RECT 52.950 177.450 55.050 177.900 ;
        RECT 46.950 176.250 55.050 177.450 ;
        RECT 46.950 175.800 49.050 176.250 ;
        RECT 52.950 175.800 55.050 176.250 ;
        RECT 58.950 177.450 61.050 177.900 ;
        RECT 64.950 177.450 67.050 177.900 ;
        RECT 58.950 176.250 67.050 177.450 ;
        RECT 58.950 175.800 61.050 176.250 ;
        RECT 64.950 175.800 67.050 176.250 ;
        RECT 70.950 177.450 73.050 177.900 ;
        RECT 82.950 177.450 85.050 178.050 ;
        RECT 100.950 177.450 103.050 177.900 ;
        RECT 70.950 176.250 103.050 177.450 ;
        RECT 70.950 175.800 73.050 176.250 ;
        RECT 82.950 175.950 85.050 176.250 ;
        RECT 100.950 175.800 103.050 176.250 ;
        RECT 169.950 177.600 172.050 177.900 ;
        RECT 179.400 177.600 180.600 179.400 ;
        RECT 169.950 176.400 180.600 177.600 ;
        RECT 194.400 177.600 195.600 179.400 ;
        RECT 214.950 177.600 217.050 177.900 ;
        RECT 194.400 176.400 217.050 177.600 ;
        RECT 218.400 177.600 219.600 179.400 ;
        RECT 223.950 177.600 226.050 178.050 ;
        RECT 263.400 177.900 264.600 184.950 ;
        RECT 935.400 184.200 936.600 185.400 ;
        RECT 997.950 184.950 1000.050 185.400 ;
        RECT 265.950 183.600 268.050 184.200 ;
        RECT 292.950 183.600 295.050 184.200 ;
        RECT 265.950 182.400 295.050 183.600 ;
        RECT 265.950 182.100 268.050 182.400 ;
        RECT 292.950 182.100 295.050 182.400 ;
        RECT 307.950 183.600 310.050 184.050 ;
        RECT 322.950 183.600 325.050 184.200 ;
        RECT 307.950 182.400 325.050 183.600 ;
        RECT 307.950 181.950 310.050 182.400 ;
        RECT 322.950 182.100 325.050 182.400 ;
        RECT 337.950 183.600 340.050 184.050 ;
        RECT 349.950 183.600 352.050 184.200 ;
        RECT 337.950 182.400 352.050 183.600 ;
        RECT 337.950 181.950 340.050 182.400 ;
        RECT 349.950 182.100 352.050 182.400 ;
        RECT 355.950 183.750 358.050 184.200 ;
        RECT 361.950 183.750 364.050 184.200 ;
        RECT 355.950 182.550 364.050 183.750 ;
        RECT 355.950 182.100 358.050 182.550 ;
        RECT 361.950 182.100 364.050 182.550 ;
        RECT 400.950 183.600 403.050 184.200 ;
        RECT 409.950 183.600 412.050 184.050 ;
        RECT 400.950 182.400 412.050 183.600 ;
        RECT 400.950 182.100 403.050 182.400 ;
        RECT 409.950 181.950 412.050 182.400 ;
        RECT 415.950 183.750 418.050 184.200 ;
        RECT 424.950 183.750 427.050 184.200 ;
        RECT 415.950 182.550 427.050 183.750 ;
        RECT 415.950 182.100 418.050 182.550 ;
        RECT 424.950 182.100 427.050 182.550 ;
        RECT 439.950 183.750 442.050 184.200 ;
        RECT 448.950 183.750 451.050 184.200 ;
        RECT 439.950 182.550 451.050 183.750 ;
        RECT 439.950 182.100 442.050 182.550 ;
        RECT 448.950 182.100 451.050 182.550 ;
        RECT 505.950 183.600 508.050 184.050 ;
        RECT 511.950 183.600 514.050 184.050 ;
        RECT 568.950 183.600 571.050 184.050 ;
        RECT 505.950 182.400 571.050 183.600 ;
        RECT 505.950 181.950 508.050 182.400 ;
        RECT 511.950 181.950 514.050 182.400 ;
        RECT 568.950 181.950 571.050 182.400 ;
        RECT 598.950 183.750 601.050 184.200 ;
        RECT 616.950 183.750 619.050 184.200 ;
        RECT 598.950 182.550 619.050 183.750 ;
        RECT 598.950 182.100 601.050 182.550 ;
        RECT 616.950 182.100 619.050 182.550 ;
        RECT 628.950 183.750 631.050 184.200 ;
        RECT 640.950 183.750 643.050 184.200 ;
        RECT 628.950 182.550 643.050 183.750 ;
        RECT 628.950 182.100 631.050 182.550 ;
        RECT 640.950 182.100 643.050 182.550 ;
        RECT 676.950 183.750 679.050 184.200 ;
        RECT 688.950 183.750 691.050 184.200 ;
        RECT 676.950 182.550 691.050 183.750 ;
        RECT 676.950 182.100 679.050 182.550 ;
        RECT 688.950 182.100 691.050 182.550 ;
        RECT 700.950 183.600 703.050 184.050 ;
        RECT 712.950 183.600 715.050 184.200 ;
        RECT 700.950 182.400 715.050 183.600 ;
        RECT 700.950 181.950 703.050 182.400 ;
        RECT 712.950 182.100 715.050 182.400 ;
        RECT 745.950 183.600 748.050 184.200 ;
        RECT 793.950 183.600 796.050 184.200 ;
        RECT 799.950 183.600 802.050 184.050 ;
        RECT 745.950 182.400 802.050 183.600 ;
        RECT 745.950 182.100 748.050 182.400 ;
        RECT 793.950 182.100 796.050 182.400 ;
        RECT 799.950 181.950 802.050 182.400 ;
        RECT 805.950 183.750 808.050 184.200 ;
        RECT 811.950 183.750 814.050 184.200 ;
        RECT 805.950 182.550 814.050 183.750 ;
        RECT 805.950 182.100 808.050 182.550 ;
        RECT 811.950 182.100 814.050 182.550 ;
        RECT 910.950 181.950 913.050 184.050 ;
        RECT 934.950 182.100 937.050 184.200 ;
        RECT 973.950 183.750 976.050 184.200 ;
        RECT 982.950 183.750 985.050 184.200 ;
        RECT 973.950 182.550 985.050 183.750 ;
        RECT 973.950 182.100 976.050 182.550 ;
        RECT 982.950 182.100 985.050 182.550 ;
        RECT 1006.950 183.750 1009.050 184.200 ;
        RECT 1015.950 183.750 1018.050 184.200 ;
        RECT 1006.950 182.550 1018.050 183.750 ;
        RECT 1006.950 182.100 1009.050 182.550 ;
        RECT 1015.950 182.100 1018.050 182.550 ;
        RECT 1021.950 183.600 1024.050 184.200 ;
        RECT 1030.950 183.600 1033.050 184.050 ;
        RECT 1021.950 182.400 1033.050 183.600 ;
        RECT 1021.950 182.100 1024.050 182.400 ;
        RECT 1030.950 181.950 1033.050 182.400 ;
        RECT 802.950 180.750 805.050 181.200 ;
        RECT 823.950 180.750 826.050 181.200 ;
        RECT 802.950 179.550 826.050 180.750 ;
        RECT 802.950 179.100 805.050 179.550 ;
        RECT 823.950 179.100 826.050 179.550 ;
        RECT 218.400 176.400 226.050 177.600 ;
        RECT 169.950 175.800 172.050 176.400 ;
        RECT 214.950 175.800 217.050 176.400 ;
        RECT 223.950 175.950 226.050 176.400 ;
        RECT 244.950 177.450 247.050 177.900 ;
        RECT 256.950 177.450 259.050 177.900 ;
        RECT 244.950 176.250 259.050 177.450 ;
        RECT 244.950 175.800 247.050 176.250 ;
        RECT 256.950 175.800 259.050 176.250 ;
        RECT 262.950 175.800 265.050 177.900 ;
        RECT 310.950 177.450 313.050 177.900 ;
        RECT 319.950 177.450 322.050 177.900 ;
        RECT 310.950 176.250 322.050 177.450 ;
        RECT 310.950 175.800 313.050 176.250 ;
        RECT 319.950 175.800 322.050 176.250 ;
        RECT 325.950 177.450 328.050 177.900 ;
        RECT 334.950 177.600 337.050 177.900 ;
        RECT 352.950 177.600 355.050 177.900 ;
        RECT 451.950 177.600 454.050 177.900 ;
        RECT 334.950 177.450 355.050 177.600 ;
        RECT 325.950 176.400 355.050 177.450 ;
        RECT 325.950 176.250 337.050 176.400 ;
        RECT 325.950 175.800 328.050 176.250 ;
        RECT 334.950 175.800 337.050 176.250 ;
        RECT 352.950 175.800 355.050 176.400 ;
        RECT 422.400 176.400 454.050 177.600 ;
        RECT 16.950 174.600 19.050 175.050 ;
        RECT 28.950 174.600 31.050 175.050 ;
        RECT 16.950 173.400 31.050 174.600 ;
        RECT 16.950 172.950 19.050 173.400 ;
        RECT 28.950 172.950 31.050 173.400 ;
        RECT 109.950 174.600 112.050 175.050 ;
        RECT 127.950 174.600 130.050 175.050 ;
        RECT 109.950 173.400 130.050 174.600 ;
        RECT 109.950 172.950 112.050 173.400 ;
        RECT 127.950 172.950 130.050 173.400 ;
        RECT 181.950 174.600 184.050 175.050 ;
        RECT 220.950 174.600 223.050 175.050 ;
        RECT 181.950 173.400 223.050 174.600 ;
        RECT 181.950 172.950 184.050 173.400 ;
        RECT 220.950 172.950 223.050 173.400 ;
        RECT 232.950 174.600 235.050 175.050 ;
        RECT 238.950 174.600 241.050 175.050 ;
        RECT 232.950 173.400 241.050 174.600 ;
        RECT 232.950 172.950 235.050 173.400 ;
        RECT 238.950 172.950 241.050 173.400 ;
        RECT 403.950 174.600 406.050 175.050 ;
        RECT 415.950 174.600 418.050 175.050 ;
        RECT 422.400 174.600 423.600 176.400 ;
        RECT 451.950 175.800 454.050 176.400 ;
        RECT 514.950 177.600 517.050 178.050 ;
        RECT 544.950 177.600 547.050 177.900 ;
        RECT 514.950 176.400 547.050 177.600 ;
        RECT 514.950 175.950 517.050 176.400 ;
        RECT 544.950 175.800 547.050 176.400 ;
        RECT 613.950 177.600 616.050 177.900 ;
        RECT 628.950 177.600 631.050 178.050 ;
        RECT 613.950 176.400 631.050 177.600 ;
        RECT 613.950 175.800 616.050 176.400 ;
        RECT 628.950 175.950 631.050 176.400 ;
        RECT 649.950 177.450 652.050 177.900 ;
        RECT 661.950 177.450 664.050 177.900 ;
        RECT 649.950 176.250 664.050 177.450 ;
        RECT 649.950 175.800 652.050 176.250 ;
        RECT 661.950 175.800 664.050 176.250 ;
        RECT 691.950 177.450 694.050 177.900 ;
        RECT 700.950 177.450 703.050 177.900 ;
        RECT 691.950 176.250 703.050 177.450 ;
        RECT 691.950 175.800 694.050 176.250 ;
        RECT 700.950 175.800 703.050 176.250 ;
        RECT 772.950 177.600 775.050 177.900 ;
        RECT 790.950 177.600 793.050 177.900 ;
        RECT 772.950 176.400 793.050 177.600 ;
        RECT 772.950 175.800 775.050 176.400 ;
        RECT 790.950 175.800 793.050 176.400 ;
        RECT 838.950 177.600 841.050 178.050 ;
        RECT 859.950 177.600 862.050 178.050 ;
        RECT 838.950 176.400 862.050 177.600 ;
        RECT 911.400 177.600 912.600 181.950 ;
        RECT 1000.950 180.600 1003.050 181.050 ;
        RECT 1000.950 179.400 1020.600 180.600 ;
        RECT 1000.950 178.950 1003.050 179.400 ;
        RECT 913.950 177.600 916.050 177.900 ;
        RECT 911.400 176.400 916.050 177.600 ;
        RECT 838.950 175.950 841.050 176.400 ;
        RECT 859.950 175.950 862.050 176.400 ;
        RECT 913.950 175.800 916.050 176.400 ;
        RECT 949.950 177.600 952.050 177.900 ;
        RECT 970.950 177.600 973.050 177.900 ;
        RECT 949.950 176.400 973.050 177.600 ;
        RECT 949.950 175.800 952.050 176.400 ;
        RECT 970.950 175.800 973.050 176.400 ;
        RECT 982.950 177.600 985.050 178.050 ;
        RECT 1019.400 177.900 1020.600 179.400 ;
        RECT 991.950 177.600 994.050 177.900 ;
        RECT 982.950 176.400 994.050 177.600 ;
        RECT 982.950 175.950 985.050 176.400 ;
        RECT 991.950 175.800 994.050 176.400 ;
        RECT 1003.950 177.450 1006.050 177.900 ;
        RECT 1012.950 177.450 1015.050 177.900 ;
        RECT 1003.950 176.250 1015.050 177.450 ;
        RECT 1003.950 175.800 1006.050 176.250 ;
        RECT 1012.950 175.800 1015.050 176.250 ;
        RECT 1018.950 175.800 1021.050 177.900 ;
        RECT 403.950 173.400 423.600 174.600 ;
        RECT 637.950 174.600 640.050 175.050 ;
        RECT 685.950 174.600 688.050 175.050 ;
        RECT 637.950 173.400 688.050 174.600 ;
        RECT 403.950 172.950 406.050 173.400 ;
        RECT 415.950 172.950 418.050 173.400 ;
        RECT 637.950 172.950 640.050 173.400 ;
        RECT 685.950 172.950 688.050 173.400 ;
        RECT 40.950 171.600 43.050 172.050 ;
        RECT 91.950 171.600 94.050 172.050 ;
        RECT 40.950 170.400 94.050 171.600 ;
        RECT 40.950 169.950 43.050 170.400 ;
        RECT 91.950 169.950 94.050 170.400 ;
        RECT 139.950 171.600 142.050 172.050 ;
        RECT 148.950 171.600 151.050 172.050 ;
        RECT 139.950 170.400 151.050 171.600 ;
        RECT 139.950 169.950 142.050 170.400 ;
        RECT 148.950 169.950 151.050 170.400 ;
        RECT 187.950 171.600 190.050 171.900 ;
        RECT 239.400 171.600 240.600 172.950 ;
        RECT 274.950 171.600 277.050 172.050 ;
        RECT 187.950 170.400 216.600 171.600 ;
        RECT 239.400 170.400 277.050 171.600 ;
        RECT 187.950 169.800 190.050 170.400 ;
        RECT 91.950 168.600 94.050 168.900 ;
        RECT 106.950 168.600 109.050 169.050 ;
        RECT 91.950 167.400 109.050 168.600 ;
        RECT 215.400 168.600 216.600 170.400 ;
        RECT 274.950 169.950 277.050 170.400 ;
        RECT 301.950 171.600 304.050 172.050 ;
        RECT 337.950 171.600 340.050 172.050 ;
        RECT 301.950 170.400 340.050 171.600 ;
        RECT 301.950 169.950 304.050 170.400 ;
        RECT 337.950 169.950 340.050 170.400 ;
        RECT 385.950 171.600 388.050 172.050 ;
        RECT 433.950 171.600 436.050 172.050 ;
        RECT 385.950 170.400 436.050 171.600 ;
        RECT 385.950 169.950 388.050 170.400 ;
        RECT 433.950 169.950 436.050 170.400 ;
        RECT 586.950 171.600 589.050 172.050 ;
        RECT 601.950 171.600 604.050 172.050 ;
        RECT 638.400 171.600 639.600 172.950 ;
        RECT 586.950 170.400 639.600 171.600 ;
        RECT 643.950 171.600 646.050 172.050 ;
        RECT 676.950 171.600 679.050 172.050 ;
        RECT 643.950 170.400 679.050 171.600 ;
        RECT 586.950 169.950 589.050 170.400 ;
        RECT 601.950 169.950 604.050 170.400 ;
        RECT 643.950 169.950 646.050 170.400 ;
        RECT 676.950 169.950 679.050 170.400 ;
        RECT 814.950 171.600 817.050 172.050 ;
        RECT 892.950 171.600 895.050 172.050 ;
        RECT 814.950 170.400 895.050 171.600 ;
        RECT 814.950 169.950 817.050 170.400 ;
        RECT 892.950 169.950 895.050 170.400 ;
        RECT 928.950 171.600 931.050 172.050 ;
        RECT 1006.950 171.600 1009.050 172.050 ;
        RECT 928.950 170.400 1009.050 171.600 ;
        RECT 928.950 169.950 931.050 170.400 ;
        RECT 1006.950 169.950 1009.050 170.400 ;
        RECT 289.950 168.600 292.050 169.050 ;
        RECT 302.400 168.600 303.600 169.950 ;
        RECT 215.400 167.400 303.600 168.600 ;
        RECT 379.950 168.600 382.050 169.050 ;
        RECT 445.950 168.600 448.050 169.050 ;
        RECT 460.950 168.600 463.050 169.050 ;
        RECT 379.950 167.400 463.050 168.600 ;
        RECT 91.950 166.800 94.050 167.400 ;
        RECT 106.950 166.950 109.050 167.400 ;
        RECT 289.950 166.950 292.050 167.400 ;
        RECT 379.950 166.950 382.050 167.400 ;
        RECT 445.950 166.950 448.050 167.400 ;
        RECT 460.950 166.950 463.050 167.400 ;
        RECT 700.950 168.600 703.050 169.050 ;
        RECT 805.950 168.600 808.050 169.050 ;
        RECT 700.950 167.400 808.050 168.600 ;
        RECT 700.950 166.950 703.050 167.400 ;
        RECT 805.950 166.950 808.050 167.400 ;
        RECT 979.950 168.600 982.050 169.050 ;
        RECT 1000.950 168.600 1003.050 169.050 ;
        RECT 979.950 167.400 1003.050 168.600 ;
        RECT 979.950 166.950 982.050 167.400 ;
        RECT 1000.950 166.950 1003.050 167.400 ;
        RECT 160.950 165.600 163.050 166.050 ;
        RECT 169.950 165.600 172.050 166.050 ;
        RECT 193.950 165.600 196.050 166.050 ;
        RECT 160.950 164.400 196.050 165.600 ;
        RECT 160.950 163.950 163.050 164.400 ;
        RECT 169.950 163.950 172.050 164.400 ;
        RECT 193.950 163.950 196.050 164.400 ;
        RECT 211.950 165.600 214.050 166.050 ;
        RECT 223.950 165.600 226.050 166.050 ;
        RECT 211.950 164.400 226.050 165.600 ;
        RECT 211.950 163.950 214.050 164.400 ;
        RECT 223.950 163.950 226.050 164.400 ;
        RECT 253.950 165.600 256.050 166.050 ;
        RECT 268.950 165.600 271.050 166.050 ;
        RECT 253.950 164.400 271.050 165.600 ;
        RECT 253.950 163.950 256.050 164.400 ;
        RECT 268.950 163.950 271.050 164.400 ;
        RECT 301.950 165.600 304.050 165.900 ;
        RECT 346.950 165.600 349.050 166.050 ;
        RECT 367.950 165.600 370.050 166.050 ;
        RECT 376.950 165.600 379.050 166.050 ;
        RECT 301.950 164.400 379.050 165.600 ;
        RECT 301.950 163.800 304.050 164.400 ;
        RECT 346.950 163.950 349.050 164.400 ;
        RECT 367.950 163.950 370.050 164.400 ;
        RECT 376.950 163.950 379.050 164.400 ;
        RECT 382.950 165.600 385.050 166.050 ;
        RECT 427.950 165.600 430.050 166.050 ;
        RECT 382.950 164.400 430.050 165.600 ;
        RECT 382.950 163.950 385.050 164.400 ;
        RECT 427.950 163.950 430.050 164.400 ;
        RECT 433.950 165.600 436.050 166.050 ;
        RECT 514.950 165.600 517.050 166.050 ;
        RECT 433.950 164.400 517.050 165.600 ;
        RECT 433.950 163.950 436.050 164.400 ;
        RECT 514.950 163.950 517.050 164.400 ;
        RECT 568.950 165.600 571.050 166.050 ;
        RECT 655.950 165.600 658.050 166.050 ;
        RECT 568.950 164.400 658.050 165.600 ;
        RECT 568.950 163.950 571.050 164.400 ;
        RECT 655.950 163.950 658.050 164.400 ;
        RECT 697.950 165.600 700.050 166.050 ;
        RECT 766.950 165.600 769.050 166.050 ;
        RECT 697.950 164.400 769.050 165.600 ;
        RECT 697.950 163.950 700.050 164.400 ;
        RECT 766.950 163.950 769.050 164.400 ;
        RECT 1006.950 165.600 1009.050 166.050 ;
        RECT 1024.950 165.600 1027.050 166.050 ;
        RECT 1006.950 164.400 1027.050 165.600 ;
        RECT 1006.950 163.950 1009.050 164.400 ;
        RECT 1024.950 163.950 1027.050 164.400 ;
        RECT 178.950 162.600 181.050 163.050 ;
        RECT 196.950 162.600 199.050 163.050 ;
        RECT 178.950 161.400 199.050 162.600 ;
        RECT 178.950 160.950 181.050 161.400 ;
        RECT 196.950 160.950 199.050 161.400 ;
        RECT 538.950 162.600 541.050 163.050 ;
        RECT 658.950 162.600 661.050 163.050 ;
        RECT 538.950 161.400 661.050 162.600 ;
        RECT 538.950 160.950 541.050 161.400 ;
        RECT 658.950 160.950 661.050 161.400 ;
        RECT 931.950 162.600 934.050 163.050 ;
        RECT 1027.950 162.600 1030.050 163.050 ;
        RECT 931.950 161.400 1030.050 162.600 ;
        RECT 931.950 160.950 934.050 161.400 ;
        RECT 1027.950 160.950 1030.050 161.400 ;
        RECT 346.950 159.600 349.050 160.050 ;
        RECT 358.950 159.600 361.050 160.050 ;
        RECT 346.950 158.400 361.050 159.600 ;
        RECT 346.950 157.950 349.050 158.400 ;
        RECT 358.950 157.950 361.050 158.400 ;
        RECT 619.950 159.600 622.050 160.050 ;
        RECT 709.950 159.600 712.050 160.050 ;
        RECT 619.950 158.400 712.050 159.600 ;
        RECT 619.950 157.950 622.050 158.400 ;
        RECT 709.950 157.950 712.050 158.400 ;
        RECT 778.950 159.600 781.050 160.050 ;
        RECT 829.950 159.600 832.050 160.050 ;
        RECT 778.950 158.400 832.050 159.600 ;
        RECT 778.950 157.950 781.050 158.400 ;
        RECT 829.950 157.950 832.050 158.400 ;
        RECT 868.950 159.600 871.050 160.050 ;
        RECT 976.950 159.600 979.050 160.050 ;
        RECT 868.950 158.400 979.050 159.600 ;
        RECT 868.950 157.950 871.050 158.400 ;
        RECT 976.950 157.950 979.050 158.400 ;
        RECT 76.950 156.600 79.050 157.050 ;
        RECT 118.950 156.600 121.050 157.050 ;
        RECT 76.950 155.400 121.050 156.600 ;
        RECT 76.950 154.950 79.050 155.400 ;
        RECT 118.950 154.950 121.050 155.400 ;
        RECT 298.950 156.600 301.050 157.050 ;
        RECT 439.950 156.600 442.050 157.050 ;
        RECT 298.950 155.400 442.050 156.600 ;
        RECT 298.950 154.950 301.050 155.400 ;
        RECT 439.950 154.950 442.050 155.400 ;
        RECT 517.950 156.600 520.050 157.050 ;
        RECT 577.950 156.600 580.050 157.050 ;
        RECT 613.950 156.600 616.050 157.050 ;
        RECT 517.950 155.400 616.050 156.600 ;
        RECT 517.950 154.950 520.050 155.400 ;
        RECT 577.950 154.950 580.050 155.400 ;
        RECT 613.950 154.950 616.050 155.400 ;
        RECT 631.950 156.600 634.050 157.050 ;
        RECT 643.950 156.600 646.050 157.050 ;
        RECT 631.950 155.400 646.050 156.600 ;
        RECT 631.950 154.950 634.050 155.400 ;
        RECT 643.950 154.950 646.050 155.400 ;
        RECT 673.950 156.600 676.050 157.050 ;
        RECT 736.950 156.600 739.050 157.050 ;
        RECT 673.950 155.400 739.050 156.600 ;
        RECT 673.950 154.950 676.050 155.400 ;
        RECT 736.950 154.950 739.050 155.400 ;
        RECT 925.950 156.600 928.050 157.050 ;
        RECT 943.950 156.600 946.050 157.050 ;
        RECT 925.950 155.400 946.050 156.600 ;
        RECT 925.950 154.950 928.050 155.400 ;
        RECT 943.950 154.950 946.050 155.400 ;
        RECT 244.950 153.600 247.050 154.050 ;
        RECT 283.950 153.600 286.050 154.050 ;
        RECT 349.950 153.600 352.050 154.050 ;
        RECT 244.950 152.400 352.050 153.600 ;
        RECT 244.950 151.950 247.050 152.400 ;
        RECT 283.950 151.950 286.050 152.400 ;
        RECT 349.950 151.950 352.050 152.400 ;
        RECT 361.950 153.600 364.050 154.050 ;
        RECT 361.950 152.400 525.600 153.600 ;
        RECT 361.950 151.950 364.050 152.400 ;
        RECT 350.400 150.600 351.600 151.950 ;
        RECT 442.950 150.600 445.050 151.050 ;
        RECT 514.950 150.600 517.050 151.050 ;
        RECT 350.400 149.400 517.050 150.600 ;
        RECT 524.400 150.600 525.600 152.400 ;
        RECT 553.950 150.600 556.050 151.050 ;
        RECT 524.400 149.400 556.050 150.600 ;
        RECT 442.950 148.950 445.050 149.400 ;
        RECT 514.950 148.950 517.050 149.400 ;
        RECT 553.950 148.950 556.050 149.400 ;
        RECT 592.950 150.600 595.050 151.050 ;
        RECT 631.950 150.600 634.050 151.050 ;
        RECT 592.950 149.400 634.050 150.600 ;
        RECT 592.950 148.950 595.050 149.400 ;
        RECT 631.950 148.950 634.050 149.400 ;
        RECT 703.950 150.600 706.050 151.050 ;
        RECT 715.950 150.600 718.050 151.050 ;
        RECT 703.950 149.400 718.050 150.600 ;
        RECT 703.950 148.950 706.050 149.400 ;
        RECT 715.950 148.950 718.050 149.400 ;
        RECT 820.950 150.600 823.050 151.050 ;
        RECT 880.950 150.600 883.050 151.050 ;
        RECT 820.950 149.400 883.050 150.600 ;
        RECT 820.950 148.950 823.050 149.400 ;
        RECT 880.950 148.950 883.050 149.400 ;
        RECT 949.950 150.600 952.050 151.050 ;
        RECT 961.950 150.600 964.050 151.050 ;
        RECT 949.950 149.400 964.050 150.600 ;
        RECT 949.950 148.950 952.050 149.400 ;
        RECT 961.950 148.950 964.050 149.400 ;
        RECT 100.950 147.600 103.050 148.050 ;
        RECT 118.950 147.600 121.050 148.050 ;
        RECT 100.950 146.400 121.050 147.600 ;
        RECT 100.950 145.950 103.050 146.400 ;
        RECT 118.950 145.950 121.050 146.400 ;
        RECT 271.950 147.600 274.050 148.050 ;
        RECT 382.950 147.600 385.050 148.050 ;
        RECT 271.950 146.400 385.050 147.600 ;
        RECT 271.950 145.950 274.050 146.400 ;
        RECT 382.950 145.950 385.050 146.400 ;
        RECT 451.950 147.600 454.050 148.050 ;
        RECT 493.950 147.600 496.050 148.050 ;
        RECT 451.950 146.400 496.050 147.600 ;
        RECT 451.950 145.950 454.050 146.400 ;
        RECT 493.950 145.950 496.050 146.400 ;
        RECT 598.950 147.600 601.050 148.050 ;
        RECT 628.950 147.600 631.050 148.050 ;
        RECT 598.950 146.400 631.050 147.600 ;
        RECT 598.950 145.950 601.050 146.400 ;
        RECT 628.950 145.950 631.050 146.400 ;
        RECT 634.950 147.600 637.050 148.050 ;
        RECT 700.950 147.600 703.050 148.050 ;
        RECT 634.950 146.400 703.050 147.600 ;
        RECT 634.950 145.950 637.050 146.400 ;
        RECT 700.950 145.950 703.050 146.400 ;
        RECT 727.950 147.600 730.050 148.050 ;
        RECT 796.950 147.600 799.050 148.050 ;
        RECT 727.950 146.400 799.050 147.600 ;
        RECT 727.950 145.950 730.050 146.400 ;
        RECT 796.950 145.950 799.050 146.400 ;
        RECT 886.950 147.600 889.050 148.050 ;
        RECT 907.950 147.600 910.050 148.050 ;
        RECT 886.950 146.400 910.050 147.600 ;
        RECT 886.950 145.950 889.050 146.400 ;
        RECT 907.950 145.950 910.050 146.400 ;
        RECT 916.950 147.600 919.050 148.050 ;
        RECT 928.950 147.600 931.050 148.050 ;
        RECT 916.950 146.400 931.050 147.600 ;
        RECT 916.950 145.950 919.050 146.400 ;
        RECT 928.950 145.950 931.050 146.400 ;
        RECT 958.950 147.600 961.050 148.050 ;
        RECT 1012.950 147.600 1015.050 148.050 ;
        RECT 958.950 146.400 1015.050 147.600 ;
        RECT 958.950 145.950 961.050 146.400 ;
        RECT 1012.950 145.950 1015.050 146.400 ;
        RECT 28.950 144.600 31.050 145.050 ;
        RECT 76.950 144.600 79.050 145.050 ;
        RECT 28.950 143.400 79.050 144.600 ;
        RECT 28.950 142.950 31.050 143.400 ;
        RECT 76.950 142.950 79.050 143.400 ;
        RECT 235.950 144.600 238.050 145.050 ;
        RECT 247.950 144.600 250.050 145.050 ;
        RECT 262.950 144.600 265.050 145.050 ;
        RECT 235.950 143.400 265.050 144.600 ;
        RECT 235.950 142.950 238.050 143.400 ;
        RECT 247.950 142.950 250.050 143.400 ;
        RECT 262.950 142.950 265.050 143.400 ;
        RECT 319.950 144.600 322.050 145.050 ;
        RECT 367.950 144.600 370.050 145.050 ;
        RECT 385.950 144.600 388.050 145.050 ;
        RECT 319.950 143.400 388.050 144.600 ;
        RECT 319.950 142.950 322.050 143.400 ;
        RECT 367.950 142.950 370.050 143.400 ;
        RECT 385.950 142.950 388.050 143.400 ;
        RECT 397.950 144.600 400.050 145.050 ;
        RECT 505.950 144.600 508.050 145.050 ;
        RECT 397.950 143.400 508.050 144.600 ;
        RECT 397.950 142.950 400.050 143.400 ;
        RECT 505.950 142.950 508.050 143.400 ;
        RECT 604.950 144.600 607.050 145.050 ;
        RECT 628.950 144.600 631.050 144.900 ;
        RECT 679.950 144.600 682.050 145.050 ;
        RECT 604.950 143.400 682.050 144.600 ;
        RECT 604.950 142.950 607.050 143.400 ;
        RECT 628.950 142.800 631.050 143.400 ;
        RECT 679.950 142.950 682.050 143.400 ;
        RECT 712.950 144.600 715.050 145.050 ;
        RECT 811.950 144.600 814.050 145.050 ;
        RECT 712.950 143.400 814.050 144.600 ;
        RECT 712.950 142.950 715.050 143.400 ;
        RECT 811.950 142.950 814.050 143.400 ;
        RECT 874.950 144.600 877.050 145.050 ;
        RECT 883.950 144.600 886.050 145.050 ;
        RECT 874.950 143.400 886.050 144.600 ;
        RECT 874.950 142.950 877.050 143.400 ;
        RECT 883.950 142.950 886.050 143.400 ;
        RECT 967.950 144.600 970.050 145.050 ;
        RECT 985.950 144.600 988.050 145.050 ;
        RECT 967.950 143.400 996.600 144.600 ;
        RECT 967.950 142.950 970.050 143.400 ;
        RECT 985.950 142.950 988.050 143.400 ;
        RECT 79.950 141.600 82.050 142.050 ;
        RECT 85.950 141.600 88.050 142.050 ;
        RECT 79.950 140.400 88.050 141.600 ;
        RECT 79.950 139.950 82.050 140.400 ;
        RECT 85.950 139.950 88.050 140.400 ;
        RECT 995.400 139.200 996.600 143.400 ;
        RECT 997.950 141.600 1000.050 142.050 ;
        RECT 1018.950 141.600 1021.050 142.050 ;
        RECT 997.950 140.400 1021.050 141.600 ;
        RECT 997.950 139.950 1000.050 140.400 ;
        RECT 1018.950 139.950 1021.050 140.400 ;
        RECT 19.950 138.750 22.050 139.200 ;
        RECT 31.950 138.750 34.050 139.200 ;
        RECT 19.950 137.550 34.050 138.750 ;
        RECT 19.950 137.100 22.050 137.550 ;
        RECT 31.950 137.100 34.050 137.550 ;
        RECT 40.950 138.750 43.050 139.200 ;
        RECT 52.950 138.750 55.050 139.200 ;
        RECT 40.950 137.550 55.050 138.750 ;
        RECT 40.950 137.100 43.050 137.550 ;
        RECT 52.950 137.100 55.050 137.550 ;
        RECT 64.950 138.750 67.050 139.200 ;
        RECT 70.950 138.750 73.050 139.200 ;
        RECT 64.950 137.550 73.050 138.750 ;
        RECT 64.950 137.100 67.050 137.550 ;
        RECT 70.950 137.100 73.050 137.550 ;
        RECT 97.950 138.600 100.050 139.200 ;
        RECT 130.950 138.600 133.050 139.200 ;
        RECT 97.950 137.400 133.050 138.600 ;
        RECT 97.950 137.100 100.050 137.400 ;
        RECT 130.950 137.100 133.050 137.400 ;
        RECT 229.950 136.950 232.050 139.050 ;
        RECT 256.950 138.750 259.050 139.200 ;
        RECT 274.950 138.750 277.050 139.200 ;
        RECT 256.950 137.550 277.050 138.750 ;
        RECT 256.950 137.100 259.050 137.550 ;
        RECT 274.950 137.100 277.050 137.550 ;
        RECT 283.950 137.100 286.050 139.200 ;
        RECT 325.950 138.750 328.050 139.200 ;
        RECT 334.950 138.750 337.050 139.200 ;
        RECT 325.950 137.550 337.050 138.750 ;
        RECT 325.950 137.100 328.050 137.550 ;
        RECT 334.950 137.100 337.050 137.550 ;
        RECT 370.950 138.600 373.050 139.050 ;
        RECT 379.950 138.600 382.050 139.200 ;
        RECT 370.950 137.400 382.050 138.600 ;
        RECT 28.950 132.600 31.050 132.900 ;
        RECT 40.950 132.600 43.050 133.050 ;
        RECT 28.950 131.400 43.050 132.600 ;
        RECT 28.950 130.800 31.050 131.400 ;
        RECT 40.950 130.950 43.050 131.400 ;
        RECT 49.950 132.600 52.050 132.900 ;
        RECT 64.950 132.600 67.050 133.050 ;
        RECT 49.950 131.400 67.050 132.600 ;
        RECT 49.950 130.800 52.050 131.400 ;
        RECT 64.950 130.950 67.050 131.400 ;
        RECT 100.950 132.600 103.050 132.900 ;
        RECT 112.800 132.600 114.900 133.050 ;
        RECT 100.950 131.400 114.900 132.600 ;
        RECT 100.950 130.800 103.050 131.400 ;
        RECT 112.800 130.950 114.900 131.400 ;
        RECT 115.950 132.600 118.050 133.050 ;
        RECT 124.950 132.600 127.050 132.900 ;
        RECT 115.950 131.400 127.050 132.600 ;
        RECT 115.950 130.950 118.050 131.400 ;
        RECT 124.950 130.800 127.050 131.400 ;
        RECT 133.950 132.600 136.050 133.050 ;
        RECT 184.950 132.600 187.050 132.900 ;
        RECT 133.950 131.400 187.050 132.600 ;
        RECT 133.950 130.950 136.050 131.400 ;
        RECT 184.950 130.800 187.050 131.400 ;
        RECT 190.950 132.450 193.050 132.900 ;
        RECT 202.950 132.450 205.050 132.900 ;
        RECT 190.950 131.250 205.050 132.450 ;
        RECT 230.400 132.600 231.600 136.950 ;
        RECT 284.400 135.600 285.600 137.100 ;
        RECT 370.950 136.950 373.050 137.400 ;
        RECT 379.950 137.100 382.050 137.400 ;
        RECT 406.950 138.600 409.050 139.200 ;
        RECT 421.950 138.600 424.050 139.050 ;
        RECT 406.950 137.400 424.050 138.600 ;
        RECT 406.950 137.100 409.050 137.400 ;
        RECT 421.950 136.950 424.050 137.400 ;
        RECT 427.950 138.600 430.050 139.200 ;
        RECT 463.950 138.600 466.050 139.050 ;
        RECT 472.950 138.600 475.050 139.200 ;
        RECT 427.950 137.400 466.050 138.600 ;
        RECT 427.950 137.100 430.050 137.400 ;
        RECT 463.950 136.950 466.050 137.400 ;
        RECT 470.400 137.400 475.050 138.600 ;
        RECT 275.400 134.400 285.600 135.600 ;
        RECT 232.950 132.600 235.050 132.900 ;
        RECT 230.400 131.400 235.050 132.600 ;
        RECT 190.950 130.800 193.050 131.250 ;
        RECT 202.950 130.800 205.050 131.250 ;
        RECT 232.950 130.800 235.050 131.400 ;
        RECT 265.950 132.600 268.050 132.900 ;
        RECT 275.400 132.600 276.600 134.400 ;
        RECT 265.950 131.400 276.600 132.600 ;
        RECT 277.950 132.600 280.050 133.050 ;
        RECT 286.950 132.600 289.050 132.900 ;
        RECT 277.950 131.400 289.050 132.600 ;
        RECT 265.950 130.800 268.050 131.400 ;
        RECT 277.950 130.950 280.050 131.400 ;
        RECT 286.950 130.800 289.050 131.400 ;
        RECT 337.950 132.600 340.050 132.900 ;
        RECT 346.950 132.600 349.050 133.050 ;
        RECT 337.950 131.400 349.050 132.600 ;
        RECT 337.950 130.800 340.050 131.400 ;
        RECT 346.950 130.950 349.050 131.400 ;
        RECT 385.950 132.450 388.050 132.900 ;
        RECT 397.950 132.450 400.050 132.900 ;
        RECT 385.950 131.250 400.050 132.450 ;
        RECT 385.950 130.800 388.050 131.250 ;
        RECT 397.950 130.800 400.050 131.250 ;
        RECT 409.950 132.450 412.050 132.900 ;
        RECT 418.800 132.450 420.900 132.900 ;
        RECT 409.950 131.250 420.900 132.450 ;
        RECT 409.950 130.800 412.050 131.250 ;
        RECT 418.800 130.800 420.900 131.250 ;
        RECT 421.950 132.450 424.050 132.900 ;
        RECT 430.950 132.600 433.050 132.900 ;
        RECT 445.950 132.600 448.050 133.050 ;
        RECT 430.950 132.450 448.050 132.600 ;
        RECT 421.950 131.400 448.050 132.450 ;
        RECT 421.950 131.250 433.050 131.400 ;
        RECT 421.950 130.800 424.050 131.250 ;
        RECT 430.950 130.800 433.050 131.250 ;
        RECT 445.950 130.950 448.050 131.400 ;
        RECT 454.950 132.600 457.050 132.900 ;
        RECT 470.400 132.600 471.600 137.400 ;
        RECT 472.950 137.100 475.050 137.400 ;
        RECT 478.950 138.600 481.050 139.200 ;
        RECT 511.950 138.600 514.050 139.200 ;
        RECT 478.950 137.400 514.050 138.600 ;
        RECT 478.950 137.100 481.050 137.400 ;
        RECT 511.950 137.100 514.050 137.400 ;
        RECT 532.950 138.750 535.050 139.200 ;
        RECT 550.950 138.750 553.050 139.200 ;
        RECT 532.950 137.550 553.050 138.750 ;
        RECT 532.950 137.100 535.050 137.550 ;
        RECT 550.950 137.100 553.050 137.550 ;
        RECT 592.950 138.600 595.050 139.200 ;
        RECT 598.950 138.600 601.050 139.050 ;
        RECT 592.950 137.400 601.050 138.600 ;
        RECT 592.950 137.100 595.050 137.400 ;
        RECT 598.950 136.950 601.050 137.400 ;
        RECT 622.950 138.750 625.050 139.200 ;
        RECT 637.950 138.750 640.050 139.200 ;
        RECT 622.950 137.550 640.050 138.750 ;
        RECT 622.950 137.100 625.050 137.550 ;
        RECT 637.950 137.100 640.050 137.550 ;
        RECT 661.950 138.750 664.050 139.200 ;
        RECT 670.950 138.750 673.050 139.200 ;
        RECT 661.950 137.550 673.050 138.750 ;
        RECT 661.950 137.100 664.050 137.550 ;
        RECT 670.950 137.100 673.050 137.550 ;
        RECT 676.950 138.600 679.050 139.200 ;
        RECT 709.950 138.600 712.050 139.200 ;
        RECT 676.950 137.400 712.050 138.600 ;
        RECT 676.950 137.100 679.050 137.400 ;
        RECT 709.950 137.100 712.050 137.400 ;
        RECT 721.950 138.750 724.050 139.200 ;
        RECT 730.950 138.750 733.050 139.200 ;
        RECT 721.950 137.550 733.050 138.750 ;
        RECT 721.950 137.100 724.050 137.550 ;
        RECT 730.950 137.100 733.050 137.550 ;
        RECT 808.950 138.750 811.050 139.200 ;
        RECT 820.950 138.750 823.050 139.200 ;
        RECT 808.950 137.550 823.050 138.750 ;
        RECT 808.950 137.100 811.050 137.550 ;
        RECT 820.950 137.100 823.050 137.550 ;
        RECT 838.950 138.600 841.050 139.050 ;
        RECT 871.950 138.600 874.050 139.050 ;
        RECT 838.950 137.400 874.050 138.600 ;
        RECT 838.950 136.950 841.050 137.400 ;
        RECT 871.950 136.950 874.050 137.400 ;
        RECT 922.950 138.750 925.050 139.200 ;
        RECT 940.950 138.750 943.050 139.200 ;
        RECT 922.950 137.550 943.050 138.750 ;
        RECT 922.950 137.100 925.050 137.550 ;
        RECT 940.950 137.100 943.050 137.550 ;
        RECT 994.950 137.100 997.050 139.200 ;
        RECT 941.400 135.600 942.600 137.100 ;
        RECT 946.950 135.600 949.050 136.050 ;
        RECT 941.400 134.400 949.050 135.600 ;
        RECT 946.950 133.950 949.050 134.400 ;
        RECT 454.950 131.400 471.600 132.600 ;
        RECT 520.950 132.450 523.050 132.900 ;
        RECT 529.950 132.450 532.050 132.900 ;
        RECT 454.950 130.800 457.050 131.400 ;
        RECT 520.950 131.250 532.050 132.450 ;
        RECT 520.950 130.800 523.050 131.250 ;
        RECT 529.950 130.800 532.050 131.250 ;
        RECT 571.950 132.450 574.050 132.900 ;
        RECT 577.950 132.450 580.050 132.900 ;
        RECT 571.950 131.250 580.050 132.450 ;
        RECT 571.950 130.800 574.050 131.250 ;
        RECT 577.950 130.800 580.050 131.250 ;
        RECT 634.950 132.450 637.050 132.900 ;
        RECT 652.950 132.450 655.050 132.900 ;
        RECT 634.950 131.250 655.050 132.450 ;
        RECT 634.950 130.800 637.050 131.250 ;
        RECT 652.950 130.800 655.050 131.250 ;
        RECT 682.950 132.450 685.050 132.900 ;
        RECT 694.950 132.450 697.050 132.900 ;
        RECT 682.950 131.250 697.050 132.450 ;
        RECT 682.950 130.800 685.050 131.250 ;
        RECT 694.950 130.800 697.050 131.250 ;
        RECT 715.950 132.450 718.050 132.900 ;
        RECT 727.950 132.450 730.050 132.900 ;
        RECT 715.950 131.250 730.050 132.450 ;
        RECT 715.950 130.800 718.050 131.250 ;
        RECT 727.950 130.800 730.050 131.250 ;
        RECT 811.950 132.600 814.050 133.050 ;
        RECT 823.950 132.600 826.050 132.900 ;
        RECT 811.950 131.400 826.050 132.600 ;
        RECT 811.950 130.950 814.050 131.400 ;
        RECT 823.950 130.800 826.050 131.400 ;
        RECT 865.950 132.600 868.050 133.050 ;
        RECT 883.950 132.600 886.050 132.900 ;
        RECT 865.950 131.400 886.050 132.600 ;
        RECT 865.950 130.950 868.050 131.400 ;
        RECT 883.950 130.800 886.050 131.400 ;
        RECT 916.950 132.450 919.050 132.900 ;
        RECT 925.950 132.600 928.050 132.900 ;
        RECT 925.950 132.450 939.600 132.600 ;
        RECT 916.950 131.400 939.600 132.450 ;
        RECT 916.950 131.250 928.050 131.400 ;
        RECT 916.950 130.800 919.050 131.250 ;
        RECT 925.950 130.800 928.050 131.250 ;
        RECT 938.400 130.050 939.600 131.400 ;
        RECT 952.950 132.450 955.050 132.900 ;
        RECT 958.950 132.450 961.050 132.900 ;
        RECT 952.950 131.250 961.050 132.450 ;
        RECT 952.950 130.800 955.050 131.250 ;
        RECT 958.950 130.800 961.050 131.250 ;
        RECT 1000.950 132.600 1003.050 133.050 ;
        RECT 1015.950 132.600 1018.050 132.900 ;
        RECT 1000.950 131.400 1018.050 132.600 ;
        RECT 1000.950 130.950 1003.050 131.400 ;
        RECT 1015.950 130.800 1018.050 131.400 ;
        RECT 127.950 129.600 130.050 130.050 ;
        RECT 139.950 129.600 142.050 130.050 ;
        RECT 127.950 128.400 142.050 129.600 ;
        RECT 127.950 127.950 130.050 128.400 ;
        RECT 139.950 127.950 142.050 128.400 ;
        RECT 307.950 129.600 310.050 130.050 ;
        RECT 331.950 129.600 334.050 130.050 ;
        RECT 307.950 128.400 334.050 129.600 ;
        RECT 307.950 127.950 310.050 128.400 ;
        RECT 331.950 127.950 334.050 128.400 ;
        RECT 448.950 129.600 451.050 130.050 ;
        RECT 454.950 129.600 457.050 130.050 ;
        RECT 448.950 128.400 457.050 129.600 ;
        RECT 448.950 127.950 451.050 128.400 ;
        RECT 454.950 127.950 457.050 128.400 ;
        RECT 460.950 129.600 463.050 130.050 ;
        RECT 469.950 129.600 472.050 130.050 ;
        RECT 460.950 128.400 472.050 129.600 ;
        RECT 460.950 127.950 463.050 128.400 ;
        RECT 469.950 127.950 472.050 128.400 ;
        RECT 505.950 129.600 508.050 130.050 ;
        RECT 517.950 129.600 520.050 130.050 ;
        RECT 505.950 128.400 520.050 129.600 ;
        RECT 505.950 127.950 508.050 128.400 ;
        RECT 517.950 127.950 520.050 128.400 ;
        RECT 616.950 129.600 619.050 130.050 ;
        RECT 628.950 129.600 631.050 130.050 ;
        RECT 616.950 128.400 631.050 129.600 ;
        RECT 616.950 127.950 619.050 128.400 ;
        RECT 628.950 127.950 631.050 128.400 ;
        RECT 664.950 129.600 667.050 130.050 ;
        RECT 676.950 129.600 679.050 130.050 ;
        RECT 664.950 128.400 679.050 129.600 ;
        RECT 664.950 127.950 667.050 128.400 ;
        RECT 676.950 127.950 679.050 128.400 ;
        RECT 796.950 129.600 799.050 130.050 ;
        RECT 808.950 129.600 811.050 130.050 ;
        RECT 796.950 128.400 811.050 129.600 ;
        RECT 938.400 128.400 943.050 130.050 ;
        RECT 796.950 127.950 799.050 128.400 ;
        RECT 808.950 127.950 811.050 128.400 ;
        RECT 939.000 127.950 943.050 128.400 ;
        RECT 91.950 126.600 94.050 127.050 ;
        RECT 100.950 126.600 103.050 127.050 ;
        RECT 91.950 125.400 103.050 126.600 ;
        RECT 91.950 124.950 94.050 125.400 ;
        RECT 100.950 124.950 103.050 125.400 ;
        RECT 118.950 126.600 121.050 127.050 ;
        RECT 154.950 126.600 157.050 127.050 ;
        RECT 118.950 125.400 157.050 126.600 ;
        RECT 118.950 124.950 121.050 125.400 ;
        RECT 154.950 124.950 157.050 125.400 ;
        RECT 166.950 126.600 169.050 127.050 ;
        RECT 217.950 126.600 220.050 127.050 ;
        RECT 166.950 125.400 220.050 126.600 ;
        RECT 166.950 124.950 169.050 125.400 ;
        RECT 217.950 124.950 220.050 125.400 ;
        RECT 244.950 126.600 247.050 127.050 ;
        RECT 259.950 126.600 262.050 127.050 ;
        RECT 244.950 125.400 262.050 126.600 ;
        RECT 244.950 124.950 247.050 125.400 ;
        RECT 259.950 124.950 262.050 125.400 ;
        RECT 268.950 126.600 271.050 127.050 ;
        RECT 283.950 126.600 286.050 127.050 ;
        RECT 301.950 126.600 304.050 127.050 ;
        RECT 268.950 125.400 304.050 126.600 ;
        RECT 268.950 124.950 271.050 125.400 ;
        RECT 283.950 124.950 286.050 125.400 ;
        RECT 301.950 124.950 304.050 125.400 ;
        RECT 349.950 126.600 352.050 127.050 ;
        RECT 358.950 126.600 361.050 127.050 ;
        RECT 349.950 125.400 361.050 126.600 ;
        RECT 349.950 124.950 352.050 125.400 ;
        RECT 358.950 124.950 361.050 125.400 ;
        RECT 490.950 126.600 493.050 127.050 ;
        RECT 592.950 126.600 595.050 127.050 ;
        RECT 490.950 125.400 595.050 126.600 ;
        RECT 490.950 124.950 493.050 125.400 ;
        RECT 592.950 124.950 595.050 125.400 ;
        RECT 691.950 126.600 694.050 127.050 ;
        RECT 700.950 126.600 703.050 127.050 ;
        RECT 720.000 126.600 724.050 127.050 ;
        RECT 691.950 125.400 703.050 126.600 ;
        RECT 691.950 124.950 694.050 125.400 ;
        RECT 700.950 124.950 703.050 125.400 ;
        RECT 719.400 124.950 724.050 126.600 ;
        RECT 811.950 126.600 814.050 127.050 ;
        RECT 853.950 126.600 856.050 127.050 ;
        RECT 811.950 125.400 856.050 126.600 ;
        RECT 811.950 124.950 814.050 125.400 ;
        RECT 853.950 124.950 856.050 125.400 ;
        RECT 871.950 126.600 874.050 127.050 ;
        RECT 904.950 126.600 907.050 127.050 ;
        RECT 871.950 125.400 907.050 126.600 ;
        RECT 871.950 124.950 874.050 125.400 ;
        RECT 904.950 124.950 907.050 125.400 ;
        RECT 1021.950 126.600 1024.050 127.050 ;
        RECT 1030.950 126.600 1033.050 127.050 ;
        RECT 1021.950 125.400 1033.050 126.600 ;
        RECT 1021.950 124.950 1024.050 125.400 ;
        RECT 1030.950 124.950 1033.050 125.400 ;
        RECT 218.400 123.600 219.600 124.950 ;
        RECT 256.950 123.600 259.050 124.050 ;
        RECT 218.400 122.400 259.050 123.600 ;
        RECT 256.950 121.950 259.050 122.400 ;
        RECT 262.950 123.600 265.050 124.050 ;
        RECT 313.950 123.600 316.050 124.050 ;
        RECT 325.950 123.600 328.050 124.050 ;
        RECT 262.950 122.400 328.050 123.600 ;
        RECT 262.950 121.950 265.050 122.400 ;
        RECT 313.950 121.950 316.050 122.400 ;
        RECT 325.950 121.950 328.050 122.400 ;
        RECT 376.950 123.600 379.050 124.050 ;
        RECT 403.950 123.600 406.050 124.050 ;
        RECT 376.950 122.400 406.050 123.600 ;
        RECT 376.950 121.950 379.050 122.400 ;
        RECT 403.950 121.950 406.050 122.400 ;
        RECT 514.950 123.600 517.050 124.050 ;
        RECT 535.950 123.600 538.050 124.050 ;
        RECT 514.950 122.400 538.050 123.600 ;
        RECT 514.950 121.950 517.050 122.400 ;
        RECT 535.950 121.950 538.050 122.400 ;
        RECT 565.950 123.600 568.050 124.050 ;
        RECT 661.950 123.600 664.050 124.050 ;
        RECT 682.950 123.600 685.050 124.050 ;
        RECT 565.950 122.400 685.050 123.600 ;
        RECT 565.950 121.950 568.050 122.400 ;
        RECT 661.950 121.950 664.050 122.400 ;
        RECT 682.950 121.950 685.050 122.400 ;
        RECT 706.950 123.600 709.050 124.050 ;
        RECT 719.400 123.600 720.600 124.950 ;
        RECT 706.950 122.400 720.600 123.600 ;
        RECT 727.950 123.600 730.050 124.050 ;
        RECT 751.950 123.600 754.050 124.050 ;
        RECT 727.950 122.400 754.050 123.600 ;
        RECT 706.950 121.950 709.050 122.400 ;
        RECT 727.950 121.950 730.050 122.400 ;
        RECT 751.950 121.950 754.050 122.400 ;
        RECT 784.950 123.600 787.050 124.050 ;
        RECT 865.950 123.600 868.050 124.050 ;
        RECT 784.950 122.400 868.050 123.600 ;
        RECT 784.950 121.950 787.050 122.400 ;
        RECT 865.950 121.950 868.050 122.400 ;
        RECT 22.950 120.600 25.050 121.050 ;
        RECT 67.950 120.600 70.050 121.050 ;
        RECT 22.950 119.400 70.050 120.600 ;
        RECT 22.950 118.950 25.050 119.400 ;
        RECT 67.950 118.950 70.050 119.400 ;
        RECT 79.950 120.600 82.050 121.050 ;
        RECT 145.950 120.600 148.050 121.050 ;
        RECT 277.950 120.600 280.050 121.050 ;
        RECT 307.950 120.600 310.050 121.050 ;
        RECT 79.950 119.400 310.050 120.600 ;
        RECT 79.950 118.950 82.050 119.400 ;
        RECT 145.950 118.950 148.050 119.400 ;
        RECT 277.950 118.950 280.050 119.400 ;
        RECT 307.950 118.950 310.050 119.400 ;
        RECT 406.950 120.600 409.050 121.050 ;
        RECT 508.950 120.600 511.050 121.050 ;
        RECT 406.950 119.400 511.050 120.600 ;
        RECT 406.950 118.950 409.050 119.400 ;
        RECT 508.950 118.950 511.050 119.400 ;
        RECT 721.950 120.600 724.050 121.050 ;
        RECT 778.950 120.600 781.050 121.050 ;
        RECT 721.950 119.400 781.050 120.600 ;
        RECT 721.950 118.950 724.050 119.400 ;
        RECT 778.950 118.950 781.050 119.400 ;
        RECT 799.950 120.600 802.050 121.050 ;
        RECT 829.950 120.600 832.050 121.050 ;
        RECT 844.950 120.600 847.050 121.050 ;
        RECT 799.950 119.400 847.050 120.600 ;
        RECT 799.950 118.950 802.050 119.400 ;
        RECT 829.950 118.950 832.050 119.400 ;
        RECT 844.950 118.950 847.050 119.400 ;
        RECT 919.950 120.600 922.050 121.050 ;
        RECT 925.950 120.600 928.050 121.050 ;
        RECT 919.950 119.400 928.050 120.600 ;
        RECT 919.950 118.950 922.050 119.400 ;
        RECT 925.950 118.950 928.050 119.400 ;
        RECT 157.950 117.600 160.050 118.050 ;
        RECT 169.950 117.600 172.050 118.050 ;
        RECT 157.950 116.400 172.050 117.600 ;
        RECT 157.950 115.950 160.050 116.400 ;
        RECT 169.950 115.950 172.050 116.400 ;
        RECT 196.950 117.600 199.050 118.050 ;
        RECT 214.950 117.600 217.050 118.050 ;
        RECT 268.950 117.600 271.050 118.050 ;
        RECT 196.950 116.400 271.050 117.600 ;
        RECT 196.950 115.950 199.050 116.400 ;
        RECT 214.950 115.950 217.050 116.400 ;
        RECT 268.950 115.950 271.050 116.400 ;
        RECT 274.950 117.600 277.050 118.050 ;
        RECT 292.950 117.600 295.050 118.050 ;
        RECT 298.950 117.600 301.050 118.050 ;
        RECT 274.950 116.400 301.050 117.600 ;
        RECT 274.950 115.950 277.050 116.400 ;
        RECT 292.950 115.950 295.050 116.400 ;
        RECT 298.950 115.950 301.050 116.400 ;
        RECT 310.950 117.600 313.050 118.050 ;
        RECT 319.950 117.600 322.050 118.050 ;
        RECT 310.950 116.400 322.050 117.600 ;
        RECT 310.950 115.950 313.050 116.400 ;
        RECT 319.950 115.950 322.050 116.400 ;
        RECT 331.950 117.600 334.050 118.050 ;
        RECT 409.950 117.600 412.050 118.050 ;
        RECT 478.950 117.600 481.050 118.050 ;
        RECT 331.950 116.400 481.050 117.600 ;
        RECT 331.950 115.950 334.050 116.400 ;
        RECT 409.950 115.950 412.050 116.400 ;
        RECT 478.950 115.950 481.050 116.400 ;
        RECT 577.950 117.600 580.050 118.050 ;
        RECT 634.950 117.600 637.050 118.050 ;
        RECT 664.950 117.600 667.050 118.050 ;
        RECT 577.950 116.400 637.050 117.600 ;
        RECT 577.950 115.950 580.050 116.400 ;
        RECT 634.950 115.950 637.050 116.400 ;
        RECT 644.400 116.400 667.050 117.600 ;
        RECT 13.950 114.600 16.050 115.050 ;
        RECT 34.950 114.600 37.050 115.050 ;
        RECT 13.950 113.400 37.050 114.600 ;
        RECT 13.950 112.950 16.050 113.400 ;
        RECT 34.950 112.950 37.050 113.400 ;
        RECT 571.950 114.600 574.050 115.050 ;
        RECT 644.400 114.600 645.600 116.400 ;
        RECT 664.950 115.950 667.050 116.400 ;
        RECT 676.950 117.600 679.050 118.050 ;
        RECT 694.950 117.600 697.050 118.050 ;
        RECT 676.950 116.400 697.050 117.600 ;
        RECT 676.950 115.950 679.050 116.400 ;
        RECT 694.950 115.950 697.050 116.400 ;
        RECT 733.950 117.600 736.050 118.050 ;
        RECT 763.950 117.600 766.050 118.050 ;
        RECT 733.950 116.400 766.050 117.600 ;
        RECT 733.950 115.950 736.050 116.400 ;
        RECT 763.950 115.950 766.050 116.400 ;
        RECT 784.950 117.600 787.050 118.050 ;
        RECT 823.950 117.600 826.050 118.050 ;
        RECT 784.950 116.400 826.050 117.600 ;
        RECT 784.950 115.950 787.050 116.400 ;
        RECT 823.950 115.950 826.050 116.400 ;
        RECT 571.950 113.400 645.600 114.600 ;
        RECT 646.950 114.600 649.050 115.050 ;
        RECT 658.950 114.600 661.050 115.050 ;
        RECT 646.950 113.400 661.050 114.600 ;
        RECT 571.950 112.950 574.050 113.400 ;
        RECT 646.950 112.950 649.050 113.400 ;
        RECT 658.950 112.950 661.050 113.400 ;
        RECT 94.950 111.600 97.050 112.050 ;
        RECT 109.950 111.600 112.050 112.050 ;
        RECT 94.950 110.400 112.050 111.600 ;
        RECT 94.950 109.950 97.050 110.400 ;
        RECT 109.950 109.950 112.050 110.400 ;
        RECT 124.950 111.600 127.050 112.050 ;
        RECT 145.950 111.600 148.050 112.050 ;
        RECT 124.950 110.400 148.050 111.600 ;
        RECT 124.950 109.950 127.050 110.400 ;
        RECT 145.950 109.950 148.050 110.400 ;
        RECT 256.950 111.600 259.050 112.050 ;
        RECT 265.950 111.600 268.050 112.050 ;
        RECT 256.950 110.400 268.050 111.600 ;
        RECT 256.950 109.950 259.050 110.400 ;
        RECT 265.950 109.950 268.050 110.400 ;
        RECT 349.950 111.600 352.050 112.050 ;
        RECT 385.950 111.600 388.050 112.050 ;
        RECT 349.950 110.400 388.050 111.600 ;
        RECT 349.950 109.950 352.050 110.400 ;
        RECT 385.950 109.950 388.050 110.400 ;
        RECT 430.950 111.600 433.050 112.050 ;
        RECT 439.950 111.600 442.050 112.050 ;
        RECT 430.950 110.400 442.050 111.600 ;
        RECT 430.950 109.950 433.050 110.400 ;
        RECT 439.950 109.950 442.050 110.400 ;
        RECT 457.950 111.600 460.050 112.050 ;
        RECT 514.950 111.600 517.050 112.050 ;
        RECT 538.950 111.600 541.050 112.050 ;
        RECT 457.950 110.400 541.050 111.600 ;
        RECT 457.950 109.950 460.050 110.400 ;
        RECT 514.950 109.950 517.050 110.400 ;
        RECT 538.950 109.950 541.050 110.400 ;
        RECT 574.950 111.600 577.050 112.050 ;
        RECT 610.950 111.600 613.050 112.050 ;
        RECT 574.950 110.400 613.050 111.600 ;
        RECT 574.950 109.950 577.050 110.400 ;
        RECT 610.950 109.950 613.050 110.400 ;
        RECT 625.950 111.600 628.050 112.050 ;
        RECT 631.950 111.600 634.050 112.050 ;
        RECT 646.950 111.600 649.050 111.900 ;
        RECT 625.950 110.400 649.050 111.600 ;
        RECT 625.950 109.950 628.050 110.400 ;
        RECT 631.950 109.950 634.050 110.400 ;
        RECT 646.950 109.800 649.050 110.400 ;
        RECT 679.950 111.600 682.050 112.050 ;
        RECT 691.950 111.600 694.050 112.050 ;
        RECT 811.950 111.600 814.050 112.050 ;
        RECT 679.950 110.400 814.050 111.600 ;
        RECT 679.950 109.950 682.050 110.400 ;
        RECT 691.950 109.950 694.050 110.400 ;
        RECT 811.950 109.950 814.050 110.400 ;
        RECT 850.950 111.600 853.050 112.050 ;
        RECT 874.950 111.600 877.050 112.050 ;
        RECT 850.950 110.400 877.050 111.600 ;
        RECT 850.950 109.950 853.050 110.400 ;
        RECT 874.950 109.950 877.050 110.400 ;
        RECT 880.950 111.600 883.050 112.050 ;
        RECT 970.950 111.600 973.050 112.050 ;
        RECT 880.950 110.400 973.050 111.600 ;
        RECT 880.950 109.950 883.050 110.400 ;
        RECT 970.950 109.950 973.050 110.400 ;
        RECT 16.950 108.600 19.050 109.050 ;
        RECT 22.950 108.600 25.050 109.050 ;
        RECT 16.950 107.400 25.050 108.600 ;
        RECT 16.950 106.950 19.050 107.400 ;
        RECT 22.950 106.950 25.050 107.400 ;
        RECT 298.950 108.600 301.050 109.050 ;
        RECT 304.950 108.600 307.050 109.050 ;
        RECT 298.950 107.400 307.050 108.600 ;
        RECT 298.950 106.950 301.050 107.400 ;
        RECT 304.950 106.950 307.050 107.400 ;
        RECT 460.950 108.600 463.050 109.050 ;
        RECT 466.950 108.600 469.050 109.050 ;
        RECT 460.950 107.400 469.050 108.600 ;
        RECT 460.950 106.950 463.050 107.400 ;
        RECT 466.950 106.950 469.050 107.400 ;
        RECT 544.950 108.600 547.050 109.050 ;
        RECT 553.950 108.600 556.050 109.050 ;
        RECT 784.950 108.600 787.050 109.050 ;
        RECT 544.950 107.400 556.050 108.600 ;
        RECT 544.950 106.950 547.050 107.400 ;
        RECT 553.950 106.950 556.050 107.400 ;
        RECT 713.400 107.400 787.050 108.600 ;
        RECT 22.950 105.750 25.050 106.200 ;
        RECT 31.950 105.750 34.050 106.200 ;
        RECT 22.950 104.550 34.050 105.750 ;
        RECT 22.950 104.100 25.050 104.550 ;
        RECT 31.950 104.100 34.050 104.550 ;
        RECT 43.950 105.600 46.050 106.200 ;
        RECT 82.950 105.600 85.050 106.050 ;
        RECT 43.950 104.400 85.050 105.600 ;
        RECT 43.950 104.100 46.050 104.400 ;
        RECT 82.950 103.950 85.050 104.400 ;
        RECT 133.950 105.750 136.050 106.200 ;
        RECT 139.950 105.750 142.050 106.200 ;
        RECT 133.950 104.550 142.050 105.750 ;
        RECT 133.950 104.100 136.050 104.550 ;
        RECT 139.950 104.100 142.050 104.550 ;
        RECT 145.950 105.600 148.050 106.050 ;
        RECT 187.950 105.600 190.050 106.200 ;
        RECT 145.950 104.400 190.050 105.600 ;
        RECT 145.950 103.950 148.050 104.400 ;
        RECT 187.950 104.100 190.050 104.400 ;
        RECT 196.950 105.750 199.050 106.200 ;
        RECT 211.950 105.750 214.050 106.200 ;
        RECT 196.950 104.550 214.050 105.750 ;
        RECT 196.950 104.100 199.050 104.550 ;
        RECT 211.950 104.100 214.050 104.550 ;
        RECT 223.950 105.600 226.050 106.050 ;
        RECT 235.950 105.600 238.050 106.200 ;
        RECT 274.950 105.600 277.050 106.050 ;
        RECT 223.950 104.400 238.050 105.600 ;
        RECT 223.950 103.950 226.050 104.400 ;
        RECT 235.950 104.100 238.050 104.400 ;
        RECT 239.400 104.400 277.050 105.600 ;
        RECT 239.400 99.900 240.600 104.400 ;
        RECT 274.950 103.950 277.050 104.400 ;
        RECT 373.950 105.750 376.050 106.200 ;
        RECT 379.950 105.750 382.050 106.200 ;
        RECT 373.950 104.550 382.050 105.750 ;
        RECT 373.950 104.100 376.050 104.550 ;
        RECT 379.950 104.100 382.050 104.550 ;
        RECT 391.950 105.750 394.050 106.200 ;
        RECT 406.950 105.750 409.050 106.200 ;
        RECT 391.950 104.550 409.050 105.750 ;
        RECT 391.950 104.100 394.050 104.550 ;
        RECT 406.950 104.100 409.050 104.550 ;
        RECT 424.950 105.750 427.050 106.200 ;
        RECT 436.950 105.750 439.050 106.200 ;
        RECT 424.950 104.550 439.050 105.750 ;
        RECT 424.950 104.100 427.050 104.550 ;
        RECT 436.950 104.100 439.050 104.550 ;
        RECT 556.950 105.750 559.050 106.200 ;
        RECT 565.950 105.750 568.050 106.200 ;
        RECT 556.950 104.550 568.050 105.750 ;
        RECT 574.950 105.600 577.050 106.050 ;
        RECT 556.950 104.100 559.050 104.550 ;
        RECT 565.950 104.100 568.050 104.550 ;
        RECT 569.400 104.400 577.050 105.600 ;
        RECT 334.950 102.450 337.050 102.900 ;
        RECT 349.950 102.450 352.050 102.900 ;
        RECT 569.400 102.600 570.600 104.400 ;
        RECT 574.950 103.950 577.050 104.400 ;
        RECT 580.950 105.600 583.050 106.050 ;
        RECT 598.950 105.600 601.050 106.050 ;
        RECT 580.950 104.400 601.050 105.600 ;
        RECT 580.950 103.950 583.050 104.400 ;
        RECT 598.950 103.950 601.050 104.400 ;
        RECT 604.950 105.600 607.050 106.050 ;
        RECT 616.950 105.600 619.050 106.200 ;
        RECT 604.950 104.400 619.050 105.600 ;
        RECT 604.950 103.950 607.050 104.400 ;
        RECT 616.950 104.100 619.050 104.400 ;
        RECT 652.950 105.750 655.050 106.200 ;
        RECT 658.950 105.750 661.050 106.200 ;
        RECT 652.950 104.550 661.050 105.750 ;
        RECT 652.950 104.100 655.050 104.550 ;
        RECT 658.950 104.100 661.050 104.550 ;
        RECT 673.950 105.600 676.050 106.200 ;
        RECT 713.400 106.050 714.600 107.400 ;
        RECT 784.950 106.950 787.050 107.400 ;
        RECT 934.950 108.600 937.050 109.050 ;
        RECT 967.950 108.600 970.050 109.050 ;
        RECT 934.950 107.400 970.050 108.600 ;
        RECT 934.950 106.950 937.050 107.400 ;
        RECT 967.950 106.950 970.050 107.400 ;
        RECT 685.950 105.600 688.050 106.050 ;
        RECT 688.950 105.600 691.050 106.050 ;
        RECT 673.950 104.400 691.050 105.600 ;
        RECT 673.950 104.100 676.050 104.400 ;
        RECT 685.950 103.950 688.050 104.400 ;
        RECT 688.950 103.950 691.050 104.400 ;
        RECT 694.950 105.600 697.050 106.050 ;
        RECT 712.950 105.600 715.050 106.050 ;
        RECT 763.950 105.600 766.050 106.050 ;
        RECT 694.950 104.400 715.050 105.600 ;
        RECT 694.950 103.950 697.050 104.400 ;
        RECT 712.950 103.950 715.050 104.400 ;
        RECT 749.400 104.400 766.050 105.600 ;
        RECT 749.400 102.900 750.600 104.400 ;
        RECT 763.950 103.950 766.050 104.400 ;
        RECT 787.950 105.750 790.050 106.200 ;
        RECT 817.950 105.750 820.050 106.200 ;
        RECT 787.950 104.550 820.050 105.750 ;
        RECT 787.950 104.100 790.050 104.550 ;
        RECT 817.950 104.100 820.050 104.550 ;
        RECT 844.950 105.600 847.050 106.200 ;
        RECT 865.950 105.600 868.050 106.200 ;
        RECT 844.950 104.400 868.050 105.600 ;
        RECT 844.950 104.100 847.050 104.400 ;
        RECT 865.950 104.100 868.050 104.400 ;
        RECT 874.950 105.750 877.050 106.200 ;
        RECT 880.950 105.750 883.050 106.200 ;
        RECT 874.950 104.550 883.050 105.750 ;
        RECT 874.950 104.100 877.050 104.550 ;
        RECT 880.950 104.100 883.050 104.550 ;
        RECT 925.950 105.600 928.050 106.050 ;
        RECT 931.950 105.600 934.050 106.050 ;
        RECT 925.950 104.400 934.050 105.600 ;
        RECT 925.950 103.950 928.050 104.400 ;
        RECT 931.950 103.950 934.050 104.400 ;
        RECT 976.950 105.750 979.050 106.200 ;
        RECT 985.950 105.750 988.050 106.200 ;
        RECT 976.950 104.550 988.050 105.750 ;
        RECT 976.950 104.100 979.050 104.550 ;
        RECT 985.950 104.100 988.050 104.550 ;
        RECT 334.950 101.250 352.050 102.450 ;
        RECT 334.950 100.800 337.050 101.250 ;
        RECT 349.950 100.800 352.050 101.250 ;
        RECT 545.400 101.400 570.600 102.600 ;
        RECT 19.950 99.600 22.050 99.900 ;
        RECT 46.950 99.600 49.050 99.900 ;
        RECT 19.950 98.400 49.050 99.600 ;
        RECT 19.950 97.800 22.050 98.400 ;
        RECT 46.950 97.800 49.050 98.400 ;
        RECT 70.950 99.600 73.050 99.900 ;
        RECT 91.950 99.600 94.050 99.900 ;
        RECT 70.950 98.400 94.050 99.600 ;
        RECT 70.950 97.800 73.050 98.400 ;
        RECT 91.950 97.800 94.050 98.400 ;
        RECT 118.950 99.450 121.050 99.900 ;
        RECT 145.950 99.450 148.050 99.900 ;
        RECT 118.950 98.250 148.050 99.450 ;
        RECT 118.950 97.800 121.050 98.250 ;
        RECT 145.950 97.800 148.050 98.250 ;
        RECT 166.950 99.600 169.050 99.900 ;
        RECT 184.950 99.600 187.050 99.900 ;
        RECT 214.950 99.600 217.050 99.900 ;
        RECT 166.950 99.450 217.050 99.600 ;
        RECT 223.950 99.450 226.050 99.900 ;
        RECT 166.950 98.400 226.050 99.450 ;
        RECT 166.950 97.800 169.050 98.400 ;
        RECT 184.950 97.800 187.050 98.400 ;
        RECT 214.950 98.250 226.050 98.400 ;
        RECT 214.950 97.800 217.050 98.250 ;
        RECT 223.950 97.800 226.050 98.250 ;
        RECT 238.950 97.800 241.050 99.900 ;
        RECT 244.950 99.450 247.050 99.900 ;
        RECT 250.950 99.450 253.050 99.900 ;
        RECT 244.950 98.250 253.050 99.450 ;
        RECT 244.950 97.800 247.050 98.250 ;
        RECT 250.950 97.800 253.050 98.250 ;
        RECT 262.950 99.450 265.050 99.900 ;
        RECT 277.950 99.450 280.050 99.900 ;
        RECT 262.950 98.250 280.050 99.450 ;
        RECT 262.950 97.800 265.050 98.250 ;
        RECT 277.950 97.800 280.050 98.250 ;
        RECT 283.950 99.600 286.050 100.050 ;
        RECT 289.950 99.600 292.050 99.900 ;
        RECT 283.950 98.400 292.050 99.600 ;
        RECT 283.950 97.950 286.050 98.400 ;
        RECT 289.950 97.800 292.050 98.400 ;
        RECT 313.950 99.600 316.050 100.050 ;
        RECT 382.950 99.600 385.050 99.900 ;
        RECT 313.950 99.450 385.050 99.600 ;
        RECT 397.950 99.450 400.050 99.900 ;
        RECT 313.950 98.400 400.050 99.450 ;
        RECT 313.950 97.950 316.050 98.400 ;
        RECT 382.950 98.250 400.050 98.400 ;
        RECT 382.950 97.800 385.050 98.250 ;
        RECT 397.950 97.800 400.050 98.250 ;
        RECT 433.950 99.600 436.050 99.900 ;
        RECT 448.950 99.600 451.050 100.050 ;
        RECT 433.950 98.400 451.050 99.600 ;
        RECT 433.950 97.800 436.050 98.400 ;
        RECT 448.950 97.950 451.050 98.400 ;
        RECT 460.950 99.450 463.050 99.900 ;
        RECT 466.950 99.450 469.050 99.900 ;
        RECT 460.950 98.250 469.050 99.450 ;
        RECT 460.950 97.800 463.050 98.250 ;
        RECT 466.950 97.800 469.050 98.250 ;
        RECT 541.950 99.600 544.050 99.900 ;
        RECT 545.400 99.600 546.600 101.400 ;
        RECT 748.950 100.800 751.050 102.900 ;
        RECT 541.950 98.400 546.600 99.600 ;
        RECT 553.950 99.450 556.050 99.900 ;
        RECT 562.950 99.450 565.050 99.900 ;
        RECT 541.950 97.800 544.050 98.400 ;
        RECT 553.950 98.250 565.050 99.450 ;
        RECT 553.950 97.800 556.050 98.250 ;
        RECT 562.950 97.800 565.050 98.250 ;
        RECT 583.950 99.450 586.050 99.900 ;
        RECT 589.950 99.450 592.050 99.900 ;
        RECT 583.950 98.250 592.050 99.450 ;
        RECT 583.950 97.800 586.050 98.250 ;
        RECT 589.950 97.800 592.050 98.250 ;
        RECT 619.950 99.450 622.050 99.900 ;
        RECT 625.950 99.450 628.050 99.900 ;
        RECT 619.950 98.250 628.050 99.450 ;
        RECT 619.950 97.800 622.050 98.250 ;
        RECT 625.950 97.800 628.050 98.250 ;
        RECT 631.950 99.450 634.050 99.900 ;
        RECT 637.950 99.450 640.050 99.900 ;
        RECT 631.950 98.250 640.050 99.450 ;
        RECT 631.950 97.800 634.050 98.250 ;
        RECT 637.950 97.800 640.050 98.250 ;
        RECT 664.950 99.450 667.050 99.900 ;
        RECT 676.950 99.450 679.050 99.900 ;
        RECT 664.950 98.250 679.050 99.450 ;
        RECT 664.950 97.800 667.050 98.250 ;
        RECT 676.950 97.800 679.050 98.250 ;
        RECT 691.950 99.450 694.050 99.900 ;
        RECT 697.950 99.450 700.050 99.900 ;
        RECT 691.950 98.250 700.050 99.450 ;
        RECT 691.950 97.800 694.050 98.250 ;
        RECT 697.950 97.800 700.050 98.250 ;
        RECT 784.950 99.450 787.050 99.900 ;
        RECT 799.950 99.450 802.050 99.900 ;
        RECT 784.950 98.250 802.050 99.450 ;
        RECT 784.950 97.800 787.050 98.250 ;
        RECT 799.950 97.800 802.050 98.250 ;
        RECT 820.950 99.600 823.050 99.900 ;
        RECT 835.950 99.600 838.050 100.050 ;
        RECT 820.950 98.400 838.050 99.600 ;
        RECT 820.950 97.800 823.050 98.400 ;
        RECT 835.950 97.950 838.050 98.400 ;
        RECT 904.950 99.600 907.050 100.050 ;
        RECT 928.950 99.600 931.050 103.050 ;
        RECT 904.950 99.000 931.050 99.600 ;
        RECT 904.950 98.400 930.600 99.000 ;
        RECT 904.950 97.950 907.050 98.400 ;
        RECT 190.950 96.600 193.050 97.050 ;
        RECT 196.950 96.600 199.050 97.050 ;
        RECT 190.950 95.400 199.050 96.600 ;
        RECT 190.950 94.950 193.050 95.400 ;
        RECT 196.950 94.950 199.050 95.400 ;
        RECT 358.950 96.450 361.050 96.900 ;
        RECT 370.950 96.450 373.050 96.900 ;
        RECT 358.950 95.250 373.050 96.450 ;
        RECT 358.950 94.800 361.050 95.250 ;
        RECT 370.950 94.800 373.050 95.250 ;
        RECT 391.950 96.600 394.050 97.050 ;
        RECT 424.950 96.600 427.050 97.050 ;
        RECT 391.950 95.400 427.050 96.600 ;
        RECT 391.950 94.950 394.050 95.400 ;
        RECT 424.950 94.950 427.050 95.400 ;
        RECT 850.950 96.450 853.050 96.900 ;
        RECT 880.950 96.450 883.050 96.900 ;
        RECT 850.950 95.250 883.050 96.450 ;
        RECT 850.950 94.800 853.050 95.250 ;
        RECT 880.950 94.800 883.050 95.250 ;
        RECT 985.950 96.600 988.050 97.050 ;
        RECT 1000.950 96.600 1003.050 97.050 ;
        RECT 985.950 95.400 1003.050 96.600 ;
        RECT 985.950 94.950 988.050 95.400 ;
        RECT 1000.950 94.950 1003.050 95.400 ;
        RECT 28.950 93.600 31.050 94.050 ;
        RECT 145.950 93.600 148.050 94.050 ;
        RECT 28.950 92.400 148.050 93.600 ;
        RECT 28.950 91.950 31.050 92.400 ;
        RECT 145.950 91.950 148.050 92.400 ;
        RECT 487.950 93.600 490.050 94.050 ;
        RECT 604.950 93.600 607.050 94.050 ;
        RECT 487.950 92.400 607.050 93.600 ;
        RECT 487.950 91.950 490.050 92.400 ;
        RECT 604.950 91.950 607.050 92.400 ;
        RECT 772.950 93.600 775.050 94.050 ;
        RECT 851.400 93.600 852.600 94.800 ;
        RECT 772.950 92.400 852.600 93.600 ;
        RECT 925.950 93.600 928.050 94.050 ;
        RECT 940.950 93.600 943.050 94.050 ;
        RECT 925.950 92.400 943.050 93.600 ;
        RECT 772.950 91.950 775.050 92.400 ;
        RECT 925.950 91.950 928.050 92.400 ;
        RECT 940.950 91.950 943.050 92.400 ;
        RECT 1006.950 93.600 1009.050 94.050 ;
        RECT 1021.950 93.600 1024.050 94.050 ;
        RECT 1006.950 92.400 1024.050 93.600 ;
        RECT 1006.950 91.950 1009.050 92.400 ;
        RECT 1021.950 91.950 1024.050 92.400 ;
        RECT 517.950 90.600 520.050 91.050 ;
        RECT 583.950 90.600 586.050 91.050 ;
        RECT 517.950 89.400 586.050 90.600 ;
        RECT 517.950 88.950 520.050 89.400 ;
        RECT 583.950 88.950 586.050 89.400 ;
        RECT 862.950 90.600 865.050 91.050 ;
        RECT 946.950 90.600 949.050 91.050 ;
        RECT 862.950 89.400 949.050 90.600 ;
        RECT 862.950 88.950 865.050 89.400 ;
        RECT 946.950 88.950 949.050 89.400 ;
        RECT 424.950 87.600 427.050 88.050 ;
        RECT 547.950 87.600 550.050 88.050 ;
        RECT 616.950 87.600 619.050 88.050 ;
        RECT 703.950 87.600 706.050 88.050 ;
        RECT 424.950 86.400 706.050 87.600 ;
        RECT 424.950 85.950 427.050 86.400 ;
        RECT 547.950 85.950 550.050 86.400 ;
        RECT 616.950 85.950 619.050 86.400 ;
        RECT 703.950 85.950 706.050 86.400 ;
        RECT 367.950 84.600 370.050 85.050 ;
        RECT 376.950 84.600 379.050 85.050 ;
        RECT 367.950 83.400 379.050 84.600 ;
        RECT 367.950 82.950 370.050 83.400 ;
        RECT 376.950 82.950 379.050 83.400 ;
        RECT 388.950 84.600 391.050 85.050 ;
        RECT 487.950 84.600 490.050 85.050 ;
        RECT 388.950 83.400 490.050 84.600 ;
        RECT 388.950 82.950 391.050 83.400 ;
        RECT 487.950 82.950 490.050 83.400 ;
        RECT 532.950 84.600 535.050 85.050 ;
        RECT 556.950 84.600 559.050 85.050 ;
        RECT 532.950 83.400 559.050 84.600 ;
        RECT 532.950 82.950 535.050 83.400 ;
        RECT 556.950 82.950 559.050 83.400 ;
        RECT 595.950 84.600 598.050 85.050 ;
        RECT 673.950 84.600 676.050 85.050 ;
        RECT 595.950 83.400 676.050 84.600 ;
        RECT 595.950 82.950 598.050 83.400 ;
        RECT 673.950 82.950 676.050 83.400 ;
        RECT 16.950 81.600 19.050 82.050 ;
        RECT 34.950 81.600 37.050 82.050 ;
        RECT 16.950 80.400 37.050 81.600 ;
        RECT 16.950 79.950 19.050 80.400 ;
        RECT 34.950 79.950 37.050 80.400 ;
        RECT 199.950 81.600 202.050 82.050 ;
        RECT 223.950 81.600 226.050 82.050 ;
        RECT 199.950 80.400 226.050 81.600 ;
        RECT 199.950 79.950 202.050 80.400 ;
        RECT 223.950 79.950 226.050 80.400 ;
        RECT 250.950 81.600 253.050 82.050 ;
        RECT 304.950 81.600 307.050 82.050 ;
        RECT 340.950 81.600 343.050 82.050 ;
        RECT 355.950 81.600 358.050 82.050 ;
        RECT 250.950 80.400 358.050 81.600 ;
        RECT 250.950 79.950 253.050 80.400 ;
        RECT 304.950 79.950 307.050 80.400 ;
        RECT 340.950 79.950 343.050 80.400 ;
        RECT 355.950 79.950 358.050 80.400 ;
        RECT 544.950 81.600 547.050 82.050 ;
        RECT 580.950 81.600 583.050 82.050 ;
        RECT 544.950 80.400 583.050 81.600 ;
        RECT 544.950 79.950 547.050 80.400 ;
        RECT 580.950 79.950 583.050 80.400 ;
        RECT 787.950 81.600 790.050 82.050 ;
        RECT 793.950 81.600 796.050 82.050 ;
        RECT 787.950 80.400 796.050 81.600 ;
        RECT 787.950 79.950 790.050 80.400 ;
        RECT 793.950 79.950 796.050 80.400 ;
        RECT 916.950 81.600 919.050 82.050 ;
        RECT 958.950 81.600 961.050 82.050 ;
        RECT 916.950 80.400 961.050 81.600 ;
        RECT 916.950 79.950 919.050 80.400 ;
        RECT 958.950 79.950 961.050 80.400 ;
        RECT 985.950 81.600 988.050 82.050 ;
        RECT 1003.950 81.600 1006.050 82.050 ;
        RECT 1018.950 81.600 1021.050 82.050 ;
        RECT 985.950 80.400 1021.050 81.600 ;
        RECT 985.950 79.950 988.050 80.400 ;
        RECT 1003.950 79.950 1006.050 80.400 ;
        RECT 1018.950 79.950 1021.050 80.400 ;
        RECT 229.950 78.600 232.050 79.050 ;
        RECT 373.950 78.600 376.050 79.050 ;
        RECT 385.950 78.600 388.050 79.050 ;
        RECT 229.950 77.400 388.050 78.600 ;
        RECT 229.950 76.950 232.050 77.400 ;
        RECT 373.950 76.950 376.050 77.400 ;
        RECT 385.950 76.950 388.050 77.400 ;
        RECT 412.950 78.600 415.050 79.050 ;
        RECT 523.950 78.600 526.050 79.050 ;
        RECT 412.950 77.400 526.050 78.600 ;
        RECT 412.950 76.950 415.050 77.400 ;
        RECT 523.950 76.950 526.050 77.400 ;
        RECT 841.950 78.600 844.050 79.050 ;
        RECT 904.950 78.600 907.050 79.050 ;
        RECT 943.950 78.600 946.050 79.050 ;
        RECT 841.950 77.400 946.050 78.600 ;
        RECT 841.950 76.950 844.050 77.400 ;
        RECT 904.950 76.950 907.050 77.400 ;
        RECT 943.950 76.950 946.050 77.400 ;
        RECT 40.950 75.600 43.050 76.050 ;
        RECT 67.950 75.600 70.050 76.050 ;
        RECT 148.950 75.600 151.050 76.050 ;
        RECT 40.950 74.400 151.050 75.600 ;
        RECT 40.950 73.950 43.050 74.400 ;
        RECT 67.950 73.950 70.050 74.400 ;
        RECT 148.950 73.950 151.050 74.400 ;
        RECT 199.950 75.600 202.050 76.050 ;
        RECT 274.950 75.600 277.050 76.050 ;
        RECT 199.950 74.400 277.050 75.600 ;
        RECT 199.950 73.950 202.050 74.400 ;
        RECT 274.950 73.950 277.050 74.400 ;
        RECT 379.950 75.600 382.050 76.050 ;
        RECT 413.400 75.600 414.600 76.950 ;
        RECT 379.950 74.400 414.600 75.600 ;
        RECT 439.950 75.600 442.050 76.050 ;
        RECT 460.950 75.600 463.050 76.050 ;
        RECT 490.950 75.600 493.050 76.050 ;
        RECT 439.950 74.400 493.050 75.600 ;
        RECT 524.400 75.600 525.600 76.950 ;
        RECT 751.950 75.600 754.050 76.050 ;
        RECT 524.400 74.400 754.050 75.600 ;
        RECT 379.950 73.950 382.050 74.400 ;
        RECT 439.950 73.950 442.050 74.400 ;
        RECT 460.950 73.950 463.050 74.400 ;
        RECT 490.950 73.950 493.050 74.400 ;
        RECT 751.950 73.950 754.050 74.400 ;
        RECT 865.950 75.600 868.050 76.050 ;
        RECT 871.950 75.600 874.050 76.050 ;
        RECT 865.950 74.400 874.050 75.600 ;
        RECT 865.950 73.950 868.050 74.400 ;
        RECT 871.950 73.950 874.050 74.400 ;
        RECT 949.950 75.600 952.050 76.050 ;
        RECT 970.950 75.600 973.050 76.050 ;
        RECT 949.950 74.400 973.050 75.600 ;
        RECT 949.950 73.950 952.050 74.400 ;
        RECT 970.950 73.950 973.050 74.400 ;
        RECT 22.950 72.600 25.050 73.050 ;
        RECT 31.950 72.600 34.050 73.050 ;
        RECT 370.950 72.600 373.050 73.050 ;
        RECT 22.950 71.400 373.050 72.600 ;
        RECT 22.950 70.950 25.050 71.400 ;
        RECT 31.950 70.950 34.050 71.400 ;
        RECT 370.950 70.950 373.050 71.400 ;
        RECT 397.950 72.600 400.050 73.050 ;
        RECT 481.950 72.600 484.050 73.050 ;
        RECT 397.950 71.400 484.050 72.600 ;
        RECT 397.950 70.950 400.050 71.400 ;
        RECT 481.950 70.950 484.050 71.400 ;
        RECT 505.950 72.600 508.050 73.050 ;
        RECT 568.950 72.600 571.050 73.050 ;
        RECT 505.950 71.400 571.050 72.600 ;
        RECT 505.950 70.950 508.050 71.400 ;
        RECT 568.950 70.950 571.050 71.400 ;
        RECT 934.950 72.600 937.050 73.050 ;
        RECT 1018.950 72.600 1021.050 73.050 ;
        RECT 934.950 71.400 1021.050 72.600 ;
        RECT 934.950 70.950 937.050 71.400 ;
        RECT 1018.950 70.950 1021.050 71.400 ;
        RECT 115.950 69.600 118.050 70.050 ;
        RECT 136.950 69.600 139.050 70.050 ;
        RECT 142.950 69.600 145.050 70.050 ;
        RECT 115.950 68.400 145.050 69.600 ;
        RECT 115.950 67.950 118.050 68.400 ;
        RECT 136.950 67.950 139.050 68.400 ;
        RECT 142.950 67.950 145.050 68.400 ;
        RECT 148.950 69.600 151.050 70.050 ;
        RECT 181.950 69.600 184.050 70.050 ;
        RECT 202.950 69.600 205.050 70.050 ;
        RECT 229.950 69.600 232.050 70.050 ;
        RECT 607.950 69.600 610.050 70.050 ;
        RECT 148.950 68.400 232.050 69.600 ;
        RECT 148.950 67.950 151.050 68.400 ;
        RECT 181.950 67.950 184.050 68.400 ;
        RECT 202.950 67.950 205.050 68.400 ;
        RECT 229.950 67.950 232.050 68.400 ;
        RECT 305.400 68.400 610.050 69.600 ;
        RECT 305.400 67.050 306.600 68.400 ;
        RECT 607.950 67.950 610.050 68.400 ;
        RECT 655.950 69.600 658.050 70.050 ;
        RECT 730.950 69.600 733.050 70.050 ;
        RECT 655.950 68.400 733.050 69.600 ;
        RECT 655.950 67.950 658.050 68.400 ;
        RECT 730.950 67.950 733.050 68.400 ;
        RECT 139.950 66.600 142.050 67.050 ;
        RECT 256.950 66.600 259.050 67.050 ;
        RECT 304.800 66.600 306.900 67.050 ;
        RECT 139.950 65.400 306.900 66.600 ;
        RECT 139.950 64.950 142.050 65.400 ;
        RECT 256.950 64.950 259.050 65.400 ;
        RECT 304.800 64.950 306.900 65.400 ;
        RECT 307.950 66.600 310.050 67.050 ;
        RECT 319.950 66.600 322.050 67.050 ;
        RECT 388.950 66.600 391.050 67.050 ;
        RECT 307.950 65.400 391.050 66.600 ;
        RECT 307.950 64.950 310.050 65.400 ;
        RECT 319.950 64.950 322.050 65.400 ;
        RECT 388.950 64.950 391.050 65.400 ;
        RECT 424.950 66.600 427.050 67.050 ;
        RECT 493.950 66.600 496.050 67.050 ;
        RECT 424.950 65.400 496.050 66.600 ;
        RECT 424.950 64.950 427.050 65.400 ;
        RECT 493.950 64.950 496.050 65.400 ;
        RECT 514.950 66.600 517.050 67.050 ;
        RECT 577.950 66.600 580.050 67.050 ;
        RECT 697.950 66.600 700.050 67.050 ;
        RECT 514.950 65.400 700.050 66.600 ;
        RECT 514.950 64.950 517.050 65.400 ;
        RECT 577.950 64.950 580.050 65.400 ;
        RECT 697.950 64.950 700.050 65.400 ;
        RECT 757.950 66.600 760.050 67.050 ;
        RECT 808.950 66.600 811.050 67.050 ;
        RECT 757.950 65.400 811.050 66.600 ;
        RECT 757.950 64.950 760.050 65.400 ;
        RECT 808.950 64.950 811.050 65.400 ;
        RECT 931.950 66.600 934.050 67.050 ;
        RECT 949.950 66.600 952.050 67.050 ;
        RECT 973.950 66.600 976.050 67.050 ;
        RECT 931.950 65.400 976.050 66.600 ;
        RECT 931.950 64.950 934.050 65.400 ;
        RECT 949.950 64.950 952.050 65.400 ;
        RECT 973.950 64.950 976.050 65.400 ;
        RECT 1015.950 66.600 1018.050 67.050 ;
        RECT 1033.950 66.600 1036.050 67.050 ;
        RECT 1015.950 65.400 1036.050 66.600 ;
        RECT 1015.950 64.950 1018.050 65.400 ;
        RECT 1033.950 64.950 1036.050 65.400 ;
        RECT 82.950 63.600 85.050 64.050 ;
        RECT 94.950 63.600 97.050 64.050 ;
        RECT 82.950 62.400 97.050 63.600 ;
        RECT 82.950 61.950 85.050 62.400 ;
        RECT 94.950 61.950 97.050 62.400 ;
        RECT 169.950 63.600 172.050 64.050 ;
        RECT 175.950 63.600 178.050 64.050 ;
        RECT 199.950 63.600 202.050 64.050 ;
        RECT 418.950 63.600 421.050 64.050 ;
        RECT 427.950 63.600 430.050 64.050 ;
        RECT 169.950 62.400 202.050 63.600 ;
        RECT 169.950 61.950 172.050 62.400 ;
        RECT 175.950 61.950 178.050 62.400 ;
        RECT 199.950 61.950 202.050 62.400 ;
        RECT 371.400 62.400 430.050 63.600 ;
        RECT 73.950 60.600 76.050 61.200 ;
        RECT 88.950 60.600 91.050 61.050 ;
        RECT 124.950 60.600 127.050 61.200 ;
        RECT 73.950 59.400 127.050 60.600 ;
        RECT 73.950 59.100 76.050 59.400 ;
        RECT 88.950 58.950 91.050 59.400 ;
        RECT 124.950 59.100 127.050 59.400 ;
        RECT 145.950 60.750 148.050 61.200 ;
        RECT 208.950 60.750 211.050 61.200 ;
        RECT 145.950 59.550 211.050 60.750 ;
        RECT 214.950 60.600 217.050 61.200 ;
        RECT 145.950 59.100 148.050 59.550 ;
        RECT 208.950 59.100 211.050 59.550 ;
        RECT 212.400 59.400 217.050 60.600 ;
        RECT 202.950 57.600 205.050 58.050 ;
        RECT 212.400 57.600 213.600 59.400 ;
        RECT 214.950 59.100 217.050 59.400 ;
        RECT 238.950 60.600 241.050 61.200 ;
        RECT 250.950 60.600 253.050 61.050 ;
        RECT 238.950 59.400 253.050 60.600 ;
        RECT 238.950 59.100 241.050 59.400 ;
        RECT 250.950 58.950 253.050 59.400 ;
        RECT 283.950 60.600 286.050 61.200 ;
        RECT 313.950 60.600 316.050 61.200 ;
        RECT 283.950 59.400 316.050 60.600 ;
        RECT 283.950 59.100 286.050 59.400 ;
        RECT 313.950 59.100 316.050 59.400 ;
        RECT 346.950 60.600 349.050 61.200 ;
        RECT 364.950 60.600 367.050 61.200 ;
        RECT 371.400 60.600 372.600 62.400 ;
        RECT 418.950 61.950 421.050 62.400 ;
        RECT 427.950 61.950 430.050 62.400 ;
        RECT 541.950 63.600 544.050 64.050 ;
        RECT 841.950 63.750 844.050 64.200 ;
        RECT 850.950 63.750 853.050 64.200 ;
        RECT 541.950 62.400 573.600 63.600 ;
        RECT 541.950 61.950 544.050 62.400 ;
        RECT 346.950 59.400 372.600 60.600 ;
        RECT 379.950 60.750 382.050 61.200 ;
        RECT 391.950 60.750 394.050 61.200 ;
        RECT 379.950 59.550 394.050 60.750 ;
        RECT 346.950 59.100 349.050 59.400 ;
        RECT 364.950 59.100 367.050 59.400 ;
        RECT 379.950 59.100 382.050 59.550 ;
        RECT 391.950 59.100 394.050 59.550 ;
        RECT 400.950 60.750 403.050 61.200 ;
        RECT 415.950 60.750 418.050 61.200 ;
        RECT 400.950 60.600 418.050 60.750 ;
        RECT 433.950 60.600 436.050 61.200 ;
        RECT 400.950 59.550 436.050 60.600 ;
        RECT 400.950 59.100 403.050 59.550 ;
        RECT 415.950 59.400 436.050 59.550 ;
        RECT 415.950 59.100 418.050 59.400 ;
        RECT 433.950 59.100 436.050 59.400 ;
        RECT 547.950 60.750 550.050 61.200 ;
        RECT 568.950 60.750 571.050 61.200 ;
        RECT 547.950 59.550 571.050 60.750 ;
        RECT 547.950 59.100 550.050 59.550 ;
        RECT 568.950 59.100 571.050 59.550 ;
        RECT 572.400 60.600 573.600 62.400 ;
        RECT 841.950 62.550 853.050 63.750 ;
        RECT 841.950 62.100 844.050 62.550 ;
        RECT 850.950 62.100 853.050 62.550 ;
        RECT 925.950 63.600 928.050 64.050 ;
        RECT 934.950 63.600 937.050 64.050 ;
        RECT 925.950 62.400 937.050 63.600 ;
        RECT 925.950 61.950 928.050 62.400 ;
        RECT 934.950 61.950 937.050 62.400 ;
        RECT 943.950 63.600 946.050 64.050 ;
        RECT 952.950 63.600 955.050 64.050 ;
        RECT 943.950 62.400 955.050 63.600 ;
        RECT 943.950 61.950 946.050 62.400 ;
        RECT 952.950 61.950 955.050 62.400 ;
        RECT 595.950 60.600 598.050 61.200 ;
        RECT 572.400 59.400 598.050 60.600 ;
        RECT 595.950 59.100 598.050 59.400 ;
        RECT 604.950 60.750 607.050 61.200 ;
        RECT 622.950 60.750 625.050 61.200 ;
        RECT 604.950 59.550 625.050 60.750 ;
        RECT 604.950 59.100 607.050 59.550 ;
        RECT 622.950 59.100 625.050 59.550 ;
        RECT 634.950 60.750 637.050 61.200 ;
        RECT 640.950 60.750 643.050 61.200 ;
        RECT 634.950 59.550 643.050 60.750 ;
        RECT 634.950 59.100 637.050 59.550 ;
        RECT 640.950 59.100 643.050 59.550 ;
        RECT 646.950 60.750 649.050 61.200 ;
        RECT 652.950 60.750 655.050 61.200 ;
        RECT 646.950 59.550 655.050 60.750 ;
        RECT 646.950 59.100 649.050 59.550 ;
        RECT 652.950 59.100 655.050 59.550 ;
        RECT 658.950 60.750 661.050 61.200 ;
        RECT 664.950 60.750 667.050 61.200 ;
        RECT 658.950 59.550 667.050 60.750 ;
        RECT 658.950 59.100 661.050 59.550 ;
        RECT 664.950 59.100 667.050 59.550 ;
        RECT 673.950 58.950 676.050 61.050 ;
        RECT 691.950 60.600 694.050 61.200 ;
        RECT 700.950 60.600 703.050 61.050 ;
        RECT 691.950 59.400 703.050 60.600 ;
        RECT 691.950 59.100 694.050 59.400 ;
        RECT 700.950 58.950 703.050 59.400 ;
        RECT 712.950 60.600 715.050 61.200 ;
        RECT 727.950 60.750 730.050 61.200 ;
        RECT 742.950 60.750 745.050 61.200 ;
        RECT 727.950 60.600 745.050 60.750 ;
        RECT 712.950 59.550 745.050 60.600 ;
        RECT 712.950 59.400 730.050 59.550 ;
        RECT 712.950 59.100 715.050 59.400 ;
        RECT 727.950 59.100 730.050 59.400 ;
        RECT 742.950 59.100 745.050 59.550 ;
        RECT 754.950 60.600 757.050 61.050 ;
        RECT 763.950 60.600 766.050 61.200 ;
        RECT 754.950 59.400 766.050 60.600 ;
        RECT 754.950 58.950 757.050 59.400 ;
        RECT 763.950 59.100 766.050 59.400 ;
        RECT 937.950 60.600 940.050 61.050 ;
        RECT 946.950 60.750 949.050 61.200 ;
        RECT 955.950 60.750 958.050 61.200 ;
        RECT 946.950 60.600 958.050 60.750 ;
        RECT 937.950 59.550 958.050 60.600 ;
        RECT 937.950 59.400 949.050 59.550 ;
        RECT 937.950 58.950 940.050 59.400 ;
        RECT 946.950 59.100 949.050 59.400 ;
        RECT 955.950 59.100 958.050 59.550 ;
        RECT 964.950 60.600 967.050 61.050 ;
        RECT 976.950 60.600 979.050 61.200 ;
        RECT 964.950 59.400 979.050 60.600 ;
        RECT 964.950 58.950 967.050 59.400 ;
        RECT 976.950 59.100 979.050 59.400 ;
        RECT 994.950 60.750 997.050 61.200 ;
        RECT 1009.950 60.750 1012.050 61.200 ;
        RECT 994.950 59.550 1012.050 60.750 ;
        RECT 994.950 59.100 997.050 59.550 ;
        RECT 1009.950 59.100 1012.050 59.550 ;
        RECT 202.950 56.400 213.600 57.600 ;
        RECT 202.950 55.950 205.050 56.400 ;
        RECT 19.950 54.600 22.050 54.900 ;
        RECT 37.950 54.600 40.050 55.050 ;
        RECT 19.950 53.400 40.050 54.600 ;
        RECT 19.950 52.800 22.050 53.400 ;
        RECT 37.950 52.950 40.050 53.400 ;
        RECT 76.950 54.600 79.050 54.900 ;
        RECT 82.950 54.600 85.050 55.050 ;
        RECT 76.950 53.400 85.050 54.600 ;
        RECT 76.950 52.800 79.050 53.400 ;
        RECT 82.950 52.950 85.050 53.400 ;
        RECT 103.950 54.600 106.050 54.900 ;
        RECT 112.800 54.600 114.900 55.050 ;
        RECT 103.950 53.400 114.900 54.600 ;
        RECT 103.950 52.800 106.050 53.400 ;
        RECT 112.800 52.950 114.900 53.400 ;
        RECT 115.950 54.450 118.050 54.900 ;
        RECT 121.950 54.450 124.050 54.900 ;
        RECT 115.950 53.250 124.050 54.450 ;
        RECT 115.950 52.800 118.050 53.250 ;
        RECT 121.950 52.800 124.050 53.250 ;
        RECT 139.950 54.600 142.050 55.050 ;
        RECT 148.950 54.600 151.050 54.900 ;
        RECT 139.950 53.400 151.050 54.600 ;
        RECT 139.950 52.950 142.050 53.400 ;
        RECT 148.950 52.800 151.050 53.400 ;
        RECT 181.950 54.450 184.050 54.900 ;
        RECT 187.950 54.450 190.050 54.900 ;
        RECT 181.950 53.250 190.050 54.450 ;
        RECT 181.950 52.800 184.050 53.250 ;
        RECT 187.950 52.800 190.050 53.250 ;
        RECT 193.950 54.450 196.050 54.900 ;
        RECT 199.950 54.450 202.050 54.900 ;
        RECT 193.950 53.250 202.050 54.450 ;
        RECT 193.950 52.800 196.050 53.250 ;
        RECT 199.950 52.800 202.050 53.250 ;
        RECT 217.950 54.450 220.050 54.900 ;
        RECT 226.800 54.450 228.900 54.900 ;
        RECT 217.950 53.250 228.900 54.450 ;
        RECT 217.950 52.800 220.050 53.250 ;
        RECT 226.800 52.800 228.900 53.250 ;
        RECT 229.950 54.600 232.050 55.050 ;
        RECT 235.950 54.600 238.050 54.900 ;
        RECT 229.950 53.400 238.050 54.600 ;
        RECT 229.950 52.950 232.050 53.400 ;
        RECT 235.950 52.800 238.050 53.400 ;
        RECT 250.950 54.450 253.050 54.900 ;
        RECT 262.950 54.450 265.050 54.900 ;
        RECT 250.950 53.250 265.050 54.450 ;
        RECT 250.950 52.800 253.050 53.250 ;
        RECT 262.950 52.800 265.050 53.250 ;
        RECT 274.950 54.450 277.050 54.900 ;
        RECT 280.950 54.450 283.050 54.900 ;
        RECT 274.950 53.250 283.050 54.450 ;
        RECT 274.950 52.800 277.050 53.250 ;
        RECT 280.950 52.800 283.050 53.250 ;
        RECT 304.950 54.450 307.050 54.900 ;
        RECT 310.950 54.450 313.050 54.900 ;
        RECT 304.950 53.250 313.050 54.450 ;
        RECT 304.950 52.800 307.050 53.250 ;
        RECT 310.950 52.800 313.050 53.250 ;
        RECT 322.950 54.450 325.050 54.900 ;
        RECT 349.950 54.450 352.050 54.900 ;
        RECT 322.950 53.250 352.050 54.450 ;
        RECT 322.950 52.800 325.050 53.250 ;
        RECT 349.950 52.800 352.050 53.250 ;
        RECT 388.950 54.600 391.050 54.900 ;
        RECT 403.950 54.600 406.050 55.050 ;
        RECT 388.950 53.400 406.050 54.600 ;
        RECT 388.950 52.800 391.050 53.400 ;
        RECT 403.950 52.950 406.050 53.400 ;
        RECT 412.950 54.600 415.050 54.900 ;
        RECT 442.950 54.600 445.050 54.900 ;
        RECT 454.950 54.600 457.050 55.050 ;
        RECT 412.950 53.400 457.050 54.600 ;
        RECT 412.950 52.800 415.050 53.400 ;
        RECT 442.950 52.800 445.050 53.400 ;
        RECT 454.950 52.950 457.050 53.400 ;
        RECT 499.950 54.600 502.050 54.900 ;
        RECT 526.950 54.600 529.050 54.900 ;
        RECT 499.950 54.450 529.050 54.600 ;
        RECT 544.950 54.450 547.050 54.900 ;
        RECT 499.950 53.400 547.050 54.450 ;
        RECT 499.950 52.800 502.050 53.400 ;
        RECT 526.950 53.250 547.050 53.400 ;
        RECT 526.950 52.800 529.050 53.250 ;
        RECT 544.950 52.800 547.050 53.250 ;
        RECT 607.950 54.450 610.050 54.900 ;
        RECT 613.950 54.450 616.050 54.900 ;
        RECT 607.950 53.250 616.050 54.450 ;
        RECT 607.950 52.800 610.050 53.250 ;
        RECT 613.950 52.800 616.050 53.250 ;
        RECT 619.950 54.600 622.050 54.900 ;
        RECT 634.950 54.600 637.050 55.050 ;
        RECT 619.950 53.400 637.050 54.600 ;
        RECT 619.950 52.800 622.050 53.400 ;
        RECT 634.950 52.950 637.050 53.400 ;
        RECT 643.950 54.600 646.050 54.900 ;
        RECT 658.950 54.600 661.050 55.050 ;
        RECT 643.950 53.400 661.050 54.600 ;
        RECT 643.950 52.800 646.050 53.400 ;
        RECT 658.950 52.950 661.050 53.400 ;
        RECT 667.950 54.600 670.050 54.900 ;
        RECT 674.400 54.600 675.600 58.950 ;
        RECT 826.950 57.450 829.050 57.900 ;
        RECT 850.950 57.450 853.050 57.900 ;
        RECT 826.950 56.250 853.050 57.450 ;
        RECT 826.950 55.800 829.050 56.250 ;
        RECT 850.950 55.800 853.050 56.250 ;
        RECT 667.950 53.400 675.600 54.600 ;
        RECT 703.950 54.450 706.050 54.900 ;
        RECT 709.950 54.450 712.050 54.900 ;
        RECT 667.950 52.800 670.050 53.400 ;
        RECT 703.950 53.250 712.050 54.450 ;
        RECT 703.950 52.800 706.050 53.250 ;
        RECT 709.950 52.800 712.050 53.250 ;
        RECT 745.950 54.450 748.050 54.900 ;
        RECT 754.950 54.450 757.050 54.900 ;
        RECT 745.950 53.250 757.050 54.450 ;
        RECT 745.950 52.800 748.050 53.250 ;
        RECT 754.950 52.800 757.050 53.250 ;
        RECT 766.950 54.600 769.050 54.900 ;
        RECT 772.950 54.600 775.050 55.050 ;
        RECT 787.950 54.600 790.050 55.050 ;
        RECT 766.950 53.400 790.050 54.600 ;
        RECT 766.950 52.800 769.050 53.400 ;
        RECT 772.950 52.950 775.050 53.400 ;
        RECT 787.950 52.950 790.050 53.400 ;
        RECT 916.950 54.600 919.050 55.050 ;
        RECT 928.950 54.600 931.050 54.900 ;
        RECT 916.950 53.400 931.050 54.600 ;
        RECT 916.950 52.950 919.050 53.400 ;
        RECT 928.950 52.800 931.050 53.400 ;
        RECT 973.950 54.600 976.050 55.050 ;
        RECT 1006.950 54.600 1009.050 54.900 ;
        RECT 973.950 53.400 1009.050 54.600 ;
        RECT 973.950 52.950 976.050 53.400 ;
        RECT 1006.950 52.800 1009.050 53.400 ;
        RECT 43.950 51.600 46.050 52.050 ;
        RECT 70.950 51.600 73.050 52.050 ;
        RECT 85.950 51.600 88.050 52.050 ;
        RECT 43.950 50.400 88.050 51.600 ;
        RECT 43.950 49.950 46.050 50.400 ;
        RECT 70.950 49.950 73.050 50.400 ;
        RECT 85.950 49.950 88.050 50.400 ;
        RECT 127.950 51.600 130.050 52.050 ;
        RECT 154.950 51.600 157.050 52.050 ;
        RECT 166.950 51.600 169.050 52.050 ;
        RECT 127.950 50.400 169.050 51.600 ;
        RECT 127.950 49.950 130.050 50.400 ;
        RECT 154.950 49.950 157.050 50.400 ;
        RECT 166.950 49.950 169.050 50.400 ;
        RECT 367.950 51.600 370.050 52.050 ;
        RECT 379.950 51.600 382.050 52.050 ;
        RECT 367.950 50.400 382.050 51.600 ;
        RECT 367.950 49.950 370.050 50.400 ;
        RECT 379.950 49.950 382.050 50.400 ;
        RECT 922.950 51.600 925.050 52.050 ;
        RECT 943.950 51.600 946.050 52.050 ;
        RECT 955.950 51.600 958.050 52.050 ;
        RECT 922.950 50.400 958.050 51.600 ;
        RECT 922.950 49.950 925.050 50.400 ;
        RECT 943.950 49.950 946.050 50.400 ;
        RECT 955.950 49.950 958.050 50.400 ;
        RECT 97.950 48.600 100.050 49.050 ;
        RECT 112.950 48.600 115.050 49.050 ;
        RECT 97.950 47.400 115.050 48.600 ;
        RECT 167.400 48.600 168.600 49.950 ;
        RECT 247.950 48.600 250.050 49.050 ;
        RECT 256.950 48.600 259.050 49.050 ;
        RECT 397.950 48.600 400.050 49.050 ;
        RECT 421.950 48.600 424.050 49.050 ;
        RECT 167.400 47.400 424.050 48.600 ;
        RECT 97.950 46.950 100.050 47.400 ;
        RECT 112.950 46.950 115.050 47.400 ;
        RECT 247.950 46.950 250.050 47.400 ;
        RECT 256.950 46.950 259.050 47.400 ;
        RECT 397.950 46.950 400.050 47.400 ;
        RECT 421.950 46.950 424.050 47.400 ;
        RECT 436.950 48.600 439.050 49.050 ;
        RECT 457.950 48.600 460.050 49.050 ;
        RECT 436.950 47.400 460.050 48.600 ;
        RECT 436.950 46.950 439.050 47.400 ;
        RECT 457.950 46.950 460.050 47.400 ;
        RECT 469.950 48.600 472.050 49.050 ;
        RECT 505.950 48.600 508.050 49.050 ;
        RECT 469.950 47.400 508.050 48.600 ;
        RECT 469.950 46.950 472.050 47.400 ;
        RECT 505.950 46.950 508.050 47.400 ;
        RECT 565.950 48.600 568.050 49.050 ;
        RECT 586.950 48.600 589.050 49.050 ;
        RECT 565.950 47.400 589.050 48.600 ;
        RECT 565.950 46.950 568.050 47.400 ;
        RECT 586.950 46.950 589.050 47.400 ;
        RECT 652.950 48.600 655.050 49.050 ;
        RECT 688.950 48.600 691.050 49.050 ;
        RECT 787.950 48.600 790.050 49.050 ;
        RECT 652.950 47.400 790.050 48.600 ;
        RECT 652.950 46.950 655.050 47.400 ;
        RECT 688.950 46.950 691.050 47.400 ;
        RECT 787.950 46.950 790.050 47.400 ;
        RECT 982.950 48.600 985.050 49.050 ;
        RECT 994.950 48.600 997.050 49.050 ;
        RECT 1006.950 48.600 1009.050 49.050 ;
        RECT 982.950 47.400 1009.050 48.600 ;
        RECT 982.950 46.950 985.050 47.400 ;
        RECT 994.950 46.950 997.050 47.400 ;
        RECT 1006.950 46.950 1009.050 47.400 ;
        RECT 1036.950 48.600 1039.050 49.050 ;
        RECT 1042.950 48.600 1045.050 49.050 ;
        RECT 1036.950 47.400 1045.050 48.600 ;
        RECT 1036.950 46.950 1039.050 47.400 ;
        RECT 1042.950 46.950 1045.050 47.400 ;
        RECT 94.950 45.600 97.050 46.050 ;
        RECT 109.950 45.600 112.050 46.050 ;
        RECT 94.950 44.400 112.050 45.600 ;
        RECT 94.950 43.950 97.050 44.400 ;
        RECT 109.950 43.950 112.050 44.400 ;
        RECT 211.950 45.600 214.050 46.050 ;
        RECT 223.950 45.600 226.050 46.050 ;
        RECT 211.950 44.400 226.050 45.600 ;
        RECT 211.950 43.950 214.050 44.400 ;
        RECT 223.950 43.950 226.050 44.400 ;
        RECT 292.950 45.600 295.050 46.050 ;
        RECT 424.950 45.600 427.050 46.050 ;
        RECT 292.950 44.400 427.050 45.600 ;
        RECT 292.950 43.950 295.050 44.400 ;
        RECT 424.950 43.950 427.050 44.400 ;
        RECT 532.950 45.600 535.050 46.050 ;
        RECT 556.950 45.600 559.050 46.050 ;
        RECT 532.950 44.400 559.050 45.600 ;
        RECT 532.950 43.950 535.050 44.400 ;
        RECT 556.950 43.950 559.050 44.400 ;
        RECT 577.950 45.600 580.050 46.050 ;
        RECT 604.950 45.600 607.050 46.050 ;
        RECT 577.950 44.400 607.050 45.600 ;
        RECT 577.950 43.950 580.050 44.400 ;
        RECT 604.950 43.950 607.050 44.400 ;
        RECT 697.950 45.600 700.050 46.050 ;
        RECT 721.950 45.600 724.050 46.050 ;
        RECT 697.950 44.400 724.050 45.600 ;
        RECT 697.950 43.950 700.050 44.400 ;
        RECT 721.950 43.950 724.050 44.400 ;
        RECT 739.950 45.600 742.050 46.050 ;
        RECT 757.950 45.600 760.050 46.050 ;
        RECT 739.950 44.400 760.050 45.600 ;
        RECT 739.950 43.950 742.050 44.400 ;
        RECT 757.950 43.950 760.050 44.400 ;
        RECT 952.950 45.600 955.050 46.050 ;
        RECT 964.950 45.600 967.050 46.050 ;
        RECT 952.950 44.400 967.050 45.600 ;
        RECT 952.950 43.950 955.050 44.400 ;
        RECT 964.950 43.950 967.050 44.400 ;
        RECT 349.950 42.600 352.050 43.050 ;
        RECT 403.950 42.600 406.050 43.050 ;
        RECT 349.950 41.400 406.050 42.600 ;
        RECT 349.950 40.950 352.050 41.400 ;
        RECT 403.950 40.950 406.050 41.400 ;
        RECT 730.950 42.600 733.050 43.050 ;
        RECT 1021.950 42.600 1024.050 43.050 ;
        RECT 1036.950 42.600 1039.050 43.050 ;
        RECT 730.950 41.400 849.600 42.600 ;
        RECT 730.950 40.950 733.050 41.400 ;
        RECT 286.950 39.600 289.050 40.050 ;
        RECT 298.950 39.600 301.050 40.050 ;
        RECT 286.950 38.400 301.050 39.600 ;
        RECT 286.950 37.950 289.050 38.400 ;
        RECT 298.950 37.950 301.050 38.400 ;
        RECT 343.950 39.600 346.050 40.050 ;
        RECT 400.950 39.600 403.050 40.050 ;
        RECT 343.950 38.400 403.050 39.600 ;
        RECT 343.950 37.950 346.050 38.400 ;
        RECT 400.950 37.950 403.050 38.400 ;
        RECT 433.950 39.600 436.050 40.050 ;
        RECT 472.950 39.600 475.050 40.050 ;
        RECT 478.950 39.600 481.050 40.050 ;
        RECT 433.950 38.400 481.050 39.600 ;
        RECT 433.950 37.950 436.050 38.400 ;
        RECT 472.950 37.950 475.050 38.400 ;
        RECT 478.950 37.950 481.050 38.400 ;
        RECT 604.950 39.600 607.050 40.050 ;
        RECT 691.950 39.600 694.050 40.050 ;
        RECT 604.950 38.400 694.050 39.600 ;
        RECT 848.400 39.600 849.600 41.400 ;
        RECT 1021.950 41.400 1039.050 42.600 ;
        RECT 1021.950 40.950 1024.050 41.400 ;
        RECT 1036.950 40.950 1039.050 41.400 ;
        RECT 880.950 39.600 883.050 40.050 ;
        RECT 848.400 38.400 883.050 39.600 ;
        RECT 604.950 37.950 607.050 38.400 ;
        RECT 691.950 37.950 694.050 38.400 ;
        RECT 880.950 37.950 883.050 38.400 ;
        RECT 955.950 39.600 958.050 40.050 ;
        RECT 982.950 39.600 985.050 40.050 ;
        RECT 955.950 38.400 985.050 39.600 ;
        RECT 955.950 37.950 958.050 38.400 ;
        RECT 982.950 37.950 985.050 38.400 ;
        RECT 364.950 36.600 367.050 37.050 ;
        RECT 391.950 36.600 394.050 37.050 ;
        RECT 364.950 35.400 394.050 36.600 ;
        RECT 364.950 34.950 367.050 35.400 ;
        RECT 391.950 34.950 394.050 35.400 ;
        RECT 403.950 36.600 406.050 37.050 ;
        RECT 517.950 36.600 520.050 37.050 ;
        RECT 403.950 35.400 520.050 36.600 ;
        RECT 403.950 34.950 406.050 35.400 ;
        RECT 517.950 34.950 520.050 35.400 ;
        RECT 781.950 36.600 784.050 37.050 ;
        RECT 808.950 36.600 811.050 37.050 ;
        RECT 892.950 36.600 895.050 37.050 ;
        RECT 943.950 36.600 946.050 37.050 ;
        RECT 781.950 35.400 946.050 36.600 ;
        RECT 781.950 34.950 784.050 35.400 ;
        RECT 808.950 34.950 811.050 35.400 ;
        RECT 892.950 34.950 895.050 35.400 ;
        RECT 943.950 34.950 946.050 35.400 ;
        RECT 22.950 33.600 25.050 34.050 ;
        RECT 46.950 33.600 49.050 34.050 ;
        RECT 64.950 33.600 67.050 34.050 ;
        RECT 202.950 33.600 205.050 34.050 ;
        RECT 22.950 32.400 205.050 33.600 ;
        RECT 22.950 31.950 25.050 32.400 ;
        RECT 46.950 31.950 49.050 32.400 ;
        RECT 64.950 31.950 67.050 32.400 ;
        RECT 202.950 31.950 205.050 32.400 ;
        RECT 427.950 33.600 430.050 34.050 ;
        RECT 442.950 33.600 445.050 34.050 ;
        RECT 514.950 33.600 517.050 34.050 ;
        RECT 427.950 32.400 517.050 33.600 ;
        RECT 427.950 31.950 430.050 32.400 ;
        RECT 442.950 31.950 445.050 32.400 ;
        RECT 514.950 31.950 517.050 32.400 ;
        RECT 586.950 33.600 589.050 34.050 ;
        RECT 670.950 33.600 673.050 34.050 ;
        RECT 586.950 32.400 673.050 33.600 ;
        RECT 586.950 31.950 589.050 32.400 ;
        RECT 670.950 31.950 673.050 32.400 ;
        RECT 676.950 33.600 679.050 34.050 ;
        RECT 697.950 33.600 700.050 34.050 ;
        RECT 676.950 32.400 700.050 33.600 ;
        RECT 676.950 31.950 679.050 32.400 ;
        RECT 697.950 31.950 700.050 32.400 ;
        RECT 739.950 33.600 742.050 34.050 ;
        RECT 757.950 33.600 760.050 34.050 ;
        RECT 739.950 32.400 760.050 33.600 ;
        RECT 739.950 31.950 742.050 32.400 ;
        RECT 757.950 31.950 760.050 32.400 ;
        RECT 952.950 33.600 955.050 34.050 ;
        RECT 970.950 33.600 973.050 34.050 ;
        RECT 952.950 32.400 973.050 33.600 ;
        RECT 952.950 31.950 955.050 32.400 ;
        RECT 970.950 31.950 973.050 32.400 ;
        RECT 82.950 30.600 85.050 31.050 ;
        RECT 109.950 30.600 112.050 31.050 ;
        RECT 82.950 29.400 112.050 30.600 ;
        RECT 82.950 28.950 85.050 29.400 ;
        RECT 109.950 28.950 112.050 29.400 ;
        RECT 367.950 30.600 370.050 31.050 ;
        RECT 376.950 30.600 379.050 31.050 ;
        RECT 367.950 29.400 379.050 30.600 ;
        RECT 367.950 28.950 370.050 29.400 ;
        RECT 376.950 28.950 379.050 29.400 ;
        RECT 490.950 30.600 493.050 31.050 ;
        RECT 526.950 30.600 529.050 31.050 ;
        RECT 538.950 30.600 541.050 31.050 ;
        RECT 490.950 29.400 541.050 30.600 ;
        RECT 490.950 28.950 493.050 29.400 ;
        RECT 526.950 28.950 529.050 29.400 ;
        RECT 538.950 28.950 541.050 29.400 ;
        RECT 637.950 30.600 640.050 31.050 ;
        RECT 655.950 30.600 658.050 31.050 ;
        RECT 637.950 29.400 658.050 30.600 ;
        RECT 637.950 28.950 640.050 29.400 ;
        RECT 655.950 28.950 658.050 29.400 ;
        RECT 694.950 30.600 697.050 31.050 ;
        RECT 700.950 30.600 703.050 31.050 ;
        RECT 706.950 30.600 709.050 31.050 ;
        RECT 694.950 29.400 709.050 30.600 ;
        RECT 694.950 28.950 697.050 29.400 ;
        RECT 700.950 28.950 703.050 29.400 ;
        RECT 706.950 28.950 709.050 29.400 ;
        RECT 1015.950 30.600 1018.050 31.050 ;
        RECT 1024.950 30.600 1027.050 31.050 ;
        RECT 1015.950 29.400 1027.050 30.600 ;
        RECT 1015.950 28.950 1018.050 29.400 ;
        RECT 1024.950 28.950 1027.050 29.400 ;
        RECT 103.950 27.600 106.050 28.050 ;
        RECT 118.950 27.600 121.050 28.200 ;
        RECT 145.950 27.600 148.050 28.200 ;
        RECT 103.950 26.400 148.050 27.600 ;
        RECT 103.950 25.950 106.050 26.400 ;
        RECT 118.950 26.100 121.050 26.400 ;
        RECT 145.950 26.100 148.050 26.400 ;
        RECT 178.950 27.600 181.050 28.050 ;
        RECT 190.950 27.750 193.050 28.200 ;
        RECT 232.950 27.750 235.050 28.200 ;
        RECT 190.950 27.600 235.050 27.750 ;
        RECT 178.950 26.550 235.050 27.600 ;
        RECT 178.950 26.400 193.050 26.550 ;
        RECT 178.950 25.950 181.050 26.400 ;
        RECT 190.950 26.100 193.050 26.400 ;
        RECT 232.950 26.100 235.050 26.550 ;
        RECT 256.950 27.600 259.050 28.050 ;
        RECT 368.400 27.600 369.600 28.950 ;
        RECT 256.950 26.400 369.600 27.600 ;
        RECT 403.950 27.600 406.050 28.200 ;
        RECT 418.950 27.600 421.050 28.050 ;
        RECT 403.950 26.400 421.050 27.600 ;
        RECT 256.950 25.950 259.050 26.400 ;
        RECT 403.950 26.100 406.050 26.400 ;
        RECT 418.950 25.950 421.050 26.400 ;
        RECT 481.950 27.600 484.050 28.200 ;
        RECT 547.950 27.600 550.050 28.200 ;
        RECT 481.950 26.400 550.050 27.600 ;
        RECT 481.950 26.100 484.050 26.400 ;
        RECT 547.950 26.100 550.050 26.400 ;
        RECT 553.950 27.600 556.050 28.200 ;
        RECT 568.950 27.600 571.050 28.050 ;
        RECT 553.950 26.400 571.050 27.600 ;
        RECT 553.950 26.100 556.050 26.400 ;
        RECT 283.950 24.450 286.050 24.900 ;
        RECT 298.950 24.450 301.050 24.900 ;
        RECT 283.950 23.250 301.050 24.450 ;
        RECT 283.950 22.800 286.050 23.250 ;
        RECT 298.950 22.800 301.050 23.250 ;
        RECT 319.950 24.450 322.050 24.900 ;
        RECT 340.950 24.450 343.050 24.900 ;
        RECT 319.950 23.250 343.050 24.450 ;
        RECT 319.950 22.800 322.050 23.250 ;
        RECT 340.950 22.800 343.050 23.250 ;
        RECT 370.950 24.750 373.050 25.200 ;
        RECT 376.950 24.750 379.050 25.200 ;
        RECT 370.950 23.550 379.050 24.750 ;
        RECT 370.950 23.100 373.050 23.550 ;
        RECT 376.950 23.100 379.050 23.550 ;
        RECT 548.400 24.600 549.600 26.100 ;
        RECT 568.950 25.950 571.050 26.400 ;
        RECT 598.950 26.100 601.050 28.200 ;
        RECT 604.950 26.100 607.050 28.200 ;
        RECT 610.950 27.750 613.050 28.200 ;
        RECT 625.950 27.750 628.050 28.200 ;
        RECT 610.950 26.550 628.050 27.750 ;
        RECT 610.950 26.100 613.050 26.550 ;
        RECT 625.950 26.100 628.050 26.550 ;
        RECT 643.950 27.750 646.050 28.200 ;
        RECT 649.950 27.750 652.050 28.200 ;
        RECT 643.950 26.550 652.050 27.750 ;
        RECT 643.950 26.100 646.050 26.550 ;
        RECT 649.950 26.100 652.050 26.550 ;
        RECT 664.950 27.600 667.050 28.050 ;
        RECT 679.950 27.600 682.050 28.200 ;
        RECT 664.950 26.400 682.050 27.600 ;
        RECT 599.400 24.600 600.600 26.100 ;
        RECT 548.400 23.400 600.600 24.600 ;
        RECT 605.400 24.600 606.600 26.100 ;
        RECT 664.950 25.950 667.050 26.400 ;
        RECT 679.950 26.100 682.050 26.400 ;
        RECT 691.950 27.600 694.050 28.050 ;
        RECT 718.950 27.600 721.050 28.050 ;
        RECT 730.950 27.600 733.050 28.200 ;
        RECT 691.950 26.400 705.600 27.600 ;
        RECT 691.950 25.950 694.050 26.400 ;
        RECT 605.400 23.400 642.600 24.600 ;
        RECT 52.950 21.450 55.050 21.900 ;
        RECT 82.950 21.450 85.050 22.050 ;
        RECT 91.950 21.450 94.050 21.900 ;
        RECT 52.950 20.250 94.050 21.450 ;
        RECT 52.950 19.800 55.050 20.250 ;
        RECT 82.950 19.950 85.050 20.250 ;
        RECT 91.950 19.800 94.050 20.250 ;
        RECT 97.950 21.450 100.050 21.900 ;
        RECT 103.950 21.450 106.050 21.900 ;
        RECT 97.950 20.250 106.050 21.450 ;
        RECT 97.950 19.800 100.050 20.250 ;
        RECT 103.950 19.800 106.050 20.250 ;
        RECT 109.950 21.450 112.050 21.900 ;
        RECT 124.950 21.450 127.050 21.900 ;
        RECT 109.950 20.250 127.050 21.450 ;
        RECT 109.950 19.800 112.050 20.250 ;
        RECT 124.950 19.800 127.050 20.250 ;
        RECT 136.950 21.450 139.050 21.900 ;
        RECT 142.950 21.450 145.050 21.900 ;
        RECT 136.950 20.250 145.050 21.450 ;
        RECT 136.950 19.800 139.050 20.250 ;
        RECT 142.950 19.800 145.050 20.250 ;
        RECT 214.950 21.600 217.050 21.900 ;
        RECT 232.950 21.600 235.050 22.050 ;
        RECT 214.950 20.400 235.050 21.600 ;
        RECT 214.950 19.800 217.050 20.400 ;
        RECT 232.950 19.950 235.050 20.400 ;
        RECT 391.950 21.450 394.050 21.900 ;
        RECT 400.950 21.450 403.050 21.900 ;
        RECT 391.950 20.250 403.050 21.450 ;
        RECT 391.950 19.800 394.050 20.250 ;
        RECT 400.950 19.800 403.050 20.250 ;
        RECT 406.950 21.450 409.050 21.900 ;
        RECT 442.950 21.450 445.050 21.900 ;
        RECT 406.950 20.250 445.050 21.450 ;
        RECT 406.950 19.800 409.050 20.250 ;
        RECT 442.950 19.800 445.050 20.250 ;
        RECT 472.950 21.450 475.050 21.900 ;
        RECT 478.950 21.450 481.050 21.900 ;
        RECT 472.950 20.250 481.050 21.450 ;
        RECT 472.950 19.800 475.050 20.250 ;
        RECT 478.950 19.800 481.050 20.250 ;
        RECT 508.950 21.600 511.050 21.900 ;
        RECT 529.950 21.600 532.050 21.900 ;
        RECT 508.950 20.400 532.050 21.600 ;
        RECT 508.950 19.800 511.050 20.400 ;
        RECT 529.950 19.800 532.050 20.400 ;
        RECT 568.950 21.450 571.050 21.900 ;
        RECT 574.950 21.450 577.050 21.900 ;
        RECT 568.950 20.250 577.050 21.450 ;
        RECT 568.950 19.800 571.050 20.250 ;
        RECT 574.950 19.800 577.050 20.250 ;
        RECT 601.950 21.600 604.050 21.900 ;
        RECT 610.950 21.600 613.050 22.050 ;
        RECT 601.950 20.400 613.050 21.600 ;
        RECT 601.950 19.800 604.050 20.400 ;
        RECT 610.950 19.950 613.050 20.400 ;
        RECT 628.950 21.450 631.050 21.900 ;
        RECT 637.950 21.450 640.050 21.900 ;
        RECT 628.950 20.250 640.050 21.450 ;
        RECT 641.400 21.600 642.600 23.400 ;
        RECT 704.400 21.900 705.600 26.400 ;
        RECT 718.950 26.400 733.050 27.600 ;
        RECT 718.950 25.950 721.050 26.400 ;
        RECT 730.950 26.100 733.050 26.400 ;
        RECT 751.950 27.600 754.050 28.200 ;
        RECT 775.950 27.600 778.050 28.050 ;
        RECT 751.950 26.400 778.050 27.600 ;
        RECT 751.950 26.100 754.050 26.400 ;
        RECT 775.950 25.950 778.050 26.400 ;
        RECT 961.950 27.600 964.050 28.050 ;
        RECT 976.950 27.600 979.050 28.200 ;
        RECT 961.950 26.400 979.050 27.600 ;
        RECT 961.950 25.950 964.050 26.400 ;
        RECT 976.950 26.100 979.050 26.400 ;
        RECT 982.950 27.600 985.050 28.200 ;
        RECT 1000.950 27.600 1003.050 28.200 ;
        RECT 982.950 26.400 1003.050 27.600 ;
        RECT 982.950 26.100 985.050 26.400 ;
        RECT 1000.950 26.100 1003.050 26.400 ;
        RECT 916.950 24.600 919.050 24.900 ;
        RECT 958.950 24.600 961.050 25.050 ;
        RECT 916.950 23.400 921.600 24.600 ;
        RECT 916.950 22.800 919.050 23.400 ;
        RECT 652.950 21.600 655.050 21.900 ;
        RECT 641.400 21.450 655.050 21.600 ;
        RECT 664.950 21.450 667.050 21.900 ;
        RECT 641.400 20.400 667.050 21.450 ;
        RECT 628.950 19.800 631.050 20.250 ;
        RECT 637.950 19.800 640.050 20.250 ;
        RECT 652.950 20.250 667.050 20.400 ;
        RECT 652.950 19.800 655.050 20.250 ;
        RECT 664.950 19.800 667.050 20.250 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 676.950 21.450 679.050 21.900 ;
        RECT 670.950 20.250 679.050 21.450 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 676.950 19.800 679.050 20.250 ;
        RECT 682.950 21.450 685.050 21.900 ;
        RECT 694.950 21.450 697.050 21.900 ;
        RECT 682.950 20.250 697.050 21.450 ;
        RECT 682.950 19.800 685.050 20.250 ;
        RECT 694.950 19.800 697.050 20.250 ;
        RECT 703.950 19.800 706.050 21.900 ;
        RECT 709.950 21.450 712.050 21.900 ;
        RECT 718.950 21.450 721.050 21.900 ;
        RECT 709.950 20.250 721.050 21.450 ;
        RECT 709.950 19.800 712.050 20.250 ;
        RECT 718.950 19.800 721.050 20.250 ;
        RECT 727.950 21.600 730.050 21.900 ;
        RECT 760.950 21.600 763.050 21.900 ;
        RECT 796.950 21.600 799.050 22.050 ;
        RECT 727.950 20.400 799.050 21.600 ;
        RECT 920.400 21.600 921.600 23.400 ;
        RECT 958.950 23.400 975.600 24.600 ;
        RECT 958.950 22.950 961.050 23.400 ;
        RECT 961.950 21.600 964.050 22.050 ;
        RECT 974.400 21.900 975.600 23.400 ;
        RECT 920.400 20.400 964.050 21.600 ;
        RECT 727.950 19.800 730.050 20.400 ;
        RECT 760.950 19.800 763.050 20.400 ;
        RECT 796.950 19.950 799.050 20.400 ;
        RECT 961.950 19.950 964.050 20.400 ;
        RECT 973.950 19.800 976.050 21.900 ;
        RECT 1027.950 21.450 1030.050 21.900 ;
        RECT 1039.950 21.450 1042.050 21.900 ;
        RECT 1027.950 20.250 1042.050 21.450 ;
        RECT 1027.950 19.800 1030.050 20.250 ;
        RECT 1039.950 19.800 1042.050 20.250 ;
        RECT 307.950 18.600 310.050 18.900 ;
        RECT 316.950 18.600 319.050 18.900 ;
        RECT 307.950 18.450 319.050 18.600 ;
        RECT 361.950 18.450 364.050 18.900 ;
        RECT 307.950 17.400 364.050 18.450 ;
        RECT 307.950 16.800 310.050 17.400 ;
        RECT 316.950 17.250 364.050 17.400 ;
        RECT 316.950 16.800 319.050 17.250 ;
        RECT 361.950 16.800 364.050 17.250 ;
        RECT 538.950 18.600 541.050 19.050 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 538.950 17.400 553.050 18.600 ;
        RECT 538.950 16.950 541.050 17.400 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 556.950 16.950 559.050 19.050 ;
        RECT 730.950 18.600 733.050 19.050 ;
        RECT 739.950 18.600 742.050 19.050 ;
        RECT 730.950 17.400 742.050 18.600 ;
        RECT 730.950 16.950 733.050 17.400 ;
        RECT 739.950 16.950 742.050 17.400 ;
        RECT 850.950 18.600 853.050 19.050 ;
        RECT 859.950 18.600 862.050 18.900 ;
        RECT 886.950 18.600 889.050 18.900 ;
        RECT 850.950 18.450 889.050 18.600 ;
        RECT 892.950 18.450 895.050 18.900 ;
        RECT 850.950 17.400 895.050 18.450 ;
        RECT 850.950 16.950 853.050 17.400 ;
        RECT 460.950 15.600 463.050 16.050 ;
        RECT 484.950 15.600 487.050 16.050 ;
        RECT 502.950 15.600 505.050 16.050 ;
        RECT 460.950 14.400 505.050 15.600 ;
        RECT 460.950 13.950 463.050 14.400 ;
        RECT 484.950 13.950 487.050 14.400 ;
        RECT 502.950 13.950 505.050 14.400 ;
        RECT 529.950 15.600 532.050 16.050 ;
        RECT 553.950 15.600 556.050 16.050 ;
        RECT 529.950 14.400 556.050 15.600 ;
        RECT 529.950 13.950 532.050 14.400 ;
        RECT 553.950 13.950 556.050 14.400 ;
        RECT 205.950 12.600 208.050 13.050 ;
        RECT 370.950 12.600 373.050 13.050 ;
        RECT 205.950 11.400 373.050 12.600 ;
        RECT 205.950 10.950 208.050 11.400 ;
        RECT 370.950 10.950 373.050 11.400 ;
        RECT 418.950 12.600 421.050 13.050 ;
        RECT 557.400 12.600 558.600 16.950 ;
        RECT 859.950 16.800 862.050 17.400 ;
        RECT 886.950 17.250 895.050 17.400 ;
        RECT 886.950 16.800 889.050 17.250 ;
        RECT 892.950 16.800 895.050 17.250 ;
        RECT 937.950 18.600 940.050 19.050 ;
        RECT 979.950 18.600 982.050 19.050 ;
        RECT 937.950 17.400 982.050 18.600 ;
        RECT 937.950 16.950 940.050 17.400 ;
        RECT 979.950 16.950 982.050 17.400 ;
        RECT 559.950 15.600 562.050 16.050 ;
        RECT 622.950 15.600 625.050 16.050 ;
        RECT 559.950 14.400 625.050 15.600 ;
        RECT 559.950 13.950 562.050 14.400 ;
        RECT 622.950 13.950 625.050 14.400 ;
        RECT 658.950 15.600 661.050 16.050 ;
        RECT 703.950 15.600 706.050 16.050 ;
        RECT 658.950 14.400 706.050 15.600 ;
        RECT 658.950 13.950 661.050 14.400 ;
        RECT 703.950 13.950 706.050 14.400 ;
        RECT 715.950 15.600 718.050 16.050 ;
        RECT 835.950 15.600 838.050 16.050 ;
        RECT 715.950 14.400 838.050 15.600 ;
        RECT 715.950 13.950 718.050 14.400 ;
        RECT 835.950 13.950 838.050 14.400 ;
        RECT 643.950 12.600 646.050 13.050 ;
        RECT 418.950 11.400 646.050 12.600 ;
        RECT 418.950 10.950 421.050 11.400 ;
        RECT 643.950 10.950 646.050 11.400 ;
        RECT 370.950 6.600 373.050 7.050 ;
        RECT 541.950 6.600 544.050 7.050 ;
        RECT 733.950 6.600 736.050 7.050 ;
        RECT 754.950 6.600 757.050 7.050 ;
        RECT 370.950 5.400 757.050 6.600 ;
        RECT 370.950 4.950 373.050 5.400 ;
        RECT 541.950 4.950 544.050 5.400 ;
        RECT 733.950 4.950 736.050 5.400 ;
        RECT 754.950 4.950 757.050 5.400 ;
  END
END pong_pt1
END LIBRARY

