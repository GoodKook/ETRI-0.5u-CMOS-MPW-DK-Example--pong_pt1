* NGSPICE file created from pong_pt1.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR D S R CLK Q vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

.subckt pong_pt1 gnd vdd clk down hsync p_tick reset rgb[11] rgb[10] rgb[9] rgb[8]
+ rgb[7] rgb[6] rgb[5] rgb[4] rgb[3] rgb[2] rgb[1] rgb[0] up vsync
XFILL_3__1606_ vdd gnd FILL
XFILL_1__1670_ vdd gnd FILL
XFILL_3__1468_ vdd gnd FILL
XFILL_3__1537_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL_3__1399_ vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_4__1715_ vdd gnd FILL
XFILL_4__1577_ vdd gnd FILL
XFILL_4__1646_ vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL_2__1144_ vdd gnd FILL
XFILL_2__1075_ vdd gnd FILL
XFILL_0_CLKBUF1_insert6 vdd gnd FILL
XFILL_3__1322_ vdd gnd FILL
X_1270_ _1270_/A _1270_/B _1270_/C _1270_/D _1304_/C vdd gnd OAI22X1
XFILL_0__1613_ vdd gnd FILL
XFILL_3__888_ vdd gnd FILL
XFILL_3__957_ vdd gnd FILL
XFILL_0__1544_ vdd gnd FILL
XFILL_3__1184_ vdd gnd FILL
XFILL_4_BUFX2_insert3 vdd gnd FILL
XFILL_3__1253_ vdd gnd FILL
XFILL_0__1475_ vdd gnd FILL
X_1606_ _979_/C _979_/B _1672_/A vdd gnd NOR2X1
XFILL_1__1722_ vdd gnd FILL
XFILL_1__1653_ vdd gnd FILL
XFILL_4__1500_ vdd gnd FILL
X_1468_ _1485_/B _1487_/A _1500_/B vdd gnd NAND2X1
X_1537_ _1537_/A _1595_/B _1537_/C _1544_/D _1685_/D vdd gnd OAI22X1
X_1399_ _1545_/A _1410_/B _1399_/C _1417_/C _1408_/B vdd gnd AOI22X1
XFILL_4__1431_ vdd gnd FILL
XFILL_4__1362_ vdd gnd FILL
XFILL_1__1584_ vdd gnd FILL
XFILL_4__1293_ vdd gnd FILL
XFILL_2__975_ vdd gnd FILL
XFILL_1__1018_ vdd gnd FILL
X_981_ _981_/A _981_/B _981_/Y vdd gnd NOR2X1
XFILL_4__1629_ vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
XFILL_2__1058_ vdd gnd FILL
XFILL_2__1127_ vdd gnd FILL
X_1322_ _1355_/C _1356_/B _1414_/B vdd gnd NAND2X1
XFILL_1__993_ vdd gnd FILL
X_1253_ _1253_/A _1253_/B _1253_/C _1267_/B vdd gnd NAND3X1
X_1184_ _1216_/B _1184_/B _1353_/B _1213_/B _1185_/A vdd gnd AOI22X1
XFILL_0__1527_ vdd gnd FILL
XFILL_3__1236_ vdd gnd FILL
XFILL_3__1305_ vdd gnd FILL
XFILL_3__1167_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_0__1458_ vdd gnd FILL
XFILL_3__1098_ vdd gnd FILL
XFILL_4__1414_ vdd gnd FILL
XFILL_4__1345_ vdd gnd FILL
XFILL_1__1636_ vdd gnd FILL
XFILL_1__1567_ vdd gnd FILL
XFILL_1__1498_ vdd gnd FILL
XFILL_4__1276_ vdd gnd FILL
XFILL_2__889_ vdd gnd FILL
XFILL_2__958_ vdd gnd FILL
X_895_ _938_/Q _895_/B _947_/D vdd gnd NOR2X1
X_964_ _964_/A _965_/C vdd gnd INVX2
XFILL_2__1676_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
XFILL_0__1243_ vdd gnd FILL
XFILL_3__1021_ vdd gnd FILL
XFILL_0__1312_ vdd gnd FILL
X_1236_ _1698_/Q _1513_/A _1236_/C _1237_/A vdd gnd OAI21X1
X_1305_ _1305_/A _1305_/B _1305_/C _1307_/A vdd gnd NAND3X1
XFILL_1__976_ vdd gnd FILL
XFILL_1__1352_ vdd gnd FILL
XFILL_3__1219_ vdd gnd FILL
XBUFX2_insert0 _859_/Y _956_/R vdd gnd BUFX2
X_1167_ _1691_/Q _1690_/Q _1692_/Q _1332_/A vdd gnd OAI21X1
XFILL_1__1421_ vdd gnd FILL
XFILL_4__1061_ vdd gnd FILL
XFILL_1__1283_ vdd gnd FILL
XFILL_4__1130_ vdd gnd FILL
X_1098_ _1427_/B _961_/B _1099_/C vdd gnd XOR2X1
XFILL_4__1328_ vdd gnd FILL
XFILL_2__1530_ vdd gnd FILL
XFILL_2__1461_ vdd gnd FILL
XFILL_2__1392_ vdd gnd FILL
XFILL_1__1619_ vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
XFILL_4__1259_ vdd gnd FILL
XFILL_1__830_ vdd gnd FILL
X_947_ _947_/D vdd _947_/R _949_/CLK _964_/A vdd gnd DFFSR
X_878_ _878_/A _878_/B _937_/B _942_/D vdd gnd AOI21X1
XFILL_3__1570_ vdd gnd FILL
XFILL_2__1659_ vdd gnd FILL
XFILL_4__972_ vdd gnd FILL
X_1021_ _1422_/A _953_/Q _968_/A _1616_/B _1022_/A vdd gnd AOI22X1
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1157_ vdd gnd FILL
XFILL_3__1004_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
X_1219_ _1696_/Q _974_/A _1227_/A vdd gnd NAND2X1
XFILL_1__1404_ vdd gnd FILL
XFILL_1__959_ vdd gnd FILL
XFILL_4__1044_ vdd gnd FILL
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL_4__1113_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
XFILL_3__990_ vdd gnd FILL
XFILL_2__1513_ vdd gnd FILL
XFILL_2__1375_ vdd gnd FILL
XFILL_2__1444_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
X_1570_ _1570_/A _1577_/C _1572_/B vdd gnd NAND2X1
XFILL_3__1622_ vdd gnd FILL
XFILL_3__1484_ vdd gnd FILL
XFILL_3__1553_ vdd gnd FILL
X_1004_ _951_/Q _1383_/B _997_/Y _1011_/A vdd gnd OAI21X1
XFILL_4__886_ vdd gnd FILL
XFILL_1__1120_ vdd gnd FILL
XFILL_0__1209_ vdd gnd FILL
XFILL_1__1051_ vdd gnd FILL
XFILL_4__1593_ vdd gnd FILL
XFILL_4__1662_ vdd gnd FILL
X_1699_ _1699_/D vdd _1702_/R _1702_/CLK _999_/A vdd gnd DFFSR
XFILL_2__1160_ vdd gnd FILL
XFILL_1__1318_ vdd gnd FILL
XFILL_0__831_ vdd gnd FILL
XFILL_0__900_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_4__1027_ vdd gnd FILL
XFILL_2__1091_ vdd gnd FILL
XFILL_3__973_ vdd gnd FILL
XFILL_0__1560_ vdd gnd FILL
XFILL_2__1358_ vdd gnd FILL
XFILL_0__1491_ vdd gnd FILL
XFILL_2__1427_ vdd gnd FILL
XFILL_2__1289_ vdd gnd FILL
X_1622_ up _1657_/A vdd gnd INVX1
XFILL_3__1605_ vdd gnd FILL
X_1484_ _1488_/A _1488_/B _1484_/C _1485_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert14 vdd gnd FILL
X_1553_ _1553_/A _1619_/A _1553_/C _1691_/D vdd gnd OAI21X1
XFILL_3__1398_ vdd gnd FILL
XFILL_3__1467_ vdd gnd FILL
XFILL_3__1536_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_4__869_ vdd gnd FILL
XFILL_2__991_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_4__1714_ vdd gnd FILL
XFILL_1_BUFX2_insert0 vdd gnd FILL
XFILL_4__1576_ vdd gnd FILL
XFILL_4__1645_ vdd gnd FILL
XFILL_2__1212_ vdd gnd FILL
XFILL_2__1143_ vdd gnd FILL
XFILL_2__1074_ vdd gnd FILL
XFILL_0_CLKBUF1_insert7 vdd gnd FILL
XFILL103350x70350 vdd gnd FILL
XFILL_3__1321_ vdd gnd FILL
XFILL_3__1252_ vdd gnd FILL
XFILL_0__1612_ vdd gnd FILL
XFILL_3__887_ vdd gnd FILL
XFILL_0__1543_ vdd gnd FILL
XFILL_3__1183_ vdd gnd FILL
XFILL_0__1474_ vdd gnd FILL
X_1605_ _1605_/A _1605_/B _1698_/D vdd gnd XOR2X1
X_1536_ _1602_/C _1536_/B _1536_/C _1537_/C vdd gnd NAND3X1
XFILL_4__1361_ vdd gnd FILL
XFILL_1__1652_ vdd gnd FILL
XFILL_4__1430_ vdd gnd FILL
X_1398_ _1398_/A _1398_/B _1398_/C _1417_/C vdd gnd AOI21X1
XFILL_1__1583_ vdd gnd FILL
X_1467_ _1488_/A _1487_/A vdd gnd INVX1
XFILL_1__1721_ vdd gnd FILL
XFILL_4__1292_ vdd gnd FILL
XFILL_3__1519_ vdd gnd FILL
XFILL_1__1017_ vdd gnd FILL
XFILL_2__974_ vdd gnd FILL
X_980_ _980_/A _980_/B _981_/B vdd gnd NOR2X1
XFILL_4__1628_ vdd gnd FILL
XFILL_4__1559_ vdd gnd FILL
XFILL_0__1190_ vdd gnd FILL
XFILL_2__1126_ vdd gnd FILL
XFILL_2__1057_ vdd gnd FILL
X_1321_ _979_/C _1400_/C _1356_/B vdd gnd NAND2X1
XFILL_1__992_ vdd gnd FILL
X_1252_ _1252_/A _1252_/B _1252_/C _1253_/C vdd gnd AOI21X1
X_1183_ _1327_/C _1327_/B _1353_/B vdd gnd AND2X2
XFILL_0__1526_ vdd gnd FILL
XFILL_3__1235_ vdd gnd FILL
XFILL_3__1304_ vdd gnd FILL
XFILL_0__1457_ vdd gnd FILL
XFILL_3__1166_ vdd gnd FILL
XFILL_0__1388_ vdd gnd FILL
XFILL_3__1097_ vdd gnd FILL
X_1519_ _1524_/A _1519_/B _1524_/B _1520_/C vdd gnd NAND3X1
XFILL_4__1413_ vdd gnd FILL
XFILL_4__1344_ vdd gnd FILL
XFILL_1__1566_ vdd gnd FILL
XFILL_1__1635_ vdd gnd FILL
XFILL_2__957_ vdd gnd FILL
XFILL_1__1497_ vdd gnd FILL
XFILL_4__1275_ vdd gnd FILL
XFILL_2__888_ vdd gnd FILL
X_894_ _894_/A _894_/B _937_/B _946_/D vdd gnd AOI21X1
X_963_ _963_/A _963_/B _966_/A vdd gnd NAND2X1
XFILL_2__1675_ vdd gnd FILL
XFILL_3__1020_ vdd gnd FILL
XFILL_0__1311_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
XFILL_0__1242_ vdd gnd FILL
XFILL_2__1109_ vdd gnd FILL
X_1166_ _1324_/A _1324_/B _952_/Q _1177_/B vdd gnd OAI21X1
XBUFX2_insert1 _859_/Y _954_/S vdd gnd BUFX2
X_1235_ _1235_/A _1254_/C _1235_/C _1236_/C vdd gnd NAND3X1
XFILL_1__975_ vdd gnd FILL
XFILL_1__1420_ vdd gnd FILL
X_1304_ _1304_/A _1304_/B _1304_/C _1305_/C vdd gnd NOR3X1
XFILL_3__1218_ vdd gnd FILL
XFILL_1__1351_ vdd gnd FILL
XFILL_3__1149_ vdd gnd FILL
XFILL_4__1060_ vdd gnd FILL
XFILL_0__1509_ vdd gnd FILL
XFILL_1__1282_ vdd gnd FILL
X_1097_ _1109_/A _1542_/A _1427_/B vdd gnd XOR2X1
XFILL_4__1327_ vdd gnd FILL
XFILL_1__1618_ vdd gnd FILL
XFILL_4__1258_ vdd gnd FILL
XFILL_1__1549_ vdd gnd FILL
XFILL_2__1391_ vdd gnd FILL
XFILL_2__1460_ vdd gnd FILL
XFILL_4__1189_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
X_1020_ _1020_/A _979_/A _1422_/A vdd gnd OR2X2
X_946_ _946_/D _948_/R vdd _949_/CLK _961_/A vdd gnd DFFSR
X_877_ _885_/A _885_/C _965_/A _878_/B vdd gnd OAI21X1
XFILL_2__1658_ vdd gnd FILL
XFILL_4__971_ vdd gnd FILL
XFILL_3__1003_ vdd gnd FILL
XFILL_2__1589_ vdd gnd FILL
XFILL_0__1225_ vdd gnd FILL
XFILL_0__1156_ vdd gnd FILL
XFILL_0__1087_ vdd gnd FILL
X_1218_ _1226_/A _1218_/B _1225_/A vdd gnd NAND2X1
X_1149_ _1696_/Q _1599_/A vdd gnd INVX2
XFILL_1__1403_ vdd gnd FILL
XFILL_1__889_ vdd gnd FILL
XFILL_1__958_ vdd gnd FILL
XFILL_4__1112_ vdd gnd FILL
XFILL_4__1043_ vdd gnd FILL
XFILL_1__1196_ vdd gnd FILL
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
XFILL_2__1512_ vdd gnd FILL
XFILL_2__1374_ vdd gnd FILL
XFILL_2__1443_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_3__1552_ vdd gnd FILL
XFILL_3__1621_ vdd gnd FILL
X_929_ _934_/A _929_/B _929_/C _930_/B vdd gnd NAND3X1
X_1003_ _1374_/B _1374_/C _1383_/B vdd gnd NAND2X1
XFILL_3__1483_ vdd gnd FILL
XFILL_1__1050_ vdd gnd FILL
XFILL_0__1208_ vdd gnd FILL
X_1698_ _1698_/D vdd _1710_/R _945_/CLK _1698_/Q vdd gnd DFFSR
XFILL_4__1661_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
XFILL_4__1592_ vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_0__830_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_4__1026_ vdd gnd FILL
XFILL_2__1090_ vdd gnd FILL
XFILL_3__972_ vdd gnd FILL
XFILL_0__1490_ vdd gnd FILL
XFILL_2__1426_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_2__1288_ vdd gnd FILL
XFILL_0__959_ vdd gnd FILL
X_1552_ _1582_/A _1582_/B _1691_/Q _1553_/C vdd gnd OAI21X1
X_1621_ _1621_/A _1621_/B _1674_/B vdd gnd NOR2X1
XFILL_2_BUFX2_insert15 vdd gnd FILL
XFILL_3__1604_ vdd gnd FILL
XFILL_3__1535_ vdd gnd FILL
X_1483_ _1483_/A _1498_/A _1541_/A vdd gnd XNOR2X1
XFILL_2__990_ vdd gnd FILL
XFILL_3__1397_ vdd gnd FILL
XFILL_3__1466_ vdd gnd FILL
XFILL_4__937_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_4__868_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
XFILL_4__1713_ vdd gnd FILL
XFILL_4__1644_ vdd gnd FILL
XFILL_1_BUFX2_insert1 vdd gnd FILL
XFILL_4__1575_ vdd gnd FILL
XFILL_2__1211_ vdd gnd FILL
XFILL_4__1009_ vdd gnd FILL
XFILL_2__1073_ vdd gnd FILL
XFILL_2__1142_ vdd gnd FILL
XFILL_0_CLKBUF1_insert8 vdd gnd FILL
XFILL_3__886_ vdd gnd FILL
XFILL103350x89850 vdd gnd FILL
XFILL_3__1182_ vdd gnd FILL
XFILL_3__1320_ vdd gnd FILL
XFILL_3__1251_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
XFILL_0__1473_ vdd gnd FILL
XFILL_0__1542_ vdd gnd FILL
XFILL_0__1611_ vdd gnd FILL
XFILL_1__1720_ vdd gnd FILL
X_1604_ _1604_/A _1604_/B _1604_/C _1605_/A vdd gnd OAI21X1
X_1535_ _1535_/A _1535_/B _1602_/C vdd gnd NOR2X1
XFILL_4__1360_ vdd gnd FILL
XFILL_1__1651_ vdd gnd FILL
X_1397_ _1397_/A _1397_/B _1397_/C _1398_/C vdd gnd NAND3X1
X_1466_ _1484_/C _1466_/B _1488_/A vdd gnd NAND2X1
XFILL_4__1291_ vdd gnd FILL
XFILL_3__1518_ vdd gnd FILL
XFILL_1__1582_ vdd gnd FILL
XFILL_2__973_ vdd gnd FILL
XFILL_3__1449_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_4__1627_ vdd gnd FILL
XFILL_4__1489_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
XFILL103950x31350 vdd gnd FILL
XFILL_2__1125_ vdd gnd FILL
XFILL103050x19650 vdd gnd FILL
X_1320_ _978_/A _1348_/B _1348_/C _1355_/C vdd gnd NAND3X1
XFILL103650x66450 vdd gnd FILL
X_1182_ _1403_/B _1351_/B _1327_/C vdd gnd NAND2X1
XFILL_3__869_ vdd gnd FILL
X_1251_ _1266_/A _1266_/B _1265_/A _1270_/C vdd gnd AOI21X1
XFILL_1__991_ vdd gnd FILL
XFILL_3__1165_ vdd gnd FILL
XFILL_0__1525_ vdd gnd FILL
XFILL_3__1234_ vdd gnd FILL
XFILL_3__1303_ vdd gnd FILL
XFILL_0__1456_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
XFILL_3__1096_ vdd gnd FILL
XFILL_4__1412_ vdd gnd FILL
X_1518_ _1518_/A _1573_/B _1519_/B vdd gnd NOR2X1
X_1449_ _1595_/B _1619_/A vdd gnd INVX2
XFILL_4__1343_ vdd gnd FILL
XFILL_1__1565_ vdd gnd FILL
XFILL_1__1634_ vdd gnd FILL
XFILL_1__1496_ vdd gnd FILL
XFILL_4__1274_ vdd gnd FILL
XFILL_2__887_ vdd gnd FILL
X_893_ _893_/A _945_/D vdd gnd INVX1
X_962_ _962_/A _962_/B _963_/B vdd gnd NOR2X1
XFILL_2__1674_ vdd gnd FILL
XFILL_0__1241_ vdd gnd FILL
XFILL103950x43050 vdd gnd FILL
XFILL_0__1310_ vdd gnd FILL
XFILL_2__1039_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
XFILL_2__1108_ vdd gnd FILL
XFILL_1__974_ vdd gnd FILL
X_1303_ _1303_/A _1303_/B _1303_/C _1304_/B vdd gnd NAND3X1
XFILL_1__1350_ vdd gnd FILL
X_1165_ _1332_/B _1693_/Q _1694_/Q _1324_/A vdd gnd AOI21X1
XBUFX2_insert2 _859_/Y _947_/R vdd gnd BUFX2
X_1234_ _1252_/C _1252_/B _1254_/C vdd gnd AND2X2
X_1096_ _1096_/A _1107_/A _1109_/A vdd gnd NAND2X1
XFILL_3__1217_ vdd gnd FILL
XFILL_3__1148_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_0__1508_ vdd gnd FILL
XFILL_3__1079_ vdd gnd FILL
XFILL_4__1326_ vdd gnd FILL
XFILL_4__1188_ vdd gnd FILL
XFILL_1__1617_ vdd gnd FILL
XFILL_4__1257_ vdd gnd FILL
XFILL_1__1479_ vdd gnd FILL
XFILL_2__1390_ vdd gnd FILL
XFILL_1__1548_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
X_945_ _945_/D vdd _947_/R _945_/CLK _961_/B vdd gnd DFFSR
X_876_ _885_/B _880_/B _878_/A vdd gnd NAND2X1
XFILL_2__1588_ vdd gnd FILL
XFILL_2__1657_ vdd gnd FILL
XFILL_0__1224_ vdd gnd FILL
XFILL_4__970_ vdd gnd FILL
XFILL_3__1002_ vdd gnd FILL
XFILL_0__1155_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
XFILL102450x70350 vdd gnd FILL
XFILL_1__957_ vdd gnd FILL
X_1217_ _1226_/B _1217_/B _1218_/B vdd gnd NOR2X1
XFILL_4__1042_ vdd gnd FILL
X_1148_ _1604_/A _1315_/B _1605_/B _1395_/B vdd gnd OAI21X1
XFILL_1__1333_ vdd gnd FILL
XFILL_1__1402_ vdd gnd FILL
X_1079_ _981_/Y _1079_/B _1079_/C _1080_/C vdd gnd OAI21X1
XFILL_1__888_ vdd gnd FILL
XFILL_4__1111_ vdd gnd FILL
XFILL_1__1195_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_2__1442_ vdd gnd FILL
XFILL_2__1511_ vdd gnd FILL
XFILL_2__1373_ vdd gnd FILL
XFILL_4__1309_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
X_928_ _928_/A _928_/B _933_/A _929_/C vdd gnd OAI21X1
XFILL_3__1551_ vdd gnd FILL
XFILL_3__1620_ vdd gnd FILL
X_859_ reset _859_/Y vdd gnd INVX8
X_1002_ _998_/A _992_/A _992_/B _1374_/B vdd gnd NAND3X1
XFILL_3__1482_ vdd gnd FILL
XFILL_0__1207_ vdd gnd FILL
XFILL_4__884_ vdd gnd FILL
X_1697_ _1697_/D vdd _1710_/R _945_/CLK _1697_/Q vdd gnd DFFSR
XFILL_4__1591_ vdd gnd FILL
XFILL_0__1069_ vdd gnd FILL
XFILL_4__1660_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_1__1316_ vdd gnd FILL
XFILL_4__1025_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_3__971_ vdd gnd FILL
XFILL_2__1356_ vdd gnd FILL
XFILL_2__1425_ vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
XFILL_2__1287_ vdd gnd FILL
XFILL_0__889_ vdd gnd FILL
X_1551_ _1555_/B _1555_/A _1553_/A vdd gnd XNOR2X1
X_1482_ _1482_/A _1482_/B _1507_/A vdd gnd XOR2X1
X_1620_ _1670_/B _999_/A _1699_/D vdd gnd XOR2X1
XFILL_3__1603_ vdd gnd FILL
XFILL_3__1534_ vdd gnd FILL
XFILL_3__1465_ vdd gnd FILL
XFILL_4__936_ vdd gnd FILL
XFILL_3__1396_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_1__1032_ vdd gnd FILL
XFILL_4__867_ vdd gnd FILL
XFILL_4__1712_ vdd gnd FILL
XFILL_4__1643_ vdd gnd FILL
XFILL_4__1574_ vdd gnd FILL
XFILL_2__1210_ vdd gnd FILL
XFILL_1_BUFX2_insert2 vdd gnd FILL
XFILL_4__1008_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_2__1072_ vdd gnd FILL
XFILL_0_CLKBUF1_insert9 vdd gnd FILL
XFILL_3__885_ vdd gnd FILL
XFILL_0__1610_ vdd gnd FILL
XFILL_3__1181_ vdd gnd FILL
XFILL_3__1250_ vdd gnd FILL
XFILL_2__1339_ vdd gnd FILL
XFILL_0__1472_ vdd gnd FILL
XFILL_0__1541_ vdd gnd FILL
XFILL_2__1408_ vdd gnd FILL
X_1603_ _1604_/B _1710_/Q _1603_/C _1604_/C vdd gnd AOI21X1
X_1534_ _1534_/A _1534_/B _1535_/B vdd gnd NAND2X1
X_1465_ _1537_/A _1473_/B _1466_/B vdd gnd NAND2X1
XFILL_1__1650_ vdd gnd FILL
X_1396_ _1428_/B _1397_/A vdd gnd INVX1
XFILL_1__1581_ vdd gnd FILL
XFILL_3__1517_ vdd gnd FILL
XFILL_4__1290_ vdd gnd FILL
XFILL_3__1448_ vdd gnd FILL
XFILL_4__919_ vdd gnd FILL
XFILL_2__972_ vdd gnd FILL
XFILL_3__1379_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_4__1557_ vdd gnd FILL
XFILL_4__1626_ vdd gnd FILL
XFILL_4__1488_ vdd gnd FILL
XFILL_2__1055_ vdd gnd FILL
XFILL_2__1124_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
X_1181_ _1694_/Q _1693_/Q _1332_/B _1351_/B vdd gnd NAND3X1
XFILL_3__937_ vdd gnd FILL
X_1250_ _1253_/A _1253_/B _1250_/C _1266_/A vdd gnd NAND3X1
XFILL_3__868_ vdd gnd FILL
XFILL_0__1524_ vdd gnd FILL
XFILL_3__1302_ vdd gnd FILL
XFILL_3__1164_ vdd gnd FILL
XFILL_0__1386_ vdd gnd FILL
XFILL_3__1233_ vdd gnd FILL
XFILL_3__1095_ vdd gnd FILL
XFILL_0__1455_ vdd gnd FILL
XFILL_4__1411_ vdd gnd FILL
XFILL_1__1633_ vdd gnd FILL
X_1517_ _1546_/B _1573_/B vdd gnd INVX1
X_1448_ _1582_/A _1582_/B _1595_/B vdd gnd NOR2X1
XFILL_4__1342_ vdd gnd FILL
X_1379_ _1379_/A _1612_/A _1379_/C _1381_/B vdd gnd NAND3X1
XFILL_4__1273_ vdd gnd FILL
XFILL_1__1564_ vdd gnd FILL
XFILL_1__1495_ vdd gnd FILL
XFILL_2__886_ vdd gnd FILL
X_961_ _961_/A _961_/B _963_/A vdd gnd NOR2X1
X_892_ _935_/A _894_/B _892_/C _893_/A vdd gnd NAND3X1
XFILL_4__1609_ vdd gnd FILL
XFILL_2__1673_ vdd gnd FILL
XFILL_0__1240_ vdd gnd FILL
XFILL_2__1038_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
XFILL_2__1107_ vdd gnd FILL
X_1233_ _1245_/B _1252_/A _1252_/C vdd gnd NOR2X1
XFILL_1__973_ vdd gnd FILL
X_1302_ _1302_/A _1302_/B _1302_/C _1303_/B vdd gnd NAND3X1
X_1164_ _1556_/A _1559_/A _1549_/A _1332_/B vdd gnd NAND3X1
XBUFX2_insert3 _859_/Y _948_/R vdd gnd BUFX2
XFILL_1__1280_ vdd gnd FILL
X_1095_ _1687_/Q _1542_/A vdd gnd INVX2
XFILL_0__1507_ vdd gnd FILL
XFILL_3__1216_ vdd gnd FILL
XFILL_3__1147_ vdd gnd FILL
XFILL_0__1438_ vdd gnd FILL
XFILL_3__1078_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_4__1325_ vdd gnd FILL
XFILL_1__1616_ vdd gnd FILL
XFILL_4__1187_ vdd gnd FILL
XFILL_1__1547_ vdd gnd FILL
XFILL_4__1256_ vdd gnd FILL
XFILL_1__1478_ vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_2__869_ vdd gnd FILL
XFILL_2__1725_ vdd gnd FILL
X_944_ _944_/D vdd _947_/R _945_/CLK _962_/A vdd gnd DFFSR
X_875_ _885_/A _885_/C _880_/B vdd gnd NOR2X1
XFILL_2__1587_ vdd gnd FILL
XFILL_2__1656_ vdd gnd FILL
XFILL_0__1223_ vdd gnd FILL
XFILL_0__1154_ vdd gnd FILL
XFILL_3__1001_ vdd gnd FILL
XFILL_0__1085_ vdd gnd FILL
X_1216_ _1694_/Q _1216_/B _1217_/B vdd gnd NOR2X1
XFILL_1__887_ vdd gnd FILL
XFILL_4__1041_ vdd gnd FILL
XFILL_1__1401_ vdd gnd FILL
X_1147_ _1696_/Q _1317_/B _1317_/A _1315_/B vdd gnd NAND3X1
XFILL_1__1332_ vdd gnd FILL
X_1078_ _1078_/A _974_/Y _1079_/B vdd gnd AND2X2
XFILL_1__1263_ vdd gnd FILL
XFILL_4__1110_ vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL_2__1441_ vdd gnd FILL
XFILL_2__1510_ vdd gnd FILL
XFILL_2__1372_ vdd gnd FILL
XFILL_4__1308_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
XFILL103950x4050 vdd gnd FILL
XFILL_4__1239_ vdd gnd FILL
X_927_ _953_/Q _933_/A vdd gnd INVX1
X_858_ _938_/D _858_/B _858_/C _858_/Y vdd gnd NOR3X1
XFILL_3__1481_ vdd gnd FILL
XFILL_3__1550_ vdd gnd FILL
X_1001_ _997_/A _1379_/A _998_/Y _1374_/C vdd gnd OAI21X1
XFILL_2__1639_ vdd gnd FILL
XCLKBUF1_insert10 clk _1689_/CLK vdd gnd CLKBUF1
XFILL_0__1206_ vdd gnd FILL
XFILL_4__883_ vdd gnd FILL
XFILL_0__1137_ vdd gnd FILL
XFILL102750x66450 vdd gnd FILL
XFILL_4__1590_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
X_1696_ _1696_/D vdd _1708_/R _945_/CLK _1696_/Q vdd gnd DFFSR
XFILL_1__1315_ vdd gnd FILL
XFILL_4__1024_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_3__970_ vdd gnd FILL
XFILL_2__1355_ vdd gnd FILL
XFILL_2__1424_ vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
XFILL_2__1286_ vdd gnd FILL
XFILL_3__1602_ vdd gnd FILL
XFILL_0__888_ vdd gnd FILL
X_1481_ _1481_/A _1481_/B _1482_/A vdd gnd NAND2X1
X_1550_ _1691_/Q _1709_/Q _1555_/B vdd gnd XOR2X1
XFILL_3__1533_ vdd gnd FILL
XFILL_3__1464_ vdd gnd FILL
XFILL_4__935_ vdd gnd FILL
XFILL_3__1395_ vdd gnd FILL
XFILL_4__866_ vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_1__1031_ vdd gnd FILL
XFILL_4__1711_ vdd gnd FILL
XFILL_1_BUFX2_insert3 vdd gnd FILL
XFILL_4__1642_ vdd gnd FILL
XFILL_4__1573_ vdd gnd FILL
X_1679_ _1679_/D _1702_/R vdd _1702_/CLK _1679_/Q vdd gnd DFFSR
XFILL_2__1140_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_4__1007_ vdd gnd FILL
XFILL_2__1071_ vdd gnd FILL
XFILL_3__884_ vdd gnd FILL
XFILL_0__1540_ vdd gnd FILL
XFILL_2__1338_ vdd gnd FILL
XFILL_3__1180_ vdd gnd FILL
XFILL_2__1407_ vdd gnd FILL
XFILL_2__1269_ vdd gnd FILL
XFILL_0__1471_ vdd gnd FILL
X_1602_ _1697_/Q _1710_/Q _1602_/C _1603_/C vdd gnd OAI21X1
X_1395_ _1395_/A _1395_/B _1674_/C _1428_/B vdd gnd AOI21X1
X_1533_ _1533_/A _1533_/B _1534_/B vdd gnd NOR2X1
X_1464_ _1685_/Q _1680_/Q _1484_/C vdd gnd NAND2X1
XFILL_3__1378_ vdd gnd FILL
XFILL_3__1516_ vdd gnd FILL
XFILL_3__1447_ vdd gnd FILL
XFILL_1__1580_ vdd gnd FILL
XFILL_0__1669_ vdd gnd FILL
XFILL_4__918_ vdd gnd FILL
XFILL_2__971_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL_4__849_ vdd gnd FILL
XFILL_4__1556_ vdd gnd FILL
XFILL_4__1487_ vdd gnd FILL
XFILL_4__1625_ vdd gnd FILL
XFILL_2__1123_ vdd gnd FILL
XFILL_2__1054_ vdd gnd FILL
XFILL_3__936_ vdd gnd FILL
X_1180_ _1695_/Q _1403_/B vdd gnd INVX2
XFILL_3__1232_ vdd gnd FILL
XFILL_3__867_ vdd gnd FILL
XFILL_0__1523_ vdd gnd FILL
XFILL_3__1301_ vdd gnd FILL
XFILL_3__1163_ vdd gnd FILL
XFILL_0__1385_ vdd gnd FILL
XFILL_0__1454_ vdd gnd FILL
XFILL_3__1094_ vdd gnd FILL
X_1516_ _1516_/A _1516_/B _1546_/B vdd gnd NOR2X1
XFILL_4__1341_ vdd gnd FILL
X_1378_ _1549_/A _999_/Y _1556_/A _1379_/C vdd gnd OAI21X1
X_1447_ _965_/C _1447_/B _1534_/A _1582_/A vdd gnd NAND3X1
XFILL_1__1632_ vdd gnd FILL
XFILL_4__1410_ vdd gnd FILL
XFILL_4__1272_ vdd gnd FILL
XFILL_1__1494_ vdd gnd FILL
XFILL_1__1563_ vdd gnd FILL
XFILL_2__885_ vdd gnd FILL
XFILL_4__1608_ vdd gnd FILL
X_891_ _891_/A _891_/B _892_/C vdd gnd NAND2X1
X_960_ _960_/A _965_/A _965_/B _967_/A vdd gnd NAND3X1
XFILL_2__1672_ vdd gnd FILL
XFILL_4__1539_ vdd gnd FILL
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1106_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
XFILL_3__919_ vdd gnd FILL
X_1232_ _1232_/A _1243_/A _1252_/A vdd gnd NAND2X1
XFILL_1__972_ vdd gnd FILL
XFILL102750x7950 vdd gnd FILL
X_1301_ _964_/A _1545_/A _1302_/A vdd gnd NAND2X1
XFILL_3__1215_ vdd gnd FILL
X_1163_ _1583_/A _1573_/A _1406_/A _1324_/B vdd gnd NOR3X1
XFILL_0__1437_ vdd gnd FILL
X_1094_ _1293_/B _1427_/A _1099_/B vdd gnd NAND2X1
XFILL_0__1506_ vdd gnd FILL
XFILL_3__1146_ vdd gnd FILL
XFILL_3__1077_ vdd gnd FILL
XFILL_0__1368_ vdd gnd FILL
XFILL_0__1299_ vdd gnd FILL
XFILL_4__1324_ vdd gnd FILL
XFILL_1__1615_ vdd gnd FILL
XFILL_1__1546_ vdd gnd FILL
XFILL_4__1186_ vdd gnd FILL
XFILL_2__937_ vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_4__1255_ vdd gnd FILL
XFILL_1__1477_ vdd gnd FILL
XFILL_2__868_ vdd gnd FILL
XFILL_2__1724_ vdd gnd FILL
X_874_ _965_/A _885_/B vdd gnd INVX1
XFILL_2__1655_ vdd gnd FILL
X_943_ _943_/D vdd _947_/R _945_/CLK _962_/B vdd gnd DFFSR
XFILL_2__1586_ vdd gnd FILL
XFILL_3__1000_ vdd gnd FILL
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1222_ vdd gnd FILL
XFILL_0__1084_ vdd gnd FILL
X_1215_ _952_/Q _1583_/A _1226_/B vdd gnd NOR2X1
XFILL_1__1400_ vdd gnd FILL
X_1146_ _1695_/Q _1694_/Q _1317_/B vdd gnd AND2X2
XFILL_1__886_ vdd gnd FILL
XFILL_1__1193_ vdd gnd FILL
XFILL_4__1040_ vdd gnd FILL
XFILL_1__1331_ vdd gnd FILL
X_1077_ _856_/Y _1306_/C vdd gnd INVX1
XFILL_1__1262_ vdd gnd FILL
XFILL_3__1129_ vdd gnd FILL
XFILL_2__1440_ vdd gnd FILL
XFILL_2__1371_ vdd gnd FILL
XFILL_1__1529_ vdd gnd FILL
XFILL_4__1307_ vdd gnd FILL
XFILL_4__1238_ vdd gnd FILL
XFILL_4__1169_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
X_1000_ _984_/B _999_/Y _1379_/A vdd gnd NAND2X1
X_926_ _953_/Q _932_/C _929_/B vdd gnd NAND2X1
X_857_ _938_/Q _938_/D vdd gnd INVX2
XFILL_3__1480_ vdd gnd FILL
XFILL_2__1638_ vdd gnd FILL
XFILL_2__1569_ vdd gnd FILL
XFILL_4__882_ vdd gnd FILL
XFILL_0__1205_ vdd gnd FILL
XFILL_0__1067_ vdd gnd FILL
XFILL_0__1136_ vdd gnd FILL
X_1695_ _1695_/D vdd _1709_/S _1709_/CLK _1695_/Q vdd gnd DFFSR
XFILL_1__869_ vdd gnd FILL
X_1129_ _958_/A _1520_/A _1260_/A vdd gnd NAND2X1
XFILL_1__1176_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_4__1023_ vdd gnd FILL
XFILL_1__1314_ vdd gnd FILL
XFILL_2__1354_ vdd gnd FILL
XFILL_2__1423_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_0__887_ vdd gnd FILL
XFILL_1_CLKBUF1_insert4 vdd gnd FILL
XFILL_3__1601_ vdd gnd FILL
XFILL_3__1532_ vdd gnd FILL
X_1480_ _1480_/A _1481_/B vdd gnd INVX1
X_909_ _915_/A _915_/B _910_/B vdd gnd NAND2X1
XFILL_3__1463_ vdd gnd FILL
XFILL_3__1394_ vdd gnd FILL
XFILL_4__934_ vdd gnd FILL
XFILL_1__1030_ vdd gnd FILL
XFILL_4__865_ vdd gnd FILL
XFILL_4__1641_ vdd gnd FILL
XFILL_0__1119_ vdd gnd FILL
X_1678_ _1678_/D vdd _1702_/R _1702_/CLK _1678_/Q vdd gnd DFFSR
XFILL_4__1572_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_4__1006_ vdd gnd FILL
XFILL_2__1070_ vdd gnd FILL
XFILL_3__883_ vdd gnd FILL
XFILL_2__1406_ vdd gnd FILL
XFILL_0__1470_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
XFILL_2__1268_ vdd gnd FILL
XFILL_2__1199_ vdd gnd FILL
X_1601_ _1601_/A _1604_/A _1697_/D vdd gnd XOR2X1
X_1532_ _968_/A _959_/A _1532_/C _1533_/B vdd gnd NAND3X1
XFILL_3__1515_ vdd gnd FILL
X_1463_ _1686_/Q _1680_/Q _1485_/B vdd gnd XOR2X1
X_1394_ _1394_/A _1394_/B _1397_/C vdd gnd NOR2X1
XFILL_2__970_ vdd gnd FILL
XFILL_3__1377_ vdd gnd FILL
XFILL_3__1446_ vdd gnd FILL
XFILL_0__1599_ vdd gnd FILL
XFILL_0__1668_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_4__917_ vdd gnd FILL
XFILL_4__848_ vdd gnd FILL
XFILL_4__1624_ vdd gnd FILL
XFILL_4__1555_ vdd gnd FILL
XFILL_4__1486_ vdd gnd FILL
XFILL_2__1053_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_3__935_ vdd gnd FILL
XFILL_3__866_ vdd gnd FILL
XFILL_3__1162_ vdd gnd FILL
XFILL_3__1231_ vdd gnd FILL
XFILL_0__1453_ vdd gnd FILL
XFILL_0__1522_ vdd gnd FILL
XFILL_3__1300_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
XFILL_3__1093_ vdd gnd FILL
X_1515_ _1534_/A _1515_/B _1516_/B vdd gnd NAND2X1
XFILL_4__1340_ vdd gnd FILL
X_1377_ _993_/A _999_/A _1612_/A vdd gnd NAND2X1
X_1446_ _1513_/C _1509_/C _1447_/B vdd gnd AND2X2
XFILL_1__1631_ vdd gnd FILL
XFILL_1__1562_ vdd gnd FILL
XFILL_3__1429_ vdd gnd FILL
XFILL_1__1493_ vdd gnd FILL
XFILL_2__884_ vdd gnd FILL
X_890_ _961_/B _890_/B _890_/C _894_/B vdd gnd NAND3X1
XFILL_4__1607_ vdd gnd FILL
XFILL_2__1671_ vdd gnd FILL
XFILL_4__1469_ vdd gnd FILL
XFILL_4__1538_ vdd gnd FILL
XFILL_2__1036_ vdd gnd FILL
XFILL_2__1105_ vdd gnd FILL
XFILL_3__918_ vdd gnd FILL
X_1162_ _1694_/Q _1583_/A vdd gnd INVX2
X_1231_ _1231_/A _1231_/B _1235_/A vdd gnd NOR2X1
XFILL_1__971_ vdd gnd FILL
XFILL_3__849_ vdd gnd FILL
X_1300_ _1300_/A _1300_/B _1302_/C vdd gnd NAND2X1
XFILL_3__1214_ vdd gnd FILL
XFILL_3__1145_ vdd gnd FILL
XFILL_0__1436_ vdd gnd FILL
X_1093_ _1394_/A _1427_/A vdd gnd INVX1
XFILL_0__1505_ vdd gnd FILL
XFILL_0__1367_ vdd gnd FILL
XFILL_3__1076_ vdd gnd FILL
XFILL_0__1298_ vdd gnd FILL
X_1429_ _1429_/A _1429_/B _1429_/C _1430_/C vdd gnd OAI21X1
XFILL_4__1323_ vdd gnd FILL
XFILL_4__1254_ vdd gnd FILL
XFILL_1__1614_ vdd gnd FILL
XFILL_1__1476_ vdd gnd FILL
XFILL_1__1545_ vdd gnd FILL
XFILL_4__1185_ vdd gnd FILL
XFILL_2__936_ vdd gnd FILL
XFILL103350x7950 vdd gnd FILL
XFILL_1_CLKBUF1_insert10 vdd gnd FILL
XFILL_2__867_ vdd gnd FILL
X_873_ _885_/A _885_/C _873_/C _941_/D vdd gnd AOI21X1
X_942_ _942_/D vdd _947_/R _945_/CLK _965_/A vdd gnd DFFSR
XFILL_2__1654_ vdd gnd FILL
XFILL_2__1585_ vdd gnd FILL
XFILL_2__1723_ vdd gnd FILL
XFILL_0__1221_ vdd gnd FILL
XFILL103350x85950 vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
XFILL_2__1019_ vdd gnd FILL
XFILL_0__1083_ vdd gnd FILL
X_1214_ _1226_/C _1214_/B _1226_/A vdd gnd NOR2X1
X_1145_ _1338_/A _1559_/A _1573_/A _1317_/A vdd gnd AOI21X1
XFILL_1__1330_ vdd gnd FILL
XFILL_1__885_ vdd gnd FILL
XFILL_1__1192_ vdd gnd FILL
XFILL_0__1419_ vdd gnd FILL
XFILL_3__1128_ vdd gnd FILL
XFILL_1__1261_ vdd gnd FILL
X_1076_ _1307_/B _1723_/A vdd gnd INVX1
XFILL_3__1059_ vdd gnd FILL
XFILL_1__1528_ vdd gnd FILL
XFILL_4__1237_ vdd gnd FILL
XFILL_4__1168_ vdd gnd FILL
XFILL_4__1306_ vdd gnd FILL
XFILL_2__1370_ vdd gnd FILL
XFILL_1__1459_ vdd gnd FILL
XFILL_2__919_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
XFILL_4__1099_ vdd gnd FILL
X_925_ _925_/A _928_/A _925_/C _932_/C vdd gnd NOR3X1
XFILL103050x15750 vdd gnd FILL
X_856_ _858_/B _858_/C _856_/Y vdd gnd NOR2X1
XFILL103650x62550 vdd gnd FILL
XFILL_2__1568_ vdd gnd FILL
XFILL_2__1637_ vdd gnd FILL
XFILL_0__1204_ vdd gnd FILL
XFILL_4__881_ vdd gnd FILL
XFILL_2__1499_ vdd gnd FILL
X_1694_ _1694_/D vdd _1709_/S _1710_/CLK _1694_/Q vdd gnd DFFSR
XFILL_0__1066_ vdd gnd FILL
XFILL_0__1135_ vdd gnd FILL
XFILL_1__937_ vdd gnd FILL
XFILL_3__1677_ vdd gnd FILL
XFILL_1__868_ vdd gnd FILL
XFILL_4__1022_ vdd gnd FILL
X_1059_ _999_/Y _982_/A _1059_/C _1060_/B vdd gnd OAI21X1
X_1128_ _1390_/B _957_/A _1128_/C _1130_/C vdd gnd OAI21X1
XFILL_1__1313_ vdd gnd FILL
XFILL_1__1175_ vdd gnd FILL
XFILL_1__1244_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_2__1353_ vdd gnd FILL
XFILL_2__1284_ vdd gnd FILL
XFILL_1_CLKBUF1_insert5 vdd gnd FILL
XFILL_0__886_ vdd gnd FILL
X_908_ _982_/A _986_/A _990_/A _925_/C vdd gnd NAND3X1
XFILL_3__1531_ vdd gnd FILL
XFILL_3__1600_ vdd gnd FILL
X_839_ _839_/A _852_/A _895_/B _850_/A vdd gnd OAI21X1
XFILL_3__1462_ vdd gnd FILL
XFILL_3__1393_ vdd gnd FILL
XFILL_4__864_ vdd gnd FILL
XFILL_0__1049_ vdd gnd FILL
X_1677_ _1677_/A _1677_/B _1677_/C _1710_/D vdd gnd OAI21X1
XFILL_4__1640_ vdd gnd FILL
XFILL_0__1118_ vdd gnd FILL
XFILL_4__1571_ vdd gnd FILL
XFILL_4__1005_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_3__882_ vdd gnd FILL
XFILL_2__1405_ vdd gnd FILL
XFILL103050x39150 vdd gnd FILL
XFILL_2__1198_ vdd gnd FILL
XFILL_2__1336_ vdd gnd FILL
XFILL_2__1267_ vdd gnd FILL
XFILL_0__869_ vdd gnd FILL
X_1531_ _952_/Q _975_/A _1532_/C vdd gnd NOR2X1
X_1600_ _1602_/C _1600_/B _1600_/C _1601_/A vdd gnd NAND3X1
X_1462_ _1490_/A _1462_/B _1489_/B _1488_/B vdd gnd AOI21X1
XFILL_3__1514_ vdd gnd FILL
XFILL_3__1445_ vdd gnd FILL
X_1393_ _1426_/B _1426_/A _1427_/B _1394_/B vdd gnd NAND3X1
XFILL_4__916_ vdd gnd FILL
XFILL_3__1376_ vdd gnd FILL
XFILL_0__1598_ vdd gnd FILL
XFILL_0__1667_ vdd gnd FILL
XFILL_1__1012_ vdd gnd FILL
XFILL_4__847_ vdd gnd FILL
XFILL_4__1623_ vdd gnd FILL
XFILL_4__1554_ vdd gnd FILL
XFILL_4__1485_ vdd gnd FILL
XFILL_2__1052_ vdd gnd FILL
XFILL_2__1121_ vdd gnd FILL
XFILL_3__934_ vdd gnd FILL
XFILL_3__865_ vdd gnd FILL
XFILL_3__1161_ vdd gnd FILL
XFILL_2__1319_ vdd gnd FILL
XFILL_3__1230_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_0__1452_ vdd gnd FILL
XFILL_3__1092_ vdd gnd FILL
XFILL_0__1521_ vdd gnd FILL
X_1514_ _1514_/A _1514_/B _1515_/B vdd gnd NOR2X1
X_1445_ _957_/A _960_/A _1509_/C vdd gnd NOR2X1
X_1376_ _1691_/Q _1376_/B _1381_/A vdd gnd NAND2X1
XFILL_4__1270_ vdd gnd FILL
XFILL_3__1428_ vdd gnd FILL
XFILL_1__1561_ vdd gnd FILL
XFILL_0__1719_ vdd gnd FILL
XFILL_1__1492_ vdd gnd FILL
XFILL_1__1630_ vdd gnd FILL
XFILL_3__1359_ vdd gnd FILL
XFILL_2__883_ vdd gnd FILL
XFILL_2__1670_ vdd gnd FILL
XFILL_4__1537_ vdd gnd FILL
XFILL_4__1468_ vdd gnd FILL
XFILL_4__1399_ vdd gnd FILL
XFILL_2__1035_ vdd gnd FILL
XFILL_2__1104_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
X_1161_ _951_/Q _1359_/B _1177_/A vdd gnd NAND2X1
XFILL_3__917_ vdd gnd FILL
X_1230_ _1230_/A _1235_/C _1230_/C _1237_/B vdd gnd AOI21X1
XFILL_3__848_ vdd gnd FILL
X_1092_ _961_/A _1293_/B vdd gnd INVX2
XFILL_3__1213_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_3__1144_ vdd gnd FILL
XFILL_3__1075_ vdd gnd FILL
XFILL_0__1435_ vdd gnd FILL
XFILL_0__1504_ vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
XFILL_1__1613_ vdd gnd FILL
X_1428_ _1428_/A _1428_/B _1428_/C _1429_/C vdd gnd NOR3X1
XFILL_4__1184_ vdd gnd FILL
XFILL_4__1322_ vdd gnd FILL
X_1359_ _998_/A _1359_/B _1361_/B vdd gnd NAND2X1
XFILL_4__1253_ vdd gnd FILL
XFILL_1__1475_ vdd gnd FILL
XFILL_1__1544_ vdd gnd FILL
XFILL_2__935_ vdd gnd FILL
XFILL_2__866_ vdd gnd FILL
XFILL_2__1722_ vdd gnd FILL
X_941_ _941_/D vdd _948_/R _949_/CLK _958_/A vdd gnd DFFSR
X_872_ _885_/A _885_/C _935_/A _873_/C vdd gnd OAI21X1
XFILL_2__1653_ vdd gnd FILL
XFILL_2__1584_ vdd gnd FILL
XFILL_0__1220_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL_2__1018_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
X_1213_ _1695_/Q _1213_/B _1214_/B vdd gnd NOR2X1
X_1144_ _1691_/Q _1690_/Q _1338_/A vdd gnd NOR2X1
X_1075_ _856_/Y _967_/Y _1075_/C _1307_/B vdd gnd NAND3X1
XFILL_1__884_ vdd gnd FILL
XFILL_1__1260_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_3__1058_ vdd gnd FILL
XFILL_3__1127_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_4__1305_ vdd gnd FILL
XFILL_1__1527_ vdd gnd FILL
XFILL_4__1236_ vdd gnd FILL
XFILL_4__1167_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_1__1458_ vdd gnd FILL
XFILL_2__918_ vdd gnd FILL
XFILL_2__849_ vdd gnd FILL
XFILL_4__1098_ vdd gnd FILL
X_924_ _938_/D _931_/B _953_/Q _930_/C vdd gnd OAI21X1
XFILL103950x46950 vdd gnd FILL
X_855_ _895_/B _855_/B _858_/C vdd gnd NAND2X1
XFILL_2__1567_ vdd gnd FILL
XFILL_2__1636_ vdd gnd FILL
XFILL_2__1498_ vdd gnd FILL
XFILL_0__1203_ vdd gnd FILL
XFILL_4__880_ vdd gnd FILL
XFILL_0__1134_ vdd gnd FILL
X_1693_ _1693_/D vdd _1710_/R _1710_/CLK _1693_/Q vdd gnd DFFSR
XFILL_0__1065_ vdd gnd FILL
XFILL_1__936_ vdd gnd FILL
XFILL_1__867_ vdd gnd FILL
XFILL_3__1676_ vdd gnd FILL
X_1058_ _1058_/A _1061_/A _1058_/C _1072_/A vdd gnd AOI21X1
XFILL_1__1243_ vdd gnd FILL
XFILL_4__1021_ vdd gnd FILL
X_1127_ _1682_/Q _959_/A _1297_/A _1128_/C vdd gnd OAI21X1
XFILL_1__1312_ vdd gnd FILL
XFILL_1__1174_ vdd gnd FILL
XFILL_2__1352_ vdd gnd FILL
XFILL_2__1421_ vdd gnd FILL
XFILL_4__1219_ vdd gnd FILL
XFILL_1_CLKBUF1_insert6 vdd gnd FILL
XFILL_2__1283_ vdd gnd FILL
XFILL103950x58650 vdd gnd FILL
XFILL_0__885_ vdd gnd FILL
X_907_ _938_/D _931_/B _990_/A _911_/C vdd gnd OAI21X1
X_838_ _964_/A _895_/B vdd gnd INVX1
XFILL_3__1530_ vdd gnd FILL
XFILL_3__1461_ vdd gnd FILL
XFILL_4__932_ vdd gnd FILL
XFILL_3__1392_ vdd gnd FILL
XFILL_2__1619_ vdd gnd FILL
XFILL_4__863_ vdd gnd FILL
XFILL_0__1117_ vdd gnd FILL
XFILL_0__1048_ vdd gnd FILL
XFILL_4__1570_ vdd gnd FILL
X_1676_ _1676_/A _1677_/B _1677_/C _1709_/D vdd gnd OAI21X1
XFILL_1__919_ vdd gnd FILL
XFILL_3__1659_ vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_4__1004_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_3__881_ vdd gnd FILL
XFILL_2__1404_ vdd gnd FILL
XFILL_2__1335_ vdd gnd FILL
XFILL_2__1197_ vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
XFILL_2__1266_ vdd gnd FILL
XFILL_0__868_ vdd gnd FILL
X_1530_ _1530_/A _965_/C _1530_/C _1533_/A vdd gnd NAND3X1
X_1461_ _1520_/A _1473_/B _1461_/C _1490_/A vdd gnd OAI21X1
X_1392_ _1392_/A _1392_/B _1426_/B vdd gnd AND2X2
XFILL_3__1513_ vdd gnd FILL
XFILL_3__1444_ vdd gnd FILL
XFILL_0__1666_ vdd gnd FILL
XFILL_4__915_ vdd gnd FILL
XFILL_3__1375_ vdd gnd FILL
XFILL_4__846_ vdd gnd FILL
XFILL_0__1597_ vdd gnd FILL
XFILL102450x85950 vdd gnd FILL
XFILL_1__1011_ vdd gnd FILL
XFILL_4__1622_ vdd gnd FILL
XFILL_4__1484_ vdd gnd FILL
X_1659_ _1659_/A _1666_/C _1666_/A vdd gnd NAND2X1
XFILL_4__1553_ vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_2__1051_ vdd gnd FILL
XFILL_2__1120_ vdd gnd FILL
XFILL_3__933_ vdd gnd FILL
XFILL_3__864_ vdd gnd FILL
XFILL_0__1520_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_3__1160_ vdd gnd FILL
XFILL_2__1249_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
XFILL_3__1091_ vdd gnd FILL
XFILL102750x62550 vdd gnd FILL
X_1375_ _1559_/A _995_/B _1382_/B vdd gnd NAND2X1
X_1513_ _1513_/A _982_/A _1513_/C _1514_/B vdd gnd NAND3X1
X_1444_ _965_/A _958_/A _1513_/C vdd gnd NOR2X1
XFILL_0__1718_ vdd gnd FILL
XFILL_3__1358_ vdd gnd FILL
XFILL_0__1649_ vdd gnd FILL
XFILL_1__1560_ vdd gnd FILL
XFILL_1__1491_ vdd gnd FILL
XFILL_3__1427_ vdd gnd FILL
XFILL_4__829_ vdd gnd FILL
XFILL_2__882_ vdd gnd FILL
XFILL_3__1289_ vdd gnd FILL
XFILL_4__1605_ vdd gnd FILL
XFILL_4__1467_ vdd gnd FILL
XFILL_4__1536_ vdd gnd FILL
XFILL_4__1398_ vdd gnd FILL
XFILL_2__1103_ vdd gnd FILL
XFILL_2__1034_ vdd gnd FILL
XFILL_3__916_ vdd gnd FILL
XFILL_3__1212_ vdd gnd FILL
X_1160_ _1330_/B _1330_/C _1359_/B vdd gnd NAND2X1
XFILL_3__847_ vdd gnd FILL
XFILL_0__1503_ vdd gnd FILL
X_1091_ _961_/A _1394_/A _1099_/A vdd gnd NAND2X1
XFILL_0__1365_ vdd gnd FILL
XFILL_3__1074_ vdd gnd FILL
XFILL_3__1143_ vdd gnd FILL
XFILL_0__1434_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
X_1358_ _1358_/A _1358_/B _1358_/C _1367_/A vdd gnd NAND3X1
XFILL_4__1321_ vdd gnd FILL
XFILL_1__1612_ vdd gnd FILL
XFILL_1_BUFX2_insert11 vdd gnd FILL
X_1427_ _1427_/A _1427_/B _1427_/C _1428_/C vdd gnd NAND3X1
XFILL_4__1183_ vdd gnd FILL
XFILL_4__1252_ vdd gnd FILL
XFILL_1__1474_ vdd gnd FILL
XFILL_1__1543_ vdd gnd FILL
X_1289_ _1289_/A _1289_/B _1289_/C _1290_/C vdd gnd OAI21X1
XFILL_2__934_ vdd gnd FILL
XFILL_2__865_ vdd gnd FILL
X_940_ _940_/D vdd _948_/R _949_/CLK _957_/A vdd gnd DFFSR
X_871_ _958_/A _885_/A vdd gnd INVX2
XFILL_2__1652_ vdd gnd FILL
XFILL_2__1721_ vdd gnd FILL
XFILL_2__1583_ vdd gnd FILL
XFILL_4__1519_ vdd gnd FILL
XFILL_0__1150_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
X_1212_ _953_/Q _1403_/B _1226_/C vdd gnd NOR2X1
XFILL_1__883_ vdd gnd FILL
X_1074_ _1074_/A _1074_/B _1080_/D _1075_/C vdd gnd OAI21X1
X_1143_ _1692_/Q _1559_/A vdd gnd INVX1
XFILL_0__1417_ vdd gnd FILL
XFILL_0__1348_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_3__1057_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_3__1126_ vdd gnd FILL
XFILL_1__1526_ vdd gnd FILL
XFILL_4__1304_ vdd gnd FILL
XFILL_4__1166_ vdd gnd FILL
XFILL_2__917_ vdd gnd FILL
XFILL_4__1235_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_4__1097_ vdd gnd FILL
XFILL_1__1457_ vdd gnd FILL
XFILL_2__848_ vdd gnd FILL
X_923_ _935_/A _923_/B _923_/C _952_/D vdd gnd OAI21X1
X_854_ _864_/B _854_/B _855_/B vdd gnd NOR2X1
XFILL_2__1635_ vdd gnd FILL
XFILL_2__1566_ vdd gnd FILL
XFILL_2__1497_ vdd gnd FILL
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
X_1692_ _1692_/D vdd _1708_/R _1709_/CLK _1692_/Q vdd gnd DFFSR
XFILL_1__935_ vdd gnd FILL
XFILL_1__866_ vdd gnd FILL
X_1126_ _960_/A _1390_/A _1297_/A vdd gnd NOR2X1
XFILL_3__1675_ vdd gnd FILL
X_1057_ _1057_/A _1057_/B _1057_/C _1058_/C vdd gnd OAI21X1
XFILL_1__1173_ vdd gnd FILL
XFILL_1__1242_ vdd gnd FILL
XFILL_4__1020_ vdd gnd FILL
XFILL_3__1109_ vdd gnd FILL
XFILL_1__1311_ vdd gnd FILL
XFILL_4__1218_ vdd gnd FILL
XFILL_2__1351_ vdd gnd FILL
XFILL_2__1420_ vdd gnd FILL
XFILL_1__1509_ vdd gnd FILL
XFILL_2__1282_ vdd gnd FILL
XFILL_4__1149_ vdd gnd FILL
XFILL_0__884_ vdd gnd FILL
XFILL_1_CLKBUF1_insert7 vdd gnd FILL
X_837_ _937_/A _853_/A _858_/B vdd gnd NAND2X1
X_906_ _935_/A _906_/B _906_/C _949_/D vdd gnd OAI21X1
XFILL_2__1618_ vdd gnd FILL
XFILL_3__1391_ vdd gnd FILL
XFILL_3__1460_ vdd gnd FILL
XFILL_4__931_ vdd gnd FILL
XFILL_4__862_ vdd gnd FILL
XFILL_2__1549_ vdd gnd FILL
XFILL_0__1047_ vdd gnd FILL
XFILL_0__1116_ vdd gnd FILL
X_1675_ _1675_/A _1675_/B _1708_/D vdd gnd NAND2X1
XFILL_1__918_ vdd gnd FILL
XFILL_1__849_ vdd gnd FILL
XFILL_3__1589_ vdd gnd FILL
X_1109_ _1109_/A _1109_/B _1110_/B vdd gnd NAND2X1
XFILL_3__1658_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1156_ vdd gnd FILL
XFILL_4__1003_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL_3__880_ vdd gnd FILL
XFILL_2__1334_ vdd gnd FILL
XFILL_2__1403_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL103950x7950 vdd gnd FILL
XFILL_2__1196_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
XFILL_0__867_ vdd gnd FILL
X_1391_ _1684_/Q _1537_/A _1392_/B vdd gnd NOR2X1
X_1460_ _1492_/B _1492_/A _1461_/C vdd gnd NAND2X1
XFILL_3__1512_ vdd gnd FILL
XFILL_3__1374_ vdd gnd FILL
XFILL_0__1596_ vdd gnd FILL
XFILL_3__1443_ vdd gnd FILL
XFILL_0__1665_ vdd gnd FILL
XFILL_4__914_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
XFILL_4__845_ vdd gnd FILL
XFILL_4__1621_ vdd gnd FILL
X_1658_ _979_/B _1672_/B _1666_/C vdd gnd NAND2X1
X_1589_ _1695_/Q _1694_/Q _1710_/Q _1590_/A vdd gnd OAI21X1
XFILL_4__1552_ vdd gnd FILL
XFILL_4__1483_ vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_2__1050_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_3__932_ vdd gnd FILL
XFILL_3__863_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_2__1317_ vdd gnd FILL
XFILL_2__1248_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
XFILL_3__1090_ vdd gnd FILL
XFILL_0__919_ vdd gnd FILL
XFILL_2__1179_ vdd gnd FILL
X_1512_ _987_/B _1512_/B _1514_/A vdd gnd NAND2X1
X_1374_ _1573_/A _1374_/B _1374_/C _1382_/A vdd gnd NAND3X1
X_1443_ _966_/A _1534_/A vdd gnd INVX1
XFILL_3__1357_ vdd gnd FILL
XFILL_0__1648_ vdd gnd FILL
XFILL_0__1579_ vdd gnd FILL
XFILL_3__1288_ vdd gnd FILL
XFILL_0__1717_ vdd gnd FILL
XFILL_1__1490_ vdd gnd FILL
XFILL_3__1426_ vdd gnd FILL
XFILL_4__828_ vdd gnd FILL
XFILL_2__881_ vdd gnd FILL
XFILL_4__1604_ vdd gnd FILL
XFILL_4__1535_ vdd gnd FILL
XFILL_4__1397_ vdd gnd FILL
XFILL_4__1466_ vdd gnd FILL
XFILL_2__1033_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_3__915_ vdd gnd FILL
XFILL_3__846_ vdd gnd FILL
XFILL_3__1211_ vdd gnd FILL
XFILL_3__1142_ vdd gnd FILL
XFILL_0__1433_ vdd gnd FILL
X_1090_ _1121_/B _1544_/A _1394_/A vdd gnd XOR2X1
XFILL_0__1502_ vdd gnd FILL
XFILL_0__1364_ vdd gnd FILL
XFILL_3__1073_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
X_1357_ _1415_/B _1415_/A _1357_/C _1430_/B vdd gnd NAND3X1
XFILL_4__1320_ vdd gnd FILL
XFILL_4__1251_ vdd gnd FILL
XFILL_1_BUFX2_insert12 vdd gnd FILL
X_1288_ _1288_/A _1297_/B _1288_/C _1290_/B vdd gnd OAI21X1
XFILL_1__1542_ vdd gnd FILL
XFILL_1__1611_ vdd gnd FILL
X_1426_ _1426_/A _1426_/B _1427_/C vdd gnd AND2X2
XFILL_4__1182_ vdd gnd FILL
XFILL_2__933_ vdd gnd FILL
XFILL_3__1409_ vdd gnd FILL
XFILL_1__1473_ vdd gnd FILL
XFILL_2__864_ vdd gnd FILL
XFILL_2__1720_ vdd gnd FILL
X_870_ _870_/A _937_/B _940_/D vdd gnd NOR2X1
XFILL_2__1651_ vdd gnd FILL
XFILL_4__1518_ vdd gnd FILL
XFILL_4__1449_ vdd gnd FILL
XFILL_2__1582_ vdd gnd FILL
XFILL_2__1016_ vdd gnd FILL
XFILL_0__1080_ vdd gnd FILL
XFILL_3__829_ vdd gnd FILL
X_1211_ _1211_/A _1211_/B _1211_/C _1230_/A vdd gnd OAI21X1
X_1142_ _1693_/Q _1573_/A vdd gnd INVX2
X_999_ _999_/A _999_/Y vdd gnd INVX2
XFILL_1__882_ vdd gnd FILL
XFILL_0__1416_ vdd gnd FILL
X_1073_ _956_/Q _1618_/B _1073_/C _1080_/D vdd gnd AOI21X1
XFILL_3__1125_ vdd gnd FILL
XFILL_0__1347_ vdd gnd FILL
XFILL_3__1056_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
X_1409_ _1679_/Q _1433_/A vdd gnd INVX1
XFILL_1__1525_ vdd gnd FILL
XFILL_4__1234_ vdd gnd FILL
XFILL_4__1303_ vdd gnd FILL
XFILL_2__916_ vdd gnd FILL
XFILL_4__1165_ vdd gnd FILL
XFILL_1__1387_ vdd gnd FILL
XFILL_4__1096_ vdd gnd FILL
XFILL_1__1456_ vdd gnd FILL
XFILL_2__847_ vdd gnd FILL
X_853_ _853_/A _853_/B _853_/Y vdd gnd NOR2X1
X_922_ _933_/B _922_/B _934_/A _923_/B vdd gnd NAND3X1
XFILL_2__1565_ vdd gnd FILL
XFILL_2__1634_ vdd gnd FILL
XFILL_0__1201_ vdd gnd FILL
XFILL_2__1496_ vdd gnd FILL
XFILL_0__1063_ vdd gnd FILL
XFILL_0__1132_ vdd gnd FILL
X_1691_ _1691_/D vdd _1708_/R _1709_/CLK _1691_/Q vdd gnd DFFSR
XFILL_1__934_ vdd gnd FILL
XFILL_3__1674_ vdd gnd FILL
XFILL_1__865_ vdd gnd FILL
X_1125_ _1125_/A _1133_/A _1134_/B vdd gnd NAND2X1
XFILL_1__1310_ vdd gnd FILL
X_1056_ _1056_/A _1056_/B _1056_/C _1057_/C vdd gnd AOI21X1
XFILL_1__1172_ vdd gnd FILL
XFILL_1__1241_ vdd gnd FILL
XFILL_3__1108_ vdd gnd FILL
XFILL_3__1039_ vdd gnd FILL
XFILL_4__1217_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_2__1281_ vdd gnd FILL
XFILL_1__1508_ vdd gnd FILL
XFILL_4__1148_ vdd gnd FILL
XFILL_1_CLKBUF1_insert8 vdd gnd FILL
XFILL_0__883_ vdd gnd FILL
X_905_ _938_/D _931_/B _986_/A _906_/C vdd gnd OAI21X1
X_836_ _975_/A _968_/A _852_/A _839_/A _853_/A vdd gnd OAI22X1
XFILL_2__1617_ vdd gnd FILL
XFILL_3__1390_ vdd gnd FILL
XFILL_2__1548_ vdd gnd FILL
XFILL_4__930_ vdd gnd FILL
XFILL_4__861_ vdd gnd FILL
XFILL_2__1479_ vdd gnd FILL
XFILL_0__1046_ vdd gnd FILL
X_1674_ _1674_/A _1674_/B _1674_/C _1707_/D vdd gnd AOI21X1
XFILL_0__1115_ vdd gnd FILL
XFILL_1__917_ vdd gnd FILL
XFILL_3__1657_ vdd gnd FILL
X_1039_ _952_/Q _1650_/A _1043_/B vdd gnd NAND2X1
XFILL_4__1002_ vdd gnd FILL
XFILL_1__848_ vdd gnd FILL
XFILL_3__1588_ vdd gnd FILL
X_1108_ _1135_/B _962_/B _1136_/C vdd gnd OR2X2
XFILL_1__1224_ vdd gnd FILL
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1086_ vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_2__1195_ vdd gnd FILL
XFILL_2__1333_ vdd gnd FILL
XFILL_2__1264_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
XFILL_0__866_ vdd gnd FILL
XFILL_3__1511_ vdd gnd FILL
X_1390_ _1390_/A _1390_/B _1520_/A _1392_/A vdd gnd OAI21X1
XFILL_3__1442_ vdd gnd FILL
XFILL_3__1373_ vdd gnd FILL
XFILL_0__1595_ vdd gnd FILL
XFILL_0__1664_ vdd gnd FILL
XFILL_4__913_ vdd gnd FILL
XFILL_4__844_ vdd gnd FILL
XFILL_0__1029_ vdd gnd FILL
X_1588_ _1588_/A _1597_/A vdd gnd INVX1
X_1657_ _1657_/A _1657_/B _1663_/A _1659_/A vdd gnd OAI21X1
XFILL_4__1620_ vdd gnd FILL
XFILL_4__1551_ vdd gnd FILL
XFILL_4__1482_ vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_3__931_ vdd gnd FILL
XFILL_3__862_ vdd gnd FILL
XFILL103050x11850 vdd gnd FILL
XFILL_2__1178_ vdd gnd FILL
XFILL_2__1316_ vdd gnd FILL
XFILL_2__1247_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
XFILL_0__918_ vdd gnd FILL
XFILL_0__849_ vdd gnd FILL
X_1442_ _1513_/A _1442_/B _1442_/C _1582_/B vdd gnd NAND3X1
X_1511_ _1511_/A _1511_/B _1516_/A vdd gnd OR2X2
XFILL_0__1716_ vdd gnd FILL
XFILL_3__1425_ vdd gnd FILL
X_1373_ _1696_/Q _1616_/B _1697_/Q _1388_/B _1389_/A vdd gnd OAI22X1
XFILL_3__1356_ vdd gnd FILL
XFILL_2__880_ vdd gnd FILL
XFILL_0__1647_ vdd gnd FILL
XFILL_0__1578_ vdd gnd FILL
XFILL_3__1287_ vdd gnd FILL
XFILL_4__1603_ vdd gnd FILL
XFILL_4__1534_ vdd gnd FILL
X_1709_ _1709_/D _1709_/S vdd _1709_/CLK _1709_/Q vdd gnd DFFSR
XFILL_4__1396_ vdd gnd FILL
XFILL_4__1465_ vdd gnd FILL
XFILL_2__1032_ vdd gnd FILL
XFILL_2__1101_ vdd gnd FILL
XFILL_3__914_ vdd gnd FILL
XFILL_3__845_ vdd gnd FILL
XFILL_3__1210_ vdd gnd FILL
XFILL103650x70350 vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_3__1141_ vdd gnd FILL
XFILL_0__1501_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XFILL_3__1072_ vdd gnd FILL
XFILL_0__1294_ vdd gnd FILL
X_1425_ _1425_/A _1425_/B _1425_/C _1429_/B vdd gnd AOI21X1
XFILL_1_BUFX2_insert13 vdd gnd FILL
X_1356_ _1356_/A _1356_/B _1415_/A vdd gnd AND2X2
XFILL_4__1181_ vdd gnd FILL
XFILL_4__1250_ vdd gnd FILL
XFILL_1__1610_ vdd gnd FILL
XFILL_1__1472_ vdd gnd FILL
XFILL_1__1541_ vdd gnd FILL
XFILL_3__1408_ vdd gnd FILL
X_1287_ _1287_/A _1289_/B _1298_/C vdd gnd NOR2X1
XFILL_2__932_ vdd gnd FILL
XFILL_2__863_ vdd gnd FILL
XFILL_3__1339_ vdd gnd FILL
XFILL_2__1650_ vdd gnd FILL
XFILL_2__1581_ vdd gnd FILL
XFILL_4__1517_ vdd gnd FILL
XFILL_4__1379_ vdd gnd FILL
XFILL_4__1448_ vdd gnd FILL
XFILL_2__1015_ vdd gnd FILL
XFILL103050x35250 vdd gnd FILL
XFILL_3__828_ vdd gnd FILL
X_1210_ _1210_/A _1248_/A _1210_/C _1211_/C vdd gnd AOI21X1
X_1141_ _1698_/Q _1605_/B vdd gnd INVX2
X_1072_ _1072_/A _1072_/B _1072_/C _1073_/C vdd gnd OAI21X1
XFILL_1__881_ vdd gnd FILL
X_998_ _998_/A _998_/Y vdd gnd INVX2
XFILL_0__1346_ vdd gnd FILL
XFILL_0__1415_ vdd gnd FILL
XFILL_3__1055_ vdd gnd FILL
XFILL_3__1124_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1677_/B _1408_/B _1408_/C _1678_/D vdd gnd OAI21X1
XFILL_4__1164_ vdd gnd FILL
XFILL_4__1233_ vdd gnd FILL
X_1339_ _1364_/A _1341_/B vdd gnd INVX1
XFILL_1__1524_ vdd gnd FILL
XFILL_1__1455_ vdd gnd FILL
XFILL_4__1302_ vdd gnd FILL
XFILL_2__915_ vdd gnd FILL
XFILL_1__1386_ vdd gnd FILL
XFILL_2__846_ vdd gnd FILL
XFILL_4__1095_ vdd gnd FILL
X_921_ _925_/A _925_/C _928_/A _922_/B vdd gnd OAI21X1
X_852_ _852_/A _852_/B _853_/B vdd gnd OR2X2
XFILL_2__1564_ vdd gnd FILL
XFILL_2__1633_ vdd gnd FILL
XFILL_0__1200_ vdd gnd FILL
XFILL_2__1495_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
X_1690_ _1690_/D vdd _1710_/R _1710_/CLK _1690_/Q vdd gnd DFFSR
XFILL_0__1131_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
XFILL_3__1673_ vdd gnd FILL
X_1055_ _1055_/A _1055_/B _1055_/C _1057_/A vdd gnd AOI21X1
XFILL_1__864_ vdd gnd FILL
X_1124_ _1523_/A _1520_/A _1124_/C _1125_/A vdd gnd NAND3X1
XFILL_0__1329_ vdd gnd FILL
XFILL_3__1038_ vdd gnd FILL
XFILL_1__1171_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
XFILL_3__1107_ vdd gnd FILL
XFILL_4__1216_ vdd gnd FILL
XFILL_4__1147_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
XFILL_2__1280_ vdd gnd FILL
XFILL_1__1507_ vdd gnd FILL
XFILL_2__829_ vdd gnd FILL
XFILL_4__1078_ vdd gnd FILL
XFILL_0__882_ vdd gnd FILL
XFILL_1_CLKBUF1_insert9 vdd gnd FILL
X_904_ _904_/A _915_/B _934_/A _906_/B vdd gnd NAND3X1
X_835_ _925_/A _915_/A _902_/A _839_/A vdd gnd NAND3X1
XFILL_2__1616_ vdd gnd FILL
XFILL_2__1547_ vdd gnd FILL
XFILL_2__1478_ vdd gnd FILL
XFILL_4__860_ vdd gnd FILL
XFILL_0__1114_ vdd gnd FILL
XFILL_0__1045_ vdd gnd FILL
X_1673_ _1673_/A _1673_/B _1673_/C _1674_/A vdd gnd OAI21X1
XFILL_1__916_ vdd gnd FILL
XFILL_3__1725_ vdd gnd FILL
XFILL_1__847_ vdd gnd FILL
XFILL_3__1587_ vdd gnd FILL
XFILL_3__1656_ vdd gnd FILL
XFILL_1__1223_ vdd gnd FILL
X_1038_ _953_/Q _1655_/A _1055_/B vdd gnd NAND2X1
XFILL_4__1001_ vdd gnd FILL
X_1107_ _1107_/A _1537_/A _1135_/B vdd gnd XOR2X1
XFILL_4__989_ vdd gnd FILL
XFILL_1__1154_ vdd gnd FILL
XFILL_1__1085_ vdd gnd FILL
XFILL_2__1401_ vdd gnd FILL
XFILL_2__1332_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_2__1194_ vdd gnd FILL
XFILL_2__1263_ vdd gnd FILL
XFILL_0__865_ vdd gnd FILL
XFILL_3__1441_ vdd gnd FILL
XFILL_3__1510_ vdd gnd FILL
XFILL_4__912_ vdd gnd FILL
XFILL_3__1372_ vdd gnd FILL
XFILL_0__1594_ vdd gnd FILL
XFILL_0__1663_ vdd gnd FILL
X_1725_ _853_/Y vsync vdd gnd BUFX2
XFILL_4__843_ vdd gnd FILL
XFILL_0__1028_ vdd gnd FILL
X_1587_ _1696_/Q _1710_/Q _1588_/A vdd gnd XOR2X1
X_1656_ _1656_/A _1656_/B _1656_/C _1673_/A vdd gnd AOI21X1
XFILL_4__1550_ vdd gnd FILL
XFILL_3__1639_ vdd gnd FILL
XFILL_4__1481_ vdd gnd FILL
XFILL_1__1206_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_3__930_ vdd gnd FILL
XFILL_3__861_ vdd gnd FILL
XFILL_2__1315_ vdd gnd FILL
XFILL_2__1177_ vdd gnd FILL
XFILL_0__917_ vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
X_1441_ _1441_/A _1441_/B _1442_/B vdd gnd NOR2X1
X_1510_ _997_/B _981_/A _1510_/C _1511_/B vdd gnd NAND3X1
XFILL_0__848_ vdd gnd FILL
XFILL_3__1424_ vdd gnd FILL
X_1372_ _980_/B _980_/A _1388_/B vdd gnd OR2X2
XFILL_0__1715_ vdd gnd FILL
XFILL_0__1646_ vdd gnd FILL
XFILL_3__1355_ vdd gnd FILL
XFILL_0__1577_ vdd gnd FILL
XFILL_3__1286_ vdd gnd FILL
X_1708_ _1708_/D vdd _1708_/R _1709_/CLK _1708_/Q vdd gnd DFFSR
XFILL_4__1602_ vdd gnd FILL
XFILL_4__1533_ vdd gnd FILL
XFILL_4__1464_ vdd gnd FILL
X_1639_ _1639_/A _1645_/B _1640_/A vdd gnd XNOR2X1
XFILL_4__1395_ vdd gnd FILL
XFILL_2__1031_ vdd gnd FILL
XFILL_2__1100_ vdd gnd FILL
XFILL_3__913_ vdd gnd FILL
XFILL_3_BUFX2_insert0 vdd gnd FILL
XFILL103950x54750 vdd gnd FILL
XFILL_3__844_ vdd gnd FILL
XFILL_0__1500_ vdd gnd FILL
XFILL103650x89850 vdd gnd FILL
XFILL_2__1229_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
XFILL_3__1140_ vdd gnd FILL
XFILL_3__1071_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
X_1355_ _979_/B _1355_/B _1355_/C _1356_/A vdd gnd NAND3X1
X_1424_ _1604_/A _981_/B _1605_/B _1424_/D _1425_/C vdd gnd OAI22X1
XFILL_1_BUFX2_insert14 vdd gnd FILL
XFILL_3__1338_ vdd gnd FILL
XFILL_4__1180_ vdd gnd FILL
XFILL_3__1407_ vdd gnd FILL
XFILL_1__1471_ vdd gnd FILL
XFILL_1__1540_ vdd gnd FILL
XFILL_0__1629_ vdd gnd FILL
X_1286_ _1286_/A _1289_/C _1289_/B vdd gnd NAND2X1
XFILL_2__931_ vdd gnd FILL
XFILL_2__862_ vdd gnd FILL
XFILL_3__1269_ vdd gnd FILL
XFILL_4__1516_ vdd gnd FILL
XFILL_4__1447_ vdd gnd FILL
XFILL_2__1580_ vdd gnd FILL
XFILL_4__1378_ vdd gnd FILL
XFILL_1__1669_ vdd gnd FILL
XFILL_2__1014_ vdd gnd FILL
XFILL103350x19650 vdd gnd FILL
XFILL103950x66450 vdd gnd FILL
X_997_ _997_/A _997_/B _997_/Y vdd gnd NAND2X1
XFILL_1__880_ vdd gnd FILL
X_1140_ _1697_/Q _1604_/A vdd gnd INVX2
X_1071_ _959_/A _959_/B _1071_/C _1072_/C vdd gnd AOI21X1
XFILL_0__1414_ vdd gnd FILL
XFILL_0__1345_ vdd gnd FILL
XFILL_3__1054_ vdd gnd FILL
XFILL_0__1276_ vdd gnd FILL
XFILL_3__1123_ vdd gnd FILL
X_1338_ _1338_/A _1338_/B _984_/B _1364_/A vdd gnd OAI21X1
X_1407_ _1407_/A _1677_/C _1677_/B vdd gnd NAND2X1
XFILL_4__1301_ vdd gnd FILL
XFILL_4__1163_ vdd gnd FILL
XFILL_4__1232_ vdd gnd FILL
XFILL_1__1385_ vdd gnd FILL
X_1269_ _1269_/A _1269_/B _1270_/B vdd gnd NAND2X1
XFILL_1__1454_ vdd gnd FILL
XFILL_4__1094_ vdd gnd FILL
XFILL_1__1523_ vdd gnd FILL
XFILL_2__914_ vdd gnd FILL
XFILL_2__845_ vdd gnd FILL
X_920_ _952_/Q _928_/A vdd gnd INVX1
X_851_ _925_/A _937_/A _852_/B vdd gnd NAND2X1
XFILL_2__1632_ vdd gnd FILL
XFILL_2__1494_ vdd gnd FILL
XFILL_2__1563_ vdd gnd FILL
XFILL_0__1130_ vdd gnd FILL
XFILL_0__1061_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
XFILL_1__863_ vdd gnd FILL
XFILL_3__1672_ vdd gnd FILL
X_1054_ _1060_/A _1054_/B _1054_/C _1058_/A vdd gnd OAI21X1
X_1123_ _1123_/A _1123_/B _1428_/A vdd gnd NAND2X1
XFILL_3__1037_ vdd gnd FILL
XFILL_0__1328_ vdd gnd FILL
XFILL_1__1170_ vdd gnd FILL
XFILL_0__1259_ vdd gnd FILL
XFILL_3__1106_ vdd gnd FILL
XFILL_1__1506_ vdd gnd FILL
XFILL_4__1215_ vdd gnd FILL
XFILL_4__1146_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_4__1077_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_2__828_ vdd gnd FILL
XFILL_0__881_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
X_903_ _982_/A _986_/A _915_/B vdd gnd NAND2X1
X_834_ _982_/A _986_/A _902_/A vdd gnd NOR2X1
XFILL_2__1615_ vdd gnd FILL
XFILL_2__1477_ vdd gnd FILL
XFILL_2__1546_ vdd gnd FILL
XFILL_0__1113_ vdd gnd FILL
XFILL_3__1724_ vdd gnd FILL
XFILL_0__1044_ vdd gnd FILL
X_1672_ _1672_/A _1672_/B _1673_/A _1673_/C vdd gnd NAND3X1
XFILL_1__915_ vdd gnd FILL
XFILL102750x70350 vdd gnd FILL
XFILL_1__846_ vdd gnd FILL
XFILL_3__1655_ vdd gnd FILL
X_1106_ _1281_/B _1426_/A _1112_/C vdd gnd NAND2X1
XFILL_3__1586_ vdd gnd FILL
XFILL_4__1000_ vdd gnd FILL
X_1037_ _971_/A _1655_/A vdd gnd INVX2
XFILL_1__1153_ vdd gnd FILL
XFILL_4__988_ vdd gnd FILL
XFILL_1__1222_ vdd gnd FILL
XFILL_1__1084_ vdd gnd FILL
XFILL_2__1400_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_2__1262_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_0__864_ vdd gnd FILL
XFILL_4__1129_ vdd gnd FILL
XFILL_3__1440_ vdd gnd FILL
XFILL_3__1371_ vdd gnd FILL
XFILL_0__1662_ vdd gnd FILL
XFILL_4__911_ vdd gnd FILL
XFILL_4__842_ vdd gnd FILL
XFILL_0__1593_ vdd gnd FILL
XFILL_2__1529_ vdd gnd FILL
X_1724_ _1724_/A rgb[9] vdd gnd BUFX2
XFILL_0__1027_ vdd gnd FILL
X_1655_ _1655_/A _1671_/C _1655_/C _1656_/C vdd gnd OAI21X1
XFILL_4__1480_ vdd gnd FILL
X_1586_ _1619_/A _1586_/B _1586_/C _1695_/D vdd gnd OAI21X1
XFILL_1__829_ vdd gnd FILL
XFILL_3__1569_ vdd gnd FILL
XFILL_3__1638_ vdd gnd FILL
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
XFILL_3__860_ vdd gnd FILL
XFILL_2__1245_ vdd gnd FILL
XFILL_2__1314_ vdd gnd FILL
XFILL_2__1176_ vdd gnd FILL
XFILL_0__916_ vdd gnd FILL
XFILL_0__847_ vdd gnd FILL
X_1440_ _982_/A _987_/B _1441_/A vdd gnd NAND2X1
X_1371_ _1429_/A _1398_/B vdd gnd INVX1
XFILL_0__1714_ vdd gnd FILL
XFILL_3__1354_ vdd gnd FILL
XFILL_3__989_ vdd gnd FILL
XFILL_3__1423_ vdd gnd FILL
XFILL_0__1645_ vdd gnd FILL
XFILL_0__1576_ vdd gnd FILL
XFILL_3__1285_ vdd gnd FILL
X_1707_ _1707_/D vdd _1710_/R _1710_/CLK _1707_/Q vdd gnd DFFSR
XFILL_4__1601_ vdd gnd FILL
X_1638_ _1671_/C _998_/Y _1645_/B vdd gnd XOR2X1
XFILL_4__1532_ vdd gnd FILL
X_1569_ _1569_/A _1577_/C vdd gnd INVX1
XFILL_4__1463_ vdd gnd FILL
XFILL_4__1394_ vdd gnd FILL
XFILL_3_BUFX2_insert1 vdd gnd FILL
XFILL_2__1030_ vdd gnd FILL
XFILL_1__1119_ vdd gnd FILL
XFILL_3__912_ vdd gnd FILL
XFILL_3__843_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_2__1228_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
XFILL_3__1070_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_2__1159_ vdd gnd FILL
X_1354_ _1354_/A _1358_/A _1358_/B _1415_/B vdd gnd NAND3X1
X_1423_ _1423_/A _1423_/B _1423_/C _1425_/A vdd gnd OAI21X1
X_1285_ _1684_/Q _1530_/A _1289_/C vdd gnd NAND2X1
XFILL_1_BUFX2_insert15 vdd gnd FILL
XFILL_2__930_ vdd gnd FILL
XFILL_3__1406_ vdd gnd FILL
XFILL_3__1337_ vdd gnd FILL
XFILL_0__1559_ vdd gnd FILL
XFILL_1__1470_ vdd gnd FILL
XFILL_0__1628_ vdd gnd FILL
XFILL_2__861_ vdd gnd FILL
XFILL_3__1199_ vdd gnd FILL
XFILL_3__1268_ vdd gnd FILL
XFILL_4__1377_ vdd gnd FILL
XFILL_4__1446_ vdd gnd FILL
XFILL_4__1515_ vdd gnd FILL
XFILL_1__1668_ vdd gnd FILL
XFILL_1__1599_ vdd gnd FILL
XFILL_2__1013_ vdd gnd FILL
X_996_ _996_/A _996_/B _996_/C _996_/Y vdd gnd AOI21X1
XFILL_0__1413_ vdd gnd FILL
X_1070_ _967_/A _963_/A _1070_/C _1071_/C vdd gnd OAI21X1
XFILL_3__1122_ vdd gnd FILL
XFILL_0__1344_ vdd gnd FILL
XFILL_3__1053_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
XFILL_4__1231_ vdd gnd FILL
X_1406_ _1406_/A _1406_/B _1406_/C _1407_/A vdd gnd NAND3X1
X_1337_ _993_/A _1337_/B _1364_/C vdd gnd NAND2X1
X_1268_ _1268_/A _1268_/B _1269_/A vdd gnd NOR2X1
XFILL_1__1522_ vdd gnd FILL
XFILL_4__1300_ vdd gnd FILL
XFILL_2__913_ vdd gnd FILL
XFILL_4__1162_ vdd gnd FILL
X_1199_ _1692_/Q _997_/B _1248_/B vdd gnd NOR2X1
XFILL_1__1384_ vdd gnd FILL
XFILL_1__1453_ vdd gnd FILL
XFILL_4__1093_ vdd gnd FILL
XFILL_2__844_ vdd gnd FILL
X_850_ _850_/A _858_/B _850_/C _850_/Y vdd gnd NOR3X1
XFILL_2__1631_ vdd gnd FILL
XFILL_4__1429_ vdd gnd FILL
XFILL_2__1493_ vdd gnd FILL
XFILL_2__1562_ vdd gnd FILL
XFILL_0__1060_ vdd gnd FILL
XFILL_2_CLKBUF1_insert4 vdd gnd FILL
XFILL_1__931_ vdd gnd FILL
XFILL_1__862_ vdd gnd FILL
X_979_ _979_/A _979_/B _979_/C _980_/A vdd gnd AOI21X1
XFILL_3__1671_ vdd gnd FILL
X_1122_ _1545_/A _1122_/B _1123_/B vdd gnd NAND2X1
X_1053_ _998_/A _1512_/B _1053_/C _1054_/C vdd gnd AOI21X1
XFILL_3__1105_ vdd gnd FILL
XFILL_0__1327_ vdd gnd FILL
XFILL_0__1189_ vdd gnd FILL
XFILL_3__1036_ vdd gnd FILL
XFILL_0__1258_ vdd gnd FILL
XFILL_4__1214_ vdd gnd FILL
XFILL_1__1505_ vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
XFILL_4__1145_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_0__880_ vdd gnd FILL
XFILL_4__1076_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
X_833_ _990_/A _915_/A vdd gnd INVX1
X_902_ _902_/A _904_/A vdd gnd INVX1
XFILL_2__1614_ vdd gnd FILL
XFILL_2__1545_ vdd gnd FILL
XFILL_2__1476_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
X_1671_ _979_/C _979_/B _1671_/C _1673_/B vdd gnd NAND3X1
XFILL_0__1112_ vdd gnd FILL
XFILL_1__914_ vdd gnd FILL
XFILL_3__1654_ vdd gnd FILL
XFILL_3__1723_ vdd gnd FILL
XFILL_1__845_ vdd gnd FILL
XFILL_3__1585_ vdd gnd FILL
X_1105_ _1109_/B _1109_/A _1426_/A vdd gnd AND2X2
XFILL102750x89850 vdd gnd FILL
XFILL_1__1221_ vdd gnd FILL
XFILL_1__1152_ vdd gnd FILL
X_1036_ _1056_/B _1036_/B _1036_/C _1057_/B vdd gnd NAND3X1
XFILL_4__987_ vdd gnd FILL
XFILL_3__1019_ vdd gnd FILL
XFILL_1__1083_ vdd gnd FILL
XFILL_2__1330_ vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_2__1261_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL_2__1192_ vdd gnd FILL
XFILL_0__863_ vdd gnd FILL
XFILL_4__1059_ vdd gnd FILL
XFILL_4__1128_ vdd gnd FILL
XFILL_2__1528_ vdd gnd FILL
XFILL_3__1370_ vdd gnd FILL
XFILL_0__1592_ vdd gnd FILL
XFILL_0__1661_ vdd gnd FILL
XFILL_4__910_ vdd gnd FILL
XFILL_4__841_ vdd gnd FILL
XFILL_2__1459_ vdd gnd FILL
XFILL_0__1026_ vdd gnd FILL
X_1654_ _1654_/A _1654_/B _1656_/B vdd gnd NOR2X1
X_1723_ _1723_/A rgb[8] vdd gnd BUFX2
XFILL102450x19650 vdd gnd FILL
X_1585_ _1585_/A _1591_/B _1586_/B vdd gnd XNOR2X1
XFILL_3__1637_ vdd gnd FILL
XFILL_1__828_ vdd gnd FILL
X_1019_ _974_/B _1616_/B vdd gnd INVX1
XFILL_3__1568_ vdd gnd FILL
XFILL_3__1499_ vdd gnd FILL
XFILL_1__1204_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_1__1135_ vdd gnd FILL
XFILL_4__1677_ vdd gnd FILL
XFILL_2__1175_ vdd gnd FILL
XFILL_2__1244_ vdd gnd FILL
XFILL_2__1313_ vdd gnd FILL
XFILL_0__915_ vdd gnd FILL
XFILL_0__846_ vdd gnd FILL
XFILL_3__988_ vdd gnd FILL
X_1370_ _1698_/Q _1618_/B _1429_/A vdd gnd NOR2X1
XFILL_0__1713_ vdd gnd FILL
XFILL_3__1353_ vdd gnd FILL
XFILL_3__1422_ vdd gnd FILL
XFILL_0__1575_ vdd gnd FILL
XFILL_3__1284_ vdd gnd FILL
XFILL_0__1644_ vdd gnd FILL
XFILL_0__1009_ vdd gnd FILL
XFILL_4__1600_ vdd gnd FILL
X_1706_ _1706_/D vdd _1709_/S _1709_/CLK _979_/C vdd gnd DFFSR
X_1637_ _992_/A _1671_/C _1637_/C _1639_/A vdd gnd OAI21X1
XFILL_4__1531_ vdd gnd FILL
X_1568_ _1573_/A _1677_/A _1569_/A vdd gnd NOR2X1
X_1499_ _1499_/A _1500_/A _1499_/C _1501_/C vdd gnd OAI21X1
XFILL_4__1393_ vdd gnd FILL
XFILL_3_BUFX2_insert2 vdd gnd FILL
XFILL_1__1049_ vdd gnd FILL
XFILL_1__1118_ vdd gnd FILL
XFILL_3__911_ vdd gnd FILL
XFILL_3__842_ vdd gnd FILL
XFILL_2__1227_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
XFILL_2__1158_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
XFILL_0__829_ vdd gnd FILL
X_1422_ _1422_/A _1695_/Q _1696_/Q _1616_/B _1423_/C vdd gnd AOI22X1
XFILL_2__1089_ vdd gnd FILL
X_1353_ _1655_/A _1353_/B _1353_/C _1354_/A vdd gnd OAI21X1
XFILL_3__1405_ vdd gnd FILL
X_1284_ _965_/A _1523_/A _1286_/A vdd gnd NAND2X1
XFILL_2__860_ vdd gnd FILL
XFILL_3__1336_ vdd gnd FILL
XFILL_3__1267_ vdd gnd FILL
XFILL_0__1558_ vdd gnd FILL
XFILL_0__1489_ vdd gnd FILL
XFILL_0__1627_ vdd gnd FILL
XFILL_3__1198_ vdd gnd FILL
XFILL_4__1514_ vdd gnd FILL
XFILL_4__1376_ vdd gnd FILL
XFILL_4__1445_ vdd gnd FILL
XFILL_1__1598_ vdd gnd FILL
XFILL_1__1667_ vdd gnd FILL
XFILL_2__1012_ vdd gnd FILL
XFILL_2__989_ vdd gnd FILL
X_995_ _997_/B _995_/B _996_/C vdd gnd NOR2X1
XFILL_0__1412_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_3__1121_ vdd gnd FILL
XFILL_3__1052_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
X_1405_ _1694_/Q _1693_/Q _1406_/B vdd gnd NOR2X1
XFILL_4__1161_ vdd gnd FILL
XFILL_4__1230_ vdd gnd FILL
X_1198_ _990_/A _1559_/A _1248_/A vdd gnd NOR2X1
X_1336_ _1338_/A _1338_/B _1337_/B vdd gnd NOR2X1
X_1267_ _1267_/A _1267_/B _1267_/C _1269_/B vdd gnd NAND3X1
XFILL_1__1452_ vdd gnd FILL
XFILL_1__1521_ vdd gnd FILL
XFILL_2__912_ vdd gnd FILL
XFILL_3__1319_ vdd gnd FILL
XFILL_1__1383_ vdd gnd FILL
XFILL_2__843_ vdd gnd FILL
XFILL_4__1092_ vdd gnd FILL
XFILL_2__1561_ vdd gnd FILL
XFILL_2__1630_ vdd gnd FILL
XFILL_4__1359_ vdd gnd FILL
XFILL_2_CLKBUF1_insert5 vdd gnd FILL
XFILL_4__1428_ vdd gnd FILL
XFILL_1__1719_ vdd gnd FILL
XFILL_2__1492_ vdd gnd FILL
XFILL_1__930_ vdd gnd FILL
XFILL_3__1670_ vdd gnd FILL
XCLKBUF1_insert4 clk _1702_/CLK vdd gnd CLKBUF1
XFILL_1__861_ vdd gnd FILL
X_1052_ _998_/Y _951_/Q _997_/Y _1053_/C vdd gnd AOI21X1
X_978_ _978_/A _978_/B _980_/B vdd gnd NOR2X1
X_1121_ _1544_/A _1121_/B _1122_/B vdd gnd NOR2X1
XFILL_0__1326_ vdd gnd FILL
XFILL_3__1035_ vdd gnd FILL
XFILL_3__1104_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
XFILL_0__1257_ vdd gnd FILL
X_1319_ _1347_/B _1347_/A _1414_/A vdd gnd NAND2X1
XFILL_4__1213_ vdd gnd FILL
XFILL_4__1144_ vdd gnd FILL
XFILL_1__1435_ vdd gnd FILL
XFILL_1__1504_ vdd gnd FILL
XFILL_1__1366_ vdd gnd FILL
XFILL_4__1075_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
X_901_ _901_/A _935_/A _901_/C _948_/D vdd gnd AOI21X1
X_832_ _951_/Q _925_/A vdd gnd INVX1
XFILL_2__1613_ vdd gnd FILL
XFILL_2__1544_ vdd gnd FILL
XFILL_2__1475_ vdd gnd FILL
XFILL_0__1042_ vdd gnd FILL
X_1670_ _978_/A _1670_/B _1670_/C _1706_/D vdd gnd OAI21X1
XFILL_0__1111_ vdd gnd FILL
XFILL_1__913_ vdd gnd FILL
XFILL_3__1722_ vdd gnd FILL
XFILL_3__1653_ vdd gnd FILL
XFILL_3__1584_ vdd gnd FILL
X_1035_ _968_/A _1663_/A _1036_/B vdd gnd NAND2X1
XFILL_1__844_ vdd gnd FILL
X_1104_ _1537_/A _1133_/A _1540_/A _1109_/B vdd gnd OAI21X1
XFILL_1__1220_ vdd gnd FILL
XFILL_1__1151_ vdd gnd FILL
XFILL_3__1018_ vdd gnd FILL
XFILL_4__986_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
XFILL_4_CLKBUF1_insert10 vdd gnd FILL
XFILL_0__1309_ vdd gnd FILL
XFILL_0__931_ vdd gnd FILL
XFILL_2__1191_ vdd gnd FILL
XFILL_1__1349_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_2__1260_ vdd gnd FILL
XFILL_0__862_ vdd gnd FILL
XFILL_4__1058_ vdd gnd FILL
XFILL103050x31350 vdd gnd FILL
XFILL_2__1527_ vdd gnd FILL
XFILL_0__1591_ vdd gnd FILL
XFILL_0__1660_ vdd gnd FILL
XFILL_2__1458_ vdd gnd FILL
XFILL_2__1389_ vdd gnd FILL
XFILL_4__840_ vdd gnd FILL
X_1722_ _1724_/A rgb[7] vdd gnd BUFX2
XFILL_0__1025_ vdd gnd FILL
X_1653_ _1653_/A _1655_/A _1670_/B _1704_/D vdd gnd MUX2X1
X_1584_ _1695_/Q _1710_/Q _1591_/B vdd gnd XOR2X1
XFILL_3__1567_ vdd gnd FILL
XFILL_3__1636_ vdd gnd FILL
XFILL_1__1203_ vdd gnd FILL
X_1018_ _1018_/A _1018_/B _1022_/B vdd gnd NAND2X1
XFILL_3__1498_ vdd gnd FILL
XFILL_4__969_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_1__1134_ vdd gnd FILL
XFILL_4__1676_ vdd gnd FILL
XFILL_2__1312_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_0__914_ vdd gnd FILL
XFILL_2__1243_ vdd gnd FILL
XFILL_0__845_ vdd gnd FILL
XFILL103050x43050 vdd gnd FILL
XFILL_0__1712_ vdd gnd FILL
XFILL_3__987_ vdd gnd FILL
XFILL_3__1421_ vdd gnd FILL
XFILL_3__1352_ vdd gnd FILL
XFILL_0__1643_ vdd gnd FILL
XFILL_0__1574_ vdd gnd FILL
XFILL_3__1283_ vdd gnd FILL
X_1705_ _1705_/D vdd _1709_/S _1710_/CLK _979_/B vdd gnd DFFSR
XFILL_0__1008_ vdd gnd FILL
X_1567_ _1577_/A _1570_/A vdd gnd INVX1
XFILL_4__1530_ vdd gnd FILL
X_1636_ _992_/A _1670_/B _1636_/C _1701_/D vdd gnd OAI21X1
X_1498_ _1498_/A _1498_/B _1500_/A vdd gnd NAND2X1
XFILL_4__1461_ vdd gnd FILL
XFILL_4__1392_ vdd gnd FILL
XFILL_3__1619_ vdd gnd FILL
XFILL_1__1048_ vdd gnd FILL
XFILL_3_BUFX2_insert3 vdd gnd FILL
XFILL_1__1117_ vdd gnd FILL
XFILL_3__910_ vdd gnd FILL
XFILL_3__841_ vdd gnd FILL
XFILL_4__1659_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
XFILL_2__1157_ vdd gnd FILL
XFILL_2__1088_ vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_0__828_ vdd gnd FILL
X_1421_ _1694_/Q _1421_/B _1695_/Q _1422_/A _1423_/A vdd gnd OAI22X1
X_1352_ _1352_/A _1413_/B _1353_/C vdd gnd NAND2X1
XFILL_3__1404_ vdd gnd FILL
X_1283_ _1283_/A _1283_/B _1295_/A _1299_/A vdd gnd NAND3X1
XFILL_0__1626_ vdd gnd FILL
XFILL_3__1197_ vdd gnd FILL
XFILL_3__1335_ vdd gnd FILL
XFILL_3__1266_ vdd gnd FILL
XFILL_0__1557_ vdd gnd FILL
XFILL_0__1488_ vdd gnd FILL
XFILL_4__1513_ vdd gnd FILL
X_1619_ _1619_/A _1621_/B _1670_/B vdd gnd NOR2X1
XFILL_4__1375_ vdd gnd FILL
XFILL_4__1444_ vdd gnd FILL
XFILL_1__1597_ vdd gnd FILL
XFILL_1__1666_ vdd gnd FILL
XFILL_2__1011_ vdd gnd FILL
XFILL_2__988_ vdd gnd FILL
X_994_ _994_/A _994_/B _995_/B vdd gnd NAND2X1
XFILL_0__1411_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_3__1051_ vdd gnd FILL
XFILL_0__1273_ vdd gnd FILL
XFILL_3__1120_ vdd gnd FILL
XFILL_2__1209_ vdd gnd FILL
X_1404_ _1404_/A _1404_/B _1406_/C vdd gnd NOR2X1
X_1335_ _1556_/A _1549_/A _1338_/B vdd gnd NOR2X1
XFILL_3__1318_ vdd gnd FILL
X_1197_ _956_/Q _1197_/B _1197_/C _1197_/D _1305_/B vdd gnd OAI22X1
XFILL_4__1160_ vdd gnd FILL
XFILL_1__1382_ vdd gnd FILL
X_1266_ _1266_/A _1266_/B _1267_/A _1270_/A vdd gnd AOI21X1
XFILL_0__1609_ vdd gnd FILL
XFILL_1__1451_ vdd gnd FILL
XFILL_1__1520_ vdd gnd FILL
XFILL_2__911_ vdd gnd FILL
XFILL_3__1249_ vdd gnd FILL
XFILL_2__842_ vdd gnd FILL
XFILL_4__1091_ vdd gnd FILL
XFILL_1__1718_ vdd gnd FILL
XFILL_2__1560_ vdd gnd FILL
XFILL_2__1491_ vdd gnd FILL
XFILL_4__1427_ vdd gnd FILL
XFILL_4__1358_ vdd gnd FILL
XFILL_2_CLKBUF1_insert6 vdd gnd FILL
XFILL_1__1649_ vdd gnd FILL
XFILL_4__1289_ vdd gnd FILL
XCLKBUF1_insert5 clk _956_/CLK vdd gnd CLKBUF1
XFILL_1__860_ vdd gnd FILL
X_977_ _979_/B _979_/A _978_/B vdd gnd NAND2X1
X_1051_ _989_/B _1059_/C _1054_/B vdd gnd NOR2X1
X_1120_ _1689_/Q _1545_/A vdd gnd INVX1
XFILL_0__1325_ vdd gnd FILL
XFILL_3__1034_ vdd gnd FILL
XFILL_0__1256_ vdd gnd FILL
XFILL_3__1103_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
X_1318_ _1400_/B _1400_/A _979_/B _1347_/A vdd gnd OAI21X1
XFILL_1__989_ vdd gnd FILL
XFILL_4__1212_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
X_1249_ _1249_/A _1250_/C vdd gnd INVX1
XFILL_4__1074_ vdd gnd FILL
XFILL_4__1143_ vdd gnd FILL
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1503_ vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
X_831_ _936_/A _968_/A _898_/B _852_/A vdd gnd NAND3X1
X_900_ _934_/A _901_/A _935_/A _901_/C vdd gnd AOI21X1
XFILL_2__1612_ vdd gnd FILL
XFILL_2__1474_ vdd gnd FILL
XFILL_2__1543_ vdd gnd FILL
XFILL103950x50850 vdd gnd FILL
XFILL_0__1110_ vdd gnd FILL
XFILL103650x85950 vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_3__1721_ vdd gnd FILL
XFILL_1__912_ vdd gnd FILL
XFILL_1__843_ vdd gnd FILL
XFILL_3__1652_ vdd gnd FILL
XFILL_3__1583_ vdd gnd FILL
X_1034_ _975_/A _978_/A _1056_/B vdd gnd NAND2X1
X_1103_ _1683_/Q _1132_/B _1684_/Q _1133_/A vdd gnd OAI21X1
XFILL_1__1150_ vdd gnd FILL
XFILL_3__1017_ vdd gnd FILL
XFILL_4__985_ vdd gnd FILL
XFILL_0__1308_ vdd gnd FILL
XFILL_1__1081_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_2__1190_ vdd gnd FILL
XFILL_4__1057_ vdd gnd FILL
XFILL_1__1417_ vdd gnd FILL
XFILL_4__1126_ vdd gnd FILL
XFILL_0__861_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
XFILL103350x15750 vdd gnd FILL
XFILL_2__1526_ vdd gnd FILL
XFILL103950x62550 vdd gnd FILL
XFILL_0__1590_ vdd gnd FILL
XFILL_2__1457_ vdd gnd FILL
XFILL_2__1388_ vdd gnd FILL
X_1721_ _1721_/A rgb[6] vdd gnd BUFX2
XFILL_0__1024_ vdd gnd FILL
X_1652_ _1652_/A _1654_/A _1653_/A vdd gnd XOR2X1
X_1583_ _1583_/A _1677_/A _1583_/C _1585_/A vdd gnd OAI21X1
XFILL_3__1566_ vdd gnd FILL
XFILL_3__1635_ vdd gnd FILL
XFILL_3__1497_ vdd gnd FILL
XFILL_4__968_ vdd gnd FILL
XFILL_1__1202_ vdd gnd FILL
X_1017_ _1386_/D _1213_/B _1216_/B _1615_/C _1018_/A vdd gnd AOI22X1
XFILL_4__899_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_1__1133_ vdd gnd FILL
XFILL_4__1675_ vdd gnd FILL
XFILL_2__1242_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_0__913_ vdd gnd FILL
XFILL_2__1173_ vdd gnd FILL
XFILL_0__844_ vdd gnd FILL
XFILL_4__1109_ vdd gnd FILL
XFILL_3__1351_ vdd gnd FILL
XFILL103950x74250 vdd gnd FILL
XFILL_0__1711_ vdd gnd FILL
XFILL_3__986_ vdd gnd FILL
XFILL_3__1420_ vdd gnd FILL
XFILL_0__1642_ vdd gnd FILL
XFILL_0_BUFX2_insert0 vdd gnd FILL
XFILL_2__1509_ vdd gnd FILL
XFILL_0__1573_ vdd gnd FILL
XFILL_3__1282_ vdd gnd FILL
XFILL_0__1007_ vdd gnd FILL
X_1704_ _1704_/D vdd _1709_/S _1710_/CLK _971_/A vdd gnd DFFSR
X_1566_ _1693_/Q _1710_/Q _1577_/A vdd gnd NOR2X1
X_1635_ _1637_/C _1635_/B _1670_/B _1636_/C vdd gnd NAND3X1
X_1497_ _1688_/Q _1687_/Q _1680_/Q _1499_/C vdd gnd OAI21X1
XFILL_4__1460_ vdd gnd FILL
XFILL_3__1618_ vdd gnd FILL
XFILL_4__1391_ vdd gnd FILL
XFILL_3__1549_ vdd gnd FILL
XFILL_1__1116_ vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
XFILL_3__840_ vdd gnd FILL
XFILL_4__1589_ vdd gnd FILL
XFILL_4__1658_ vdd gnd FILL
XFILL_2__1225_ vdd gnd FILL
XFILL_2__1156_ vdd gnd FILL
XFILL103350x39150 vdd gnd FILL
XFILL_2__1087_ vdd gnd FILL
X_1351_ _1351_/A _1351_/B _1650_/A _1352_/A vdd gnd AOI21X1
X_1420_ _1420_/A _1420_/B _1423_/B vdd gnd AND2X2
XFILL_3__1334_ vdd gnd FILL
XFILL_3__1403_ vdd gnd FILL
XFILL_3__969_ vdd gnd FILL
X_1282_ _1291_/B _1291_/C _1283_/B vdd gnd AND2X2
XFILL_0__1625_ vdd gnd FILL
XFILL_3__1196_ vdd gnd FILL
XFILL_3__1265_ vdd gnd FILL
XFILL_0__1556_ vdd gnd FILL
XFILL_0__1487_ vdd gnd FILL
X_1618_ _1618_/A _1618_/B _1672_/B _1621_/B vdd gnd AOI21X1
XFILL_4__1512_ vdd gnd FILL
XFILL_4__1443_ vdd gnd FILL
X_1549_ _1549_/A _1675_/A _1555_/A vdd gnd NOR2X1
XFILL_1__1665_ vdd gnd FILL
XFILL_4__1374_ vdd gnd FILL
XFILL_1__1596_ vdd gnd FILL
XFILL_2__1010_ vdd gnd FILL
XFILL_2__987_ vdd gnd FILL
X_993_ _993_/A _999_/A _997_/A _994_/A vdd gnd OAI21X1
XFILL_0__1410_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
XFILL_2__1208_ vdd gnd FILL
XFILL_3__1050_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_2__1139_ vdd gnd FILL
X_1334_ _1359_/B _998_/A _1360_/A _1345_/B vdd gnd AOI21X1
X_1403_ _1599_/A _1403_/B _1404_/B vdd gnd NAND2X1
X_1265_ _1265_/A _1267_/A vdd gnd INVX1
X_1196_ _1513_/A _1401_/B _1196_/C _1197_/C vdd gnd OAI21X1
XFILL_2__910_ vdd gnd FILL
XFILL_3__1317_ vdd gnd FILL
XFILL_1__1381_ vdd gnd FILL
XFILL_0__1608_ vdd gnd FILL
XFILL_0__1539_ vdd gnd FILL
XFILL_4__1090_ vdd gnd FILL
XFILL_1__1450_ vdd gnd FILL
XFILL_3__1179_ vdd gnd FILL
XFILL_3__1248_ vdd gnd FILL
XFILL_2__841_ vdd gnd FILL
XFILL_4__1357_ vdd gnd FILL
XFILL_1__1648_ vdd gnd FILL
XFILL_1__1717_ vdd gnd FILL
XFILL_2__1490_ vdd gnd FILL
XFILL_4__1426_ vdd gnd FILL
XFILL_1__1579_ vdd gnd FILL
XFILL_4__1288_ vdd gnd FILL
XFILL_2_CLKBUF1_insert7 vdd gnd FILL
XCLKBUF1_insert6 clk _1710_/CLK vdd gnd CLKBUF1
X_976_ _979_/C _978_/A vdd gnd INVX2
X_1050_ _999_/Y _982_/A _1050_/C _1059_/C vdd gnd AOI21X1
XFILL_3__1102_ vdd gnd FILL
XFILL_0__1186_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
XFILL_3__1033_ vdd gnd FILL
XFILL_0__1255_ vdd gnd FILL
XFILL_4_BUFX2_insert11 vdd gnd FILL
X_1317_ _1317_/A _1317_/B _1696_/Q _1400_/B vdd gnd AOI21X1
XFILL_4__1211_ vdd gnd FILL
XFILL_1__988_ vdd gnd FILL
X_1248_ _1248_/A _1248_/B _1248_/C _1253_/A vdd gnd OAI21X1
XFILL_1__1502_ vdd gnd FILL
X_1179_ _1693_/Q _1317_/B _1332_/B _1327_/B vdd gnd NAND3X1
XFILL_1__1364_ vdd gnd FILL
XFILL_4__1073_ vdd gnd FILL
XFILL_4__1142_ vdd gnd FILL
XFILL_1__1433_ vdd gnd FILL
XFILL_1__1295_ vdd gnd FILL
X_830_ _953_/Q _952_/Q _898_/B vdd gnd NOR2X1
XFILL_2__1611_ vdd gnd FILL
XFILL_4__1409_ vdd gnd FILL
XFILL_2__1473_ vdd gnd FILL
XFILL_2__1542_ vdd gnd FILL
XFILL_0__1040_ vdd gnd FILL
XFILL_3__1720_ vdd gnd FILL
XFILL_1__911_ vdd gnd FILL
XFILL_1__842_ vdd gnd FILL
XFILL_3__1651_ vdd gnd FILL
X_959_ _959_/A _959_/B _965_/B vdd gnd NOR2X1
X_1102_ _1390_/A _1390_/B _1132_/B vdd gnd NAND2X1
XFILL_3__1582_ vdd gnd FILL
X_1033_ _1056_/C _1056_/A _1036_/C vdd gnd NOR2X1
XFILL_4__984_ vdd gnd FILL
XFILL_0__1169_ vdd gnd FILL
XFILL_3__1016_ vdd gnd FILL
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_4__1056_ vdd gnd FILL
XFILL_0__860_ vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
XFILL_4__1125_ vdd gnd FILL
XFILL_2__1525_ vdd gnd FILL
XFILL_2__1387_ vdd gnd FILL
XFILL_2__1456_ vdd gnd FILL
X_1720_ _1724_/A rgb[5] vdd gnd BUFX2
XFILL_0__989_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
X_1651_ _1671_/C _971_/A _1654_/A vdd gnd XOR2X1
XFILL_3__1634_ vdd gnd FILL
X_1582_ _1582_/A _1582_/B _1695_/Q _1586_/C vdd gnd OAI21X1
XFILL_3__1565_ vdd gnd FILL
XFILL_3__1496_ vdd gnd FILL
XFILL_4__898_ vdd gnd FILL
XFILL_1__1201_ vdd gnd FILL
X_1016_ _979_/A _1020_/A _1386_/D vdd gnd NOR2X1
XFILL_4__967_ vdd gnd FILL
XFILL_1__1132_ vdd gnd FILL
XFILL_1__1063_ vdd gnd FILL
XFILL_4__1674_ vdd gnd FILL
XFILL_2__1241_ vdd gnd FILL
XFILL_2__1310_ vdd gnd FILL
XFILL_0__912_ vdd gnd FILL
XFILL_4__1039_ vdd gnd FILL
XFILL_2__1172_ vdd gnd FILL
XFILL_0__843_ vdd gnd FILL
XFILL_4__1108_ vdd gnd FILL
XFILL_3__985_ vdd gnd FILL
XFILL_3__1350_ vdd gnd FILL
XFILL_0__1641_ vdd gnd FILL
XFILL_0__1572_ vdd gnd FILL
XFILL_3__1281_ vdd gnd FILL
XFILL_2__1508_ vdd gnd FILL
XFILL_0_BUFX2_insert1 vdd gnd FILL
XFILL_2__1439_ vdd gnd FILL
XFILL_0__1006_ vdd gnd FILL
X_1703_ _1703_/D vdd _1710_/R _1710_/CLK _971_/B vdd gnd DFFSR
X_1634_ _1634_/A _1645_/A _1635_/B vdd gnd OR2X2
XFILL_3__1617_ vdd gnd FILL
X_1565_ _1577_/B _1572_/A vdd gnd INVX1
X_1496_ _1507_/A _1496_/B _1543_/B _1524_/B vdd gnd OAI21X1
XFILL_4__1390_ vdd gnd FILL
XFILL_3__1479_ vdd gnd FILL
XFILL_3__1548_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_4__1588_ vdd gnd FILL
XFILL_4__1657_ vdd gnd FILL
XFILL_2__1224_ vdd gnd FILL
XFILL_2__1155_ vdd gnd FILL
XFILL_2__1086_ vdd gnd FILL
XFILL_3__968_ vdd gnd FILL
X_1350_ _1350_/A _1350_/B _1358_/B vdd gnd NAND2X1
X_1281_ _1686_/Q _1281_/B _1291_/C vdd gnd NAND2X1
XFILL_3__899_ vdd gnd FILL
XFILL_3__1333_ vdd gnd FILL
XFILL_3__1402_ vdd gnd FILL
XFILL_3__1264_ vdd gnd FILL
XFILL_0__1555_ vdd gnd FILL
XFILL_0__1624_ vdd gnd FILL
XFILL_3__1195_ vdd gnd FILL
XFILL_0__1486_ vdd gnd FILL
XFILL102750x85950 vdd gnd FILL
X_1617_ _981_/B _1617_/B _1618_/A vdd gnd NOR2X1
XFILL_4__1442_ vdd gnd FILL
XFILL_4__1373_ vdd gnd FILL
XFILL_4__1511_ vdd gnd FILL
XFILL_1__1664_ vdd gnd FILL
X_1479_ _1479_/A _1479_/B _1543_/B vdd gnd NAND2X1
X_1548_ _1708_/Q _1675_/A vdd gnd INVX1
XFILL_1__1595_ vdd gnd FILL
XFILL_2__986_ vdd gnd FILL
XFILL_1__1029_ vdd gnd FILL
XBUFX2_insert11 _1308_/Y _1702_/R vdd gnd BUFX2
X_992_ _992_/A _992_/B _994_/B vdd gnd NAND2X1
XFILL_2__1207_ vdd gnd FILL
XFILL_0__1340_ vdd gnd FILL
XFILL_0__1271_ vdd gnd FILL
XFILL_2__1138_ vdd gnd FILL
X_1402_ _1604_/A _1605_/B _1404_/A vdd gnd NAND2X1
XFILL_2__1069_ vdd gnd FILL
X_1333_ _992_/A _1333_/B _1360_/A vdd gnd NOR2X1
X_1264_ _1268_/B _1268_/A _1264_/C _1270_/D vdd gnd NAND3X1
XFILL102450x15750 vdd gnd FILL
XFILL_3__1316_ vdd gnd FILL
X_1195_ _975_/A _1400_/C _1196_/C vdd gnd NAND2X1
XFILL_3__1247_ vdd gnd FILL
XFILL_1__1380_ vdd gnd FILL
XFILL_0__1607_ vdd gnd FILL
XFILL_0__1469_ vdd gnd FILL
XFILL_0__1538_ vdd gnd FILL
XFILL_3__1178_ vdd gnd FILL
XFILL_2__840_ vdd gnd FILL
XFILL_4__1356_ vdd gnd FILL
XFILL_1__1716_ vdd gnd FILL
XFILL_4__1425_ vdd gnd FILL
XFILL_1__1647_ vdd gnd FILL
XFILL_1__1578_ vdd gnd FILL
XFILL_2__969_ vdd gnd FILL
XFILL_2_CLKBUF1_insert8 vdd gnd FILL
XFILL_4__1287_ vdd gnd FILL
XCLKBUF1_insert7 clk _945_/CLK vdd gnd CLKBUF1
X_975_ _975_/A _981_/A vdd gnd INVX1
XFILL_0__1323_ vdd gnd FILL
XFILL_3__1101_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
XFILL_3__1032_ vdd gnd FILL
XFILL_0__1254_ vdd gnd FILL
XFILL_4_BUFX2_insert12 vdd gnd FILL
X_1178_ _1324_/A _1324_/B _1184_/B vdd gnd NOR2X1
X_1316_ _1599_/A _1327_/B _1400_/A vdd gnd NOR2X1
XFILL_4__1210_ vdd gnd FILL
XFILL_1__987_ vdd gnd FILL
X_1247_ _1556_/A _986_/A _1247_/C _1248_/C vdd gnd OAI21X1
XFILL_1__1501_ vdd gnd FILL
XFILL_1__1432_ vdd gnd FILL
XFILL_1__1363_ vdd gnd FILL
XFILL_4__1141_ vdd gnd FILL
XFILL_4__1072_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
XFILL_2__1610_ vdd gnd FILL
XFILL_2__1541_ vdd gnd FILL
XFILL_4__1339_ vdd gnd FILL
XFILL_2__1472_ vdd gnd FILL
XFILL_4__1408_ vdd gnd FILL
XFILL_1__910_ vdd gnd FILL
XFILL_3__1650_ vdd gnd FILL
X_1032_ _968_/A _1663_/A _1056_/A vdd gnd NOR2X1
X_889_ _889_/A _944_/D vdd gnd INVX1
XFILL_1__841_ vdd gnd FILL
X_958_ _958_/A _959_/B vdd gnd INVX1
XFILL_3__1581_ vdd gnd FILL
X_1101_ _1682_/Q _1390_/B vdd gnd INVX1
XFILL_3__1015_ vdd gnd FILL
XFILL_0__1306_ vdd gnd FILL
XFILL102450x39150 vdd gnd FILL
XFILL_4__983_ vdd gnd FILL
XFILL_0__1237_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
XFILL_0__1099_ vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_4__1124_ vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_4__1055_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
XFILL_2__1524_ vdd gnd FILL
XFILL_2__1386_ vdd gnd FILL
XFILL_2__1455_ vdd gnd FILL
XFILL_0__988_ vdd gnd FILL
XFILL_0__1022_ vdd gnd FILL
X_1650_ _1650_/A _1671_/C _1650_/C _1652_/A vdd gnd OAI21X1
X_1581_ _1583_/A _1595_/B _1581_/C _1694_/D vdd gnd OAI21X1
XFILL_3__1633_ vdd gnd FILL
X_1015_ _971_/A _1015_/B _1020_/A vdd gnd NOR2X1
XFILL_3__1564_ vdd gnd FILL
XFILL_3__1495_ vdd gnd FILL
XFILL_4__897_ vdd gnd FILL
XFILL_1__1200_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
XFILL_4__966_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
XFILL_4__1673_ vdd gnd FILL
XFILL_2__1171_ vdd gnd FILL
XFILL_2__1240_ vdd gnd FILL
XFILL_4__1107_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_0__911_ vdd gnd FILL
XFILL_4__1038_ vdd gnd FILL
XFILL_0__842_ vdd gnd FILL
XFILL_3__984_ vdd gnd FILL
XFILL_0_BUFX2_insert2 vdd gnd FILL
XFILL_2__1438_ vdd gnd FILL
XFILL_0__1571_ vdd gnd FILL
XFILL_3__1280_ vdd gnd FILL
XFILL_2__1507_ vdd gnd FILL
XFILL_0__1640_ vdd gnd FILL
XFILL_2__1369_ vdd gnd FILL
XFILL_0__1005_ vdd gnd FILL
X_1564_ _1564_/A _1564_/B _1564_/C _1577_/B vdd gnd AOI21X1
X_1633_ _1645_/A _1634_/A _1637_/C vdd gnd NAND2X1
X_1702_ _1702_/D vdd _1702_/R _1702_/CLK _998_/A vdd gnd DFFSR
XFILL_3__1616_ vdd gnd FILL
XFILL_3__1547_ vdd gnd FILL
X_1495_ _1495_/A _1541_/A _1539_/A _1496_/B vdd gnd NAND3X1
XFILL_3__1478_ vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_4__1725_ vdd gnd FILL
XFILL_4__1656_ vdd gnd FILL
XFILL_4__1587_ vdd gnd FILL
XFILL_2__1223_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
XFILL_2__1085_ vdd gnd FILL
XFILL_3__898_ vdd gnd FILL
XFILL_3__1401_ vdd gnd FILL
XFILL_3__967_ vdd gnd FILL
X_1280_ _1537_/A _962_/B _1291_/B vdd gnd OR2X2
XFILL_3__1194_ vdd gnd FILL
XFILL_3__1332_ vdd gnd FILL
XFILL_3__1263_ vdd gnd FILL
XFILL_0__1623_ vdd gnd FILL
XFILL_0__1485_ vdd gnd FILL
XFILL_0__1554_ vdd gnd FILL
X_1616_ down _1616_/B _1616_/C _1617_/B vdd gnd NAND3X1
X_1547_ _1547_/A _1549_/A _1690_/D vdd gnd XOR2X1
XFILL_4__1441_ vdd gnd FILL
XFILL_4__1372_ vdd gnd FILL
XFILL_1__1594_ vdd gnd FILL
XFILL_1__1663_ vdd gnd FILL
X_1478_ _1478_/A _1498_/B _1478_/C _1479_/A vdd gnd NAND3X1
XFILL_2__985_ vdd gnd FILL
XFILL_1__1028_ vdd gnd FILL
XBUFX2_insert12 _1308_/Y _1709_/S vdd gnd BUFX2
XFILL_4__1639_ vdd gnd FILL
X_991_ _997_/A _992_/A vdd gnd INVX2
XFILL_2__1206_ vdd gnd FILL
XFILL_0__1270_ vdd gnd FILL
XFILL_2__1068_ vdd gnd FILL
XFILL_2__1137_ vdd gnd FILL
X_1401_ _1401_/A _1401_/B _1677_/C vdd gnd NOR2X1
X_1194_ _1197_/B _1401_/B vdd gnd INVX1
XFILL_0__1606_ vdd gnd FILL
X_1332_ _1332_/A _1332_/B _1333_/B vdd gnd NAND2X1
X_1263_ _1297_/B _1297_/A _1268_/A vdd gnd XOR2X1
XFILL_3__1177_ vdd gnd FILL
XFILL_3__1315_ vdd gnd FILL
XFILL_3__1246_ vdd gnd FILL
XFILL_0__1468_ vdd gnd FILL
XFILL_0__1537_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL_1__1715_ vdd gnd FILL
XFILL_4__1355_ vdd gnd FILL
XFILL_4__1424_ vdd gnd FILL
XFILL_1__1577_ vdd gnd FILL
XFILL_1__1646_ vdd gnd FILL
XFILL_4__1286_ vdd gnd FILL
XFILL_2__968_ vdd gnd FILL
XFILL_2_CLKBUF1_insert9 vdd gnd FILL
XFILL_2__899_ vdd gnd FILL
XCLKBUF1_insert8 clk _949_/CLK vdd gnd CLKBUF1
X_974_ _974_/A _974_/B _974_/Y vdd gnd NAND2X1
XFILL_0__1322_ vdd gnd FILL
XFILL_3__1031_ vdd gnd FILL
XFILL_3__1100_ vdd gnd FILL
XFILL_0__1184_ vdd gnd FILL
XFILL_0__1253_ vdd gnd FILL
XFILL_4_BUFX2_insert13 vdd gnd FILL
X_1315_ _1663_/A _1315_/B _1315_/C _1347_/B vdd gnd NAND3X1
XFILL_1__986_ vdd gnd FILL
X_1177_ _1177_/A _1177_/B _1177_/C _1185_/B vdd gnd NAND3X1
X_1246_ _1254_/A _1254_/B _1249_/A _1266_/B vdd gnd OAI21X1
XFILL_1__1362_ vdd gnd FILL
XFILL_4__1140_ vdd gnd FILL
XFILL_1__1500_ vdd gnd FILL
XFILL_1__1431_ vdd gnd FILL
XFILL_3__1229_ vdd gnd FILL
XFILL_4__1071_ vdd gnd FILL
XFILL_1__1293_ vdd gnd FILL
XFILL_4__1407_ vdd gnd FILL
XFILL_2__1471_ vdd gnd FILL
XFILL_2__1540_ vdd gnd FILL
XFILL_4__1338_ vdd gnd FILL
XFILL_4__1269_ vdd gnd FILL
XFILL_1__1629_ vdd gnd FILL
XFILL_1__840_ vdd gnd FILL
X_957_ _957_/A _959_/A vdd gnd INVX1
XFILL_3__1580_ vdd gnd FILL
X_1031_ _979_/B _1663_/A vdd gnd INVX1
X_888_ _935_/A _891_/B _888_/C _889_/A vdd gnd NAND3X1
X_1100_ _1681_/Q _1390_/A vdd gnd INVX1
XFILL_2__1669_ vdd gnd FILL
XFILL_4__982_ vdd gnd FILL
XFILL_0__1236_ vdd gnd FILL
XFILL_3__1014_ vdd gnd FILL
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
XFILL_0__1098_ vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_0_BUFX2_insert11 vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
X_1229_ _1229_/A _1229_/B _1229_/C _1230_/C vdd gnd OAI21X1
XFILL_1__1345_ vdd gnd FILL
XFILL_4__1054_ vdd gnd FILL
XFILL_4__1123_ vdd gnd FILL
XFILL_1__1276_ vdd gnd FILL
XFILL_2__1454_ vdd gnd FILL
XFILL_2__1523_ vdd gnd FILL
XFILL_2__1385_ vdd gnd FILL
XFILL_0__987_ vdd gnd FILL
XFILL_0__1021_ vdd gnd FILL
X_1580_ _1595_/B _1583_/C _1580_/C _1581_/C vdd gnd NAND3X1
XFILL_3__1632_ vdd gnd FILL
XFILL_3__1563_ vdd gnd FILL
X_1014_ _1421_/B _1615_/C vdd gnd INVX1
XFILL_3__1494_ vdd gnd FILL
XFILL_0__1219_ vdd gnd FILL
XFILL_4__896_ vdd gnd FILL
XFILL_1__1061_ vdd gnd FILL
XFILL_4__965_ vdd gnd FILL
XFILL_1__1130_ vdd gnd FILL
XFILL_4__1672_ vdd gnd FILL
XFILL_4__1037_ vdd gnd FILL
XFILL_1__1328_ vdd gnd FILL
XFILL_0__910_ vdd gnd FILL
XFILL_2__1170_ vdd gnd FILL
XFILL_4__1106_ vdd gnd FILL
XFILL_0__841_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL_3__983_ vdd gnd FILL
XFILL_0_BUFX2_insert3 vdd gnd FILL
XFILL_2__1437_ vdd gnd FILL
XFILL_0__1570_ vdd gnd FILL
XFILL_2__1506_ vdd gnd FILL
XFILL_2__1368_ vdd gnd FILL
X_1701_ _1701_/D vdd _1702_/R _1702_/CLK _997_/A vdd gnd DFFSR
XFILL_2__1299_ vdd gnd FILL
XFILL_0__1004_ vdd gnd FILL
X_1632_ _1671_/C _992_/A _1645_/A vdd gnd XOR2X1
X_1494_ _1536_/C _1536_/B _1494_/C _1495_/A vdd gnd AOI21X1
X_1563_ _1563_/A _1619_/A _1563_/C _1692_/D vdd gnd OAI21X1
XFILL_3__1615_ vdd gnd FILL
XFILL_3__1477_ vdd gnd FILL
XFILL_3__1546_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_4__879_ vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL_4__1724_ vdd gnd FILL
XFILL_4__1655_ vdd gnd FILL
XFILL_4__1586_ vdd gnd FILL
XFILL_2__1222_ vdd gnd FILL
XFILL_2__1153_ vdd gnd FILL
XFILL_2__1084_ vdd gnd FILL
XFILL_3__1400_ vdd gnd FILL
XFILL_3__897_ vdd gnd FILL
XFILL_3__1331_ vdd gnd FILL
XFILL_3__966_ vdd gnd FILL
XFILL_0__1622_ vdd gnd FILL
XFILL_3__1193_ vdd gnd FILL
XFILL_3__1262_ vdd gnd FILL
XFILL_0__1484_ vdd gnd FILL
XFILL_0__1553_ vdd gnd FILL
XFILL_4__1440_ vdd gnd FILL
X_1615_ _971_/A _1615_/B _1615_/C _1616_/C vdd gnd NAND3X1
X_1477_ _1477_/A _1498_/B vdd gnd INVX1
X_1546_ _1708_/Q _1546_/B _1547_/A vdd gnd NAND2X1
XFILL_4__1371_ vdd gnd FILL
XFILL_1__1593_ vdd gnd FILL
XFILL_3__1529_ vdd gnd FILL
XFILL_1__1662_ vdd gnd FILL
XFILL_2__984_ vdd gnd FILL
XBUFX2_insert13 _1308_/Y _1710_/R vdd gnd BUFX2
X_990_ _990_/A _997_/B vdd gnd INVX2
XFILL_1__1027_ vdd gnd FILL
XFILL_4__1569_ vdd gnd FILL
XFILL_4__1638_ vdd gnd FILL
XFILL_2__1205_ vdd gnd FILL
XFILL103350x11850 vdd gnd FILL
XFILL103050x46950 vdd gnd FILL
XFILL_2__1067_ vdd gnd FILL
XFILL_2__1136_ vdd gnd FILL
XFILL103650x93750 vdd gnd FILL
X_1400_ _1400_/A _1400_/B _1400_/C _1401_/A vdd gnd OAI21X1
X_1331_ _1361_/A _1345_/A vdd gnd INVX1
X_1193_ _1193_/A _1193_/B _1193_/C _1197_/D vdd gnd AOI21X1
XFILL_0__1605_ vdd gnd FILL
X_1262_ _1262_/A _1262_/B _1268_/B vdd gnd XOR2X1
XFILL_3__1314_ vdd gnd FILL
XFILL_3__1176_ vdd gnd FILL
XFILL_3__1245_ vdd gnd FILL
XFILL_0__1398_ vdd gnd FILL
XFILL_0__1467_ vdd gnd FILL
XFILL_0__1536_ vdd gnd FILL
XFILL_1__1714_ vdd gnd FILL
XFILL_4__1423_ vdd gnd FILL
X_1529_ _960_/A _958_/A _1530_/C vdd gnd NOR2X1
XFILL_1__1645_ vdd gnd FILL
XFILL_4__1354_ vdd gnd FILL
XFILL_1__1576_ vdd gnd FILL
XFILL_4__1285_ vdd gnd FILL
XFILL_2__898_ vdd gnd FILL
XFILL_2__967_ vdd gnd FILL
X_973_ _979_/A _979_/B _974_/B vdd gnd XOR2X1
XCLKBUF1_insert9 clk _1709_/CLK vdd gnd CLKBUF1
XFILL_0__1321_ vdd gnd FILL
XFILL_3__1030_ vdd gnd FILL
XFILL103950x70350 vdd gnd FILL
XFILL_0__1252_ vdd gnd FILL
XFILL_4_BUFX2_insert14 vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
XFILL_2__1119_ vdd gnd FILL
XFILL_1__985_ vdd gnd FILL
X_1314_ _1314_/A _1314_/B _1314_/C _1410_/B vdd gnd AOI21X1
X_1176_ _951_/Q _1359_/B _1176_/C _1177_/C vdd gnd OAI21X1
XFILL_1__1361_ vdd gnd FILL
X_1245_ _1252_/A _1245_/B _1249_/A vdd gnd XOR2X1
XFILL_1__1430_ vdd gnd FILL
XFILL_4__1070_ vdd gnd FILL
XFILL_0__1519_ vdd gnd FILL
XFILL_3__1228_ vdd gnd FILL
XFILL_3__1159_ vdd gnd FILL
XFILL_1__1292_ vdd gnd FILL
XFILL_4__1406_ vdd gnd FILL
XFILL_2__1470_ vdd gnd FILL
XFILL_1__1628_ vdd gnd FILL
XFILL_4__1337_ vdd gnd FILL
XFILL_4__1199_ vdd gnd FILL
XFILL_4__1268_ vdd gnd FILL
XFILL_1__1559_ vdd gnd FILL
XFILL103350x35250 vdd gnd FILL
X_956_ _956_/D vdd _956_/R _956_/CLK _956_/Q vdd gnd DFFSR
X_1030_ _975_/A _978_/A _1056_/C vdd gnd NOR2X1
XFILL_4__981_ vdd gnd FILL
X_887_ _890_/B _890_/C _891_/B vdd gnd NAND2X1
XFILL_2__1599_ vdd gnd FILL
XFILL_2__1668_ vdd gnd FILL
XFILL_0__1166_ vdd gnd FILL
XFILL_3__1013_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
XFILL_0__1304_ vdd gnd FILL
XFILL_0__1097_ vdd gnd FILL
X_1228_ _1228_/A _1228_/B _1229_/C vdd gnd NOR2X1
XFILL_1__968_ vdd gnd FILL
XFILL_1__899_ vdd gnd FILL
XFILL_0_BUFX2_insert12 vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
X_1159_ _1573_/A _1406_/A _1330_/B vdd gnd NAND2X1
XFILL_1__1344_ vdd gnd FILL
XFILL_4__1053_ vdd gnd FILL
XFILL_1__1275_ vdd gnd FILL
XFILL_4__1122_ vdd gnd FILL
XFILL_2__1384_ vdd gnd FILL
XFILL_2__1453_ vdd gnd FILL
XFILL_2__1522_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
XFILL_0__1020_ vdd gnd FILL
X_939_ _939_/D vdd _956_/R _949_/CLK _960_/A vdd gnd DFFSR
XFILL_3__1631_ vdd gnd FILL
XFILL_3__1493_ vdd gnd FILL
XFILL_3__1562_ vdd gnd FILL
X_1013_ _952_/Q _1216_/B vdd gnd INVX1
XFILL_4__964_ vdd gnd FILL
XFILL_0__1218_ vdd gnd FILL
XFILL_0__1149_ vdd gnd FILL
XFILL_4__895_ vdd gnd FILL
XFILL_1__1060_ vdd gnd FILL
XFILL_4__1671_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_4__1036_ vdd gnd FILL
XFILL_0__840_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_4__1105_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
XFILL_3__982_ vdd gnd FILL
XFILL_2__1367_ vdd gnd FILL
XFILL_2__1436_ vdd gnd FILL
XFILL_2__1505_ vdd gnd FILL
XFILL_0__969_ vdd gnd FILL
XFILL_0__1003_ vdd gnd FILL
X_1631_ _1646_/A _1634_/A vdd gnd INVX1
X_1700_ _1700_/D vdd _1709_/S _1702_/CLK _993_/A vdd gnd DFFSR
XFILL_2__1298_ vdd gnd FILL
XFILL_3__1614_ vdd gnd FILL
X_1493_ _1493_/A _1518_/A _1521_/A _1494_/C vdd gnd NAND3X1
X_1562_ _1582_/A _1582_/B _1692_/Q _1563_/C vdd gnd OAI21X1
XFILL_3__1476_ vdd gnd FILL
XFILL_3__1545_ vdd gnd FILL
XFILL_4__878_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
XFILL_1__1043_ vdd gnd FILL
XFILL_4__1723_ vdd gnd FILL
XFILL_4__1585_ vdd gnd FILL
XFILL_2__1221_ vdd gnd FILL
XFILL_2__1152_ vdd gnd FILL
XFILL_4__1019_ vdd gnd FILL
XFILL_2__1083_ vdd gnd FILL
XFILL_3__965_ vdd gnd FILL
XFILL_3__1330_ vdd gnd FILL
XFILL_3__896_ vdd gnd FILL
XFILL_0__1552_ vdd gnd FILL
XFILL_0__1621_ vdd gnd FILL
XFILL_3__1192_ vdd gnd FILL
XFILL_2__1419_ vdd gnd FILL
XFILL_3__1261_ vdd gnd FILL
XFILL_0__1483_ vdd gnd FILL
X_1614_ _998_/A _994_/B _1614_/C _1615_/B vdd gnd OAI21X1
XFILL_4__1370_ vdd gnd FILL
XFILL_1__1661_ vdd gnd FILL
X_1476_ _1687_/Q _1680_/Q _1478_/A vdd gnd NAND2X1
X_1545_ _1545_/A _1595_/B _1689_/D vdd gnd NOR2X1
XFILL_3__1528_ vdd gnd FILL
XFILL_1__1592_ vdd gnd FILL
XFILL_3__1459_ vdd gnd FILL
XFILL_2__983_ vdd gnd FILL
XBUFX2_insert14 _1308_/Y _1689_/R vdd gnd BUFX2
XFILL_1__1026_ vdd gnd FILL
XFILL_4__1568_ vdd gnd FILL
XFILL_4__1637_ vdd gnd FILL
XFILL_4__1499_ vdd gnd FILL
XFILL_3_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__1204_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
XFILL_2__1066_ vdd gnd FILL
X_1330_ _998_/Y _1330_/B _1330_/C _1361_/A vdd gnd NAND3X1
X_1261_ _1287_/A _1262_/B vdd gnd INVX1
X_1192_ _975_/A _1400_/C _968_/A _1355_/B _1193_/C vdd gnd OAI22X1
XFILL_3__1244_ vdd gnd FILL
XFILL_0__1604_ vdd gnd FILL
XFILL_0__1535_ vdd gnd FILL
XFILL_3__879_ vdd gnd FILL
XFILL_3__1313_ vdd gnd FILL
XFILL_3__1175_ vdd gnd FILL
XFILL_0__1397_ vdd gnd FILL
XFILL_0__1466_ vdd gnd FILL
XFILL_4__1353_ vdd gnd FILL
X_1528_ _1528_/A _1528_/B _1528_/C _1535_/A vdd gnd NAND3X1
XFILL_4__1422_ vdd gnd FILL
XFILL_1__1713_ vdd gnd FILL
X_1459_ _1683_/Q _1680_/Q _1492_/B vdd gnd XOR2X1
XFILL_1__1644_ vdd gnd FILL
XFILL_1__1575_ vdd gnd FILL
XFILL_4__1284_ vdd gnd FILL
XFILL_2__897_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
XFILL_2__966_ vdd gnd FILL
X_972_ _992_/B _972_/B _972_/C _979_/A vdd gnd AOI21X1
XFILL103950x89850 vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_0__1320_ vdd gnd FILL
XFILL_0__1251_ vdd gnd FILL
XFILL_4_BUFX2_insert15 vdd gnd FILL
XFILL_2__1118_ vdd gnd FILL
XFILL_2__1049_ vdd gnd FILL
XFILL_1__984_ vdd gnd FILL
X_1244_ _1253_/B _1254_/B vdd gnd INVX1
X_1313_ _1544_/A _1542_/A _1313_/C _1314_/C vdd gnd NAND3X1
X_1175_ _1175_/A _1175_/B _1175_/C _1176_/C vdd gnd AOI21X1
XFILL_3__1227_ vdd gnd FILL
XFILL_1__1360_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
XFILL_0__1518_ vdd gnd FILL
XFILL_3__1158_ vdd gnd FILL
XFILL_3__1089_ vdd gnd FILL
XFILL_0__1449_ vdd gnd FILL
XFILL_4__1405_ vdd gnd FILL
XFILL_4__1336_ vdd gnd FILL
XFILL_1__1558_ vdd gnd FILL
XFILL_1__1627_ vdd gnd FILL
XFILL_4__1198_ vdd gnd FILL
XFILL_4__1267_ vdd gnd FILL
XFILL_1__1489_ vdd gnd FILL
XFILL103650x19650 vdd gnd FILL
X_955_ _955_/D vdd _956_/R _956_/CLK _975_/A vdd gnd DFFSR
X_886_ _886_/A _886_/B _890_/B vdd gnd NOR2X1
XFILL_2__1667_ vdd gnd FILL
XFILL_4__980_ vdd gnd FILL
XFILL_2__1598_ vdd gnd FILL
XFILL_0__1303_ vdd gnd FILL
XFILL_3__1012_ vdd gnd FILL
XFILL_0__1165_ vdd gnd FILL
XFILL_0__1234_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
XFILL_1__1412_ vdd gnd FILL
X_1227_ _1227_/A _1227_/B _1228_/B vdd gnd NOR2X1
XFILL_1__898_ vdd gnd FILL
X_1158_ _1691_/Q _1692_/Q _1690_/Q _1406_/A vdd gnd NOR3X1
XFILL_1__967_ vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_1__1343_ vdd gnd FILL
XFILL_4__1052_ vdd gnd FILL
X_1089_ _1687_/Q _1096_/A _1107_/A _1121_/B vdd gnd NAND3X1
XFILL_1__1274_ vdd gnd FILL
XFILL_4__1121_ vdd gnd FILL
XFILL_2__1521_ vdd gnd FILL
XFILL_2__1383_ vdd gnd FILL
XFILL_2__1452_ vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
XFILL_3__1630_ vdd gnd FILL
X_1012_ _953_/Q _1213_/B vdd gnd INVX1
X_938_ _938_/D vdd _956_/R _956_/CLK _938_/Q vdd gnd DFFSR
X_869_ _885_/C _869_/B _870_/A vdd gnd NAND2X1
XFILL_3__1561_ vdd gnd FILL
XFILL_2__1719_ vdd gnd FILL
XFILL_3__1492_ vdd gnd FILL
XFILL102450x11850 vdd gnd FILL
XFILL_4__894_ vdd gnd FILL
XFILL_4__963_ vdd gnd FILL
XFILL_0__1217_ vdd gnd FILL
XFILL_0__1148_ vdd gnd FILL
XFILL_0__1079_ vdd gnd FILL
XFILL_4__1670_ vdd gnd FILL
XFILL_4__1104_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
XFILL_4__1035_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_3__981_ vdd gnd FILL
XFILL_2__1504_ vdd gnd FILL
XFILL_2__1366_ vdd gnd FILL
XFILL_2__1297_ vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_0__968_ vdd gnd FILL
XFILL_0__899_ vdd gnd FILL
XFILL_0__1002_ vdd gnd FILL
X_1630_ _1630_/A _999_/A _1630_/C _1646_/A vdd gnd AOI21X1
XFILL_3__1613_ vdd gnd FILL
X_1561_ _1564_/A _1564_/B _1563_/A vdd gnd XNOR2X1
X_1492_ _1492_/A _1492_/B _1518_/A vdd gnd XNOR2X1
XFILL_3__1475_ vdd gnd FILL
XFILL_3__1544_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL_4__877_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
XFILL_4__1722_ vdd gnd FILL
XFILL_4__1653_ vdd gnd FILL
XFILL_4__1584_ vdd gnd FILL
XFILL_2__1220_ vdd gnd FILL
XFILL_2__1151_ vdd gnd FILL
XFILL_4__1018_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_3__895_ vdd gnd FILL
XFILL_3__964_ vdd gnd FILL
XFILL_0__1551_ vdd gnd FILL
XFILL_0__1482_ vdd gnd FILL
XFILL_0__1620_ vdd gnd FILL
XFILL_2__1418_ vdd gnd FILL
XFILL_3__1260_ vdd gnd FILL
XFILL_3__1191_ vdd gnd FILL
XFILL_2__1349_ vdd gnd FILL
X_1613_ _998_/A _997_/A _1613_/C _1614_/C vdd gnd NAND3X1
X_1544_ _1544_/A _1595_/B _1544_/C _1544_/D _1688_/D vdd gnd OAI22X1
XFILL_3__1527_ vdd gnd FILL
XFILL_1__1591_ vdd gnd FILL
XFILL_1__1660_ vdd gnd FILL
X_1475_ _1477_/A _1475_/B _1479_/B vdd gnd NAND2X1
XFILL_2__982_ vdd gnd FILL
XFILL_3__1389_ vdd gnd FILL
XFILL_3__1458_ vdd gnd FILL
XFILL_4__929_ vdd gnd FILL
XFILL_1__1025_ vdd gnd FILL
XBUFX2_insert15 _1308_/Y _1708_/R vdd gnd BUFX2
XFILL_4__1636_ vdd gnd FILL
XFILL_3_CLKBUF1_insert5 vdd gnd FILL
XFILL_4__1567_ vdd gnd FILL
XFILL_4__1498_ vdd gnd FILL
XFILL_2__1203_ vdd gnd FILL
XFILL_2__1134_ vdd gnd FILL
XFILL_2__1065_ vdd gnd FILL
X_1191_ _1348_/B _1348_/C _1400_/C vdd gnd NAND2X1
XFILL_3__878_ vdd gnd FILL
X_1260_ _1260_/A _1289_/A _1287_/A vdd gnd NAND2X1
XFILL_3__1174_ vdd gnd FILL
XFILL_3__1243_ vdd gnd FILL
XFILL_0__1603_ vdd gnd FILL
XFILL_0__1534_ vdd gnd FILL
XFILL_0__1465_ vdd gnd FILL
XFILL_3__1312_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ _990_/A _953_/Q _1528_/B vdd gnd NOR2X1
XFILL_4__1352_ vdd gnd FILL
XFILL_1__1712_ vdd gnd FILL
XFILL_4__1421_ vdd gnd FILL
X_1389_ _1389_/A _1389_/B _1389_/C _1398_/A vdd gnd OAI21X1
XFILL_1__1643_ vdd gnd FILL
XFILL_1__1574_ vdd gnd FILL
XFILL_4__1283_ vdd gnd FILL
X_1458_ _1482_/B _1480_/A _1481_/A _1492_/A vdd gnd OAI21X1
XFILL_2__965_ vdd gnd FILL
XFILL_2__896_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
X_971_ _971_/A _971_/B _972_/C vdd gnd NAND2X1
XFILL_4__1619_ vdd gnd FILL
XFILL_0__1181_ vdd gnd FILL
XFILL_2__1048_ vdd gnd FILL
XFILL_0__1250_ vdd gnd FILL
XFILL_2__1117_ vdd gnd FILL
X_1174_ _990_/A _1342_/B _1175_/B vdd gnd NAND2X1
X_1243_ _1243_/A _1247_/C _1243_/C _1253_/B vdd gnd NAND3X1
XFILL_1__983_ vdd gnd FILL
X_1312_ _1686_/Q _1685_/Q _1313_/C vdd gnd NOR2X1
XFILL_3__1226_ vdd gnd FILL
XFILL_3__1157_ vdd gnd FILL
XFILL_0__1517_ vdd gnd FILL
XFILL_1__1290_ vdd gnd FILL
XFILL_0__1448_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_3__1088_ vdd gnd FILL
XFILL_4__1404_ vdd gnd FILL
XFILL_4__1335_ vdd gnd FILL
XFILL_4__1266_ vdd gnd FILL
XFILL_1__1557_ vdd gnd FILL
XFILL_1__1626_ vdd gnd FILL
XFILL_4__1197_ vdd gnd FILL
XFILL_1__1488_ vdd gnd FILL
XFILL_2__879_ vdd gnd FILL
X_954_ _954_/D _954_/S vdd _956_/CLK _968_/A vdd gnd DFFSR
X_885_ _885_/A _885_/B _885_/C _890_/C vdd gnd NOR3X1
XFILL_2__1597_ vdd gnd FILL
XFILL_2__1666_ vdd gnd FILL
XFILL_3__1011_ vdd gnd FILL
XFILL_0__1302_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
XFILL_0__1233_ vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
XFILL_2_CLKBUF1_insert10 vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_1__1411_ vdd gnd FILL
X_1226_ _1226_/A _1226_/B _1226_/C _1229_/B vdd gnd AOI21X1
XFILL_1__897_ vdd gnd FILL
XFILL_1__1342_ vdd gnd FILL
X_1157_ _1692_/Q _1173_/A _1693_/Q _1330_/C vdd gnd OAI21X1
XFILL_0_BUFX2_insert14 vdd gnd FILL
XFILL_4__1120_ vdd gnd FILL
XFILL_3__1209_ vdd gnd FILL
XFILL_4__1051_ vdd gnd FILL
XFILL_1__1273_ vdd gnd FILL
X_1088_ _1540_/A _1537_/A _1096_/A vdd gnd NOR2X1
XFILL_2__1451_ vdd gnd FILL
XFILL_2__1520_ vdd gnd FILL
XFILL_4__1318_ vdd gnd FILL
XFILL_4__1249_ vdd gnd FILL
XFILL_2__1382_ vdd gnd FILL
XFILL_1__1609_ vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_3__1560_ vdd gnd FILL
XFILL_2__1718_ vdd gnd FILL
X_937_ _937_/A _937_/B _956_/D vdd gnd NOR2X1
X_1011_ _1011_/A _996_/Y _1011_/C _1018_/B vdd gnd OAI21X1
X_868_ _957_/A _960_/A _938_/Q _885_/C vdd gnd NAND3X1
XFILL_2__1649_ vdd gnd FILL
XFILL_3__1491_ vdd gnd FILL
XFILL_0__1216_ vdd gnd FILL
XFILL_4__893_ vdd gnd FILL
XFILL_4__962_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
XFILL_0__1078_ vdd gnd FILL
XFILL_1__1325_ vdd gnd FILL
X_1209_ _1209_/A _1210_/A vdd gnd INVX1
XFILL_4__1034_ vdd gnd FILL
XFILL_4__1103_ vdd gnd FILL
XFILL_1__1187_ vdd gnd FILL
XFILL_1__1256_ vdd gnd FILL
XFILL_3__980_ vdd gnd FILL
XFILL_2__1434_ vdd gnd FILL
XFILL_2__1503_ vdd gnd FILL
XFILL_2__1365_ vdd gnd FILL
XFILL_2__1296_ vdd gnd FILL
XFILL_0__898_ vdd gnd FILL
XFILL_0__1001_ vdd gnd FILL
XFILL_0__967_ vdd gnd FILL
X_1560_ _1560_/A _1564_/C _1564_/B vdd gnd NOR2X1
XFILL_3__1612_ vdd gnd FILL
XFILL_3__1543_ vdd gnd FILL
X_1491_ _1504_/A _1493_/A vdd gnd INVX1
XFILL_3__1474_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
XFILL_4__876_ vdd gnd FILL
XFILL_1__1110_ vdd gnd FILL
XFILL_4__1652_ vdd gnd FILL
XFILL_4__1721_ vdd gnd FILL
X_1689_ _1689_/D vdd _1689_/R _1689_/CLK _1689_/Q vdd gnd DFFSR
XFILL_4__1583_ vdd gnd FILL
XFILL_2__1150_ vdd gnd FILL
XFILL_4__1017_ vdd gnd FILL
XFILL_1__1308_ vdd gnd FILL
XFILL_2__1081_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_3__894_ vdd gnd FILL
XFILL_3__963_ vdd gnd FILL
XFILL_3__1190_ vdd gnd FILL
XFILL_2__1417_ vdd gnd FILL
XFILL_0__1481_ vdd gnd FILL
XFILL_0__1550_ vdd gnd FILL
XFILL_2__1348_ vdd gnd FILL
XFILL_2__1279_ vdd gnd FILL
X_1612_ _1612_/A _1613_/C vdd gnd INVX1
X_1474_ _1688_/Q _1680_/Q _1477_/A vdd gnd XNOR2X1
X_1543_ _1602_/C _1543_/B _1544_/C vdd gnd NAND2X1
XFILL102750x19650 vdd gnd FILL
XFILL_3__1526_ vdd gnd FILL
XFILL_1__1590_ vdd gnd FILL
XFILL_4__928_ vdd gnd FILL
XFILL_2__981_ vdd gnd FILL
XFILL_3__1388_ vdd gnd FILL
XFILL_3__1457_ vdd gnd FILL
XFILL_4__859_ vdd gnd FILL
XFILL_1__1024_ vdd gnd FILL
XFILL_4__1566_ vdd gnd FILL
XFILL_4__1635_ vdd gnd FILL
XFILL_3_CLKBUF1_insert6 vdd gnd FILL
XFILL_4__1497_ vdd gnd FILL
XFILL_2__1202_ vdd gnd FILL
XFILL_2__1064_ vdd gnd FILL
XFILL_2__1133_ vdd gnd FILL
X_1190_ _1599_/A _1327_/B _1604_/A _1348_/C vdd gnd OAI21X1
XFILL_3__877_ vdd gnd FILL
XFILL_0__1602_ vdd gnd FILL
XFILL_3__1311_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
XFILL_3__1173_ vdd gnd FILL
XFILL_3__1242_ vdd gnd FILL
XFILL_0__1533_ vdd gnd FILL
XFILL_0__1464_ vdd gnd FILL
X_1526_ _951_/Q _985_/B _1528_/C vdd gnd NOR2X1
XFILL_1__1711_ vdd gnd FILL
XFILL_4__1420_ vdd gnd FILL
X_1457_ _1682_/Q _1679_/Q _1480_/A vdd gnd NOR2X1
XFILL_4__1351_ vdd gnd FILL
X_1388_ _1697_/Q _1388_/B _1618_/B _1698_/Q _1389_/C vdd gnd AOI22X1
XFILL_3__1509_ vdd gnd FILL
XFILL_1__1642_ vdd gnd FILL
XFILL_1__1573_ vdd gnd FILL
XFILL_4__1282_ vdd gnd FILL
XFILL_2__895_ vdd gnd FILL
XFILL_2__964_ vdd gnd FILL
X_970_ _998_/A _997_/A _972_/B vdd gnd NOR2X1
XFILL_1__1007_ vdd gnd FILL
XFILL_4__1618_ vdd gnd FILL
XFILL_4__1549_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
XFILL_2__1047_ vdd gnd FILL
XFILL_2__1116_ vdd gnd FILL
XFILL_1__982_ vdd gnd FILL
X_1311_ _1390_/A _1390_/B _1314_/B _1314_/A vdd gnd OAI21X1
XFILL_3__929_ vdd gnd FILL
X_1173_ _1173_/A _1243_/A _1247_/C _1175_/A vdd gnd NAND3X1
X_1242_ _1247_/C _1243_/A _1243_/C _1254_/A vdd gnd AOI21X1
XFILL_3__1225_ vdd gnd FILL
XFILL_3__1156_ vdd gnd FILL
XFILL_0__1378_ vdd gnd FILL
XFILL_0__1516_ vdd gnd FILL
XFILL_0__1447_ vdd gnd FILL
XFILL_3__1087_ vdd gnd FILL
XFILL_4__1403_ vdd gnd FILL
X_1509_ _968_/A _965_/C _1509_/C _1511_/A vdd gnd NAND3X1
XFILL_4__1196_ vdd gnd FILL
XFILL_4__1334_ vdd gnd FILL
XFILL_4__1265_ vdd gnd FILL
XFILL_1__1556_ vdd gnd FILL
XFILL_1__1487_ vdd gnd FILL
XFILL_1__1625_ vdd gnd FILL
XFILL_2__878_ vdd gnd FILL
X_953_ _953_/D vdd _954_/S _956_/CLK _953_/Q vdd gnd DFFSR
XFILL_2__1596_ vdd gnd FILL
X_884_ _886_/B _884_/B _886_/A _888_/C vdd gnd OAI21X1
XFILL_2__1665_ vdd gnd FILL
XFILL_0__1232_ vdd gnd FILL
XFILL_3__1010_ vdd gnd FILL
XFILL_0__1301_ vdd gnd FILL
XFILL_0__1163_ vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
XFILL_1__965_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
X_1225_ _1225_/A _1229_/A _1235_/C vdd gnd NOR2X1
XFILL_1__1341_ vdd gnd FILL
X_1156_ _1556_/A _1549_/A _1173_/A vdd gnd NAND2X1
XFILL_1__896_ vdd gnd FILL
XFILL_4__1050_ vdd gnd FILL
X_1087_ _1685_/Q _1537_/A vdd gnd INVX2
XFILL_1__1410_ vdd gnd FILL
XFILL_3__1208_ vdd gnd FILL
XFILL_1__1272_ vdd gnd FILL
XFILL_3__1139_ vdd gnd FILL
XFILL_1__1608_ vdd gnd FILL
XFILL_2__1450_ vdd gnd FILL
XFILL_4__1317_ vdd gnd FILL
XFILL_4__1179_ vdd gnd FILL
XFILL_4__1248_ vdd gnd FILL
XFILL_2__1381_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
XFILL_1__1539_ vdd gnd FILL
X_936_ _936_/A _937_/B _955_/D vdd gnd NOR2X1
XFILL_2__1717_ vdd gnd FILL
XFILL_3__1490_ vdd gnd FILL
X_867_ _867_/A _938_/D _867_/C _869_/B vdd gnd OAI21X1
X_1010_ _951_/Q _1383_/B _1421_/B _952_/Q _1011_/C vdd gnd AOI22X1
XFILL_2__1648_ vdd gnd FILL
XFILL_4__961_ vdd gnd FILL
XFILL_2__1579_ vdd gnd FILL
XFILL102450x7950 vdd gnd FILL
XFILL_0__1215_ vdd gnd FILL
XFILL_4__892_ vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
XFILL_0__1077_ vdd gnd FILL
X_1208_ _1252_/B _1208_/B _1232_/A _1211_/A vdd gnd OAI21X1
XFILL_1__879_ vdd gnd FILL
XFILL_1__1324_ vdd gnd FILL
XFILL_4__1033_ vdd gnd FILL
XFILL_1__1255_ vdd gnd FILL
XFILL_4__1102_ vdd gnd FILL
X_1139_ _1139_/A _1139_/B _1305_/A vdd gnd NAND2X1
XFILL_1__1186_ vdd gnd FILL
XFILL_2__1364_ vdd gnd FILL
XFILL_2__1433_ vdd gnd FILL
XFILL_2__1502_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_2__1295_ vdd gnd FILL
XFILL_0__897_ vdd gnd FILL
X_1490_ _1490_/A _1490_/B _1521_/A vdd gnd XNOR2X1
X_919_ _951_/Q _952_/Q _919_/C _933_/B vdd gnd NAND3X1
XFILL_3__1473_ vdd gnd FILL
XFILL_3__1542_ vdd gnd FILL
XFILL_3__1611_ vdd gnd FILL
XFILL_1__1040_ vdd gnd FILL
XFILL_4__875_ vdd gnd FILL
XFILL_0__1129_ vdd gnd FILL
XFILL_4__1720_ vdd gnd FILL
XFILL_4__1651_ vdd gnd FILL
X_1688_ _1688_/D vdd _1689_/R _1689_/CLK _1688_/Q vdd gnd DFFSR
XFILL_4__1582_ vdd gnd FILL
XFILL_4__1016_ vdd gnd FILL
XFILL_2__1080_ vdd gnd FILL
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_3__893_ vdd gnd FILL
XFILL_3__962_ vdd gnd FILL
XFILL103350x31350 vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
XFILL_2__1347_ vdd gnd FILL
XFILL_0__1480_ vdd gnd FILL
XFILL103050x66450 vdd gnd FILL
XFILL_2__1278_ vdd gnd FILL
X_1611_ _1671_/C _1672_/B vdd gnd INVX1
X_1473_ _1542_/A _1473_/B _1478_/C _1475_/B vdd gnd OAI21X1
X_1542_ _1542_/A _1595_/B _1542_/C _1544_/D _1687_/D vdd gnd OAI22X1
XFILL_3__1525_ vdd gnd FILL
XFILL_3__1456_ vdd gnd FILL
XFILL_4__927_ vdd gnd FILL
XFILL_3__1387_ vdd gnd FILL
XFILL_2__980_ vdd gnd FILL
XFILL_4__858_ vdd gnd FILL
XFILL_1__1023_ vdd gnd FILL
XFILL_4__1565_ vdd gnd FILL
XFILL_4__1634_ vdd gnd FILL
XFILL_2__1201_ vdd gnd FILL
XFILL_3_CLKBUF1_insert7 vdd gnd FILL
XFILL_4__1496_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_2__1132_ vdd gnd FILL
XFILL103350x43050 vdd gnd FILL
XFILL_3__876_ vdd gnd FILL
XFILL_0__1601_ vdd gnd FILL
XFILL_0__1532_ vdd gnd FILL
XFILL_3__1310_ vdd gnd FILL
XFILL_3__1172_ vdd gnd FILL
XFILL_3__1241_ vdd gnd FILL
XFILL_0__1463_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
XFILL_4__1350_ vdd gnd FILL
X_1525_ _956_/Q _986_/A _1528_/A vdd gnd NOR2X1
X_1387_ _1387_/A _1387_/B _1387_/C _1389_/B vdd gnd AOI21X1
XFILL_1__1641_ vdd gnd FILL
X_1456_ _1681_/Q _1678_/Q _1482_/B vdd gnd NAND2X1
XFILL_3__1439_ vdd gnd FILL
XFILL_1__1572_ vdd gnd FILL
XFILL_4__1281_ vdd gnd FILL
XFILL_3__1508_ vdd gnd FILL
XFILL_2__894_ vdd gnd FILL
XFILL_2__963_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_4__1617_ vdd gnd FILL
XFILL_4__1479_ vdd gnd FILL
XFILL_4__1548_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
XFILL_2__1046_ vdd gnd FILL
XFILL_3__928_ vdd gnd FILL
X_1241_ _1248_/A _1248_/B _1243_/C vdd gnd NOR2X1
XFILL_1__981_ vdd gnd FILL
X_1310_ _1523_/A _1520_/A _1314_/B vdd gnd NOR2X1
XFILL_3__859_ vdd gnd FILL
XFILL_3__1224_ vdd gnd FILL
X_1172_ _1691_/Q _987_/B _1245_/B _1247_/C vdd gnd OAI21X1
XFILL_0__1515_ vdd gnd FILL
XFILL_0__1377_ vdd gnd FILL
XFILL_0__1446_ vdd gnd FILL
XFILL_3__1155_ vdd gnd FILL
XFILL_3__1086_ vdd gnd FILL
XFILL_4__1333_ vdd gnd FILL
XFILL_4__1402_ vdd gnd FILL
X_1439_ _1512_/B _997_/B _1441_/B vdd gnd NAND2X1
X_1508_ _1619_/A _1508_/B _1508_/C _1682_/D vdd gnd OAI21X1
XFILL_1__1624_ vdd gnd FILL
XFILL_4__1195_ vdd gnd FILL
XFILL_4__1264_ vdd gnd FILL
XFILL_1__1555_ vdd gnd FILL
XFILL_1__1486_ vdd gnd FILL
XFILL_2__877_ vdd gnd FILL
X_952_ _952_/D vdd _954_/S _956_/CLK _952_/Q vdd gnd DFFSR
X_883_ _962_/A _886_/A vdd gnd INVX1
XFILL_2__1595_ vdd gnd FILL
XFILL_2__1664_ vdd gnd FILL
XFILL_0__1162_ vdd gnd FILL
XFILL_0__1231_ vdd gnd FILL
XFILL_0__1300_ vdd gnd FILL
XFILL_2__1029_ vdd gnd FILL
XFILL_0__1093_ vdd gnd FILL
X_1224_ _1227_/A _1224_/B _1224_/C _1229_/A vdd gnd NAND3X1
XFILL_1__895_ vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
XFILL_3__1207_ vdd gnd FILL
XFILL_1__1340_ vdd gnd FILL
X_1155_ _1690_/Q _1549_/A vdd gnd INVX2
XFILL_1__1271_ vdd gnd FILL
X_1086_ _1686_/Q _1540_/A vdd gnd INVX1
XFILL_0__1429_ vdd gnd FILL
XFILL_3__1069_ vdd gnd FILL
XFILL_3__1138_ vdd gnd FILL
XFILL_4__1316_ vdd gnd FILL
XFILL_2__1380_ vdd gnd FILL
XFILL_1__1607_ vdd gnd FILL
XFILL_1__1538_ vdd gnd FILL
XFILL_4__1178_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
XFILL_4__1247_ vdd gnd FILL
XFILL_1__1469_ vdd gnd FILL
XFILL_2__929_ vdd gnd FILL
X_935_ _935_/A _935_/B _935_/C _954_/D vdd gnd OAI21X1
X_866_ _957_/A _867_/C vdd gnd INVX1
XFILL_2__1716_ vdd gnd FILL
XFILL_2__1647_ vdd gnd FILL
XFILL_4__891_ vdd gnd FILL
XFILL_4__960_ vdd gnd FILL
XFILL_2__1578_ vdd gnd FILL
XFILL_0__1214_ vdd gnd FILL
XFILL_0__1145_ vdd gnd FILL
XFILL_0__1076_ vdd gnd FILL
X_1207_ _982_/A _1549_/A _1252_/B vdd gnd NAND2X1
XFILL_1__878_ vdd gnd FILL
XFILL_1__1323_ vdd gnd FILL
XFILL_4__1032_ vdd gnd FILL
XFILL_1__1254_ vdd gnd FILL
X_1069_ _1069_/A _1069_/B _1070_/C vdd gnd NOR2X1
XFILL_4__1101_ vdd gnd FILL
X_1138_ _965_/C _1428_/A _1138_/C _1138_/D _1139_/A vdd gnd AOI22X1
XFILL_1__1185_ vdd gnd FILL
XFILL103050x7950 vdd gnd FILL
XFILL_2__1501_ vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_2__1294_ vdd gnd FILL
XFILL_2__1432_ vdd gnd FILL
XFILL_0__896_ vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
XFILL103950x85950 vdd gnd FILL
XFILL_3__1610_ vdd gnd FILL
X_918_ _938_/D _931_/B _952_/Q _923_/C vdd gnd OAI21X1
X_849_ _864_/B _854_/B _849_/C _850_/C vdd gnd OAI21X1
XFILL_3__1472_ vdd gnd FILL
XFILL_3__1541_ vdd gnd FILL
XFILL_4__874_ vdd gnd FILL
XFILL_0__1059_ vdd gnd FILL
XFILL_0__1128_ vdd gnd FILL
XFILL_4__1650_ vdd gnd FILL
XFILL_4__1581_ vdd gnd FILL
X_1687_ _1687_/D vdd _1689_/R _1689_/CLK _1687_/Q vdd gnd DFFSR
XFILL_1__1237_ vdd gnd FILL
XFILL_1__1168_ vdd gnd FILL
XFILL_4__1015_ vdd gnd FILL
XFILL_1__1306_ vdd gnd FILL
XFILL_3__961_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_3__892_ vdd gnd FILL
XFILL103650x15750 vdd gnd FILL
XFILL_2__1346_ vdd gnd FILL
XFILL_2__1415_ vdd gnd FILL
XFILL_2__1277_ vdd gnd FILL
XFILL_0__879_ vdd gnd FILL
X_1610_ _1623_/A _1623_/B up _1671_/C vdd gnd OAI21X1
X_1472_ _1498_/A _1483_/A _1478_/C vdd gnd NAND2X1
X_1541_ _1541_/A _1621_/A _1542_/C vdd gnd OR2X2
XFILL_3__1386_ vdd gnd FILL
XFILL_0__1677_ vdd gnd FILL
XFILL_3__1524_ vdd gnd FILL
XFILL_3__1455_ vdd gnd FILL
XFILL_4__926_ vdd gnd FILL
XFILL_4__857_ vdd gnd FILL
XFILL_1__1022_ vdd gnd FILL
XFILL_3_CLKBUF1_insert8 vdd gnd FILL
XFILL_4__1564_ vdd gnd FILL
XFILL_4__1633_ vdd gnd FILL
XFILL_4__1495_ vdd gnd FILL
XFILL_2__1200_ vdd gnd FILL
XFILL_2__1131_ vdd gnd FILL
XFILL_2__1062_ vdd gnd FILL
XFILL103650x27450 vdd gnd FILL
XFILL_0__1531_ vdd gnd FILL
XFILL_3__875_ vdd gnd FILL
XFILL_0__1600_ vdd gnd FILL
XFILL_3__1240_ vdd gnd FILL
XFILL_0__1462_ vdd gnd FILL
XFILL_2__1329_ vdd gnd FILL
XFILL_3__1171_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
X_1524_ _1524_/A _1524_/B _1544_/D vdd gnd NAND2X1
X_1386_ _1599_/A _974_/B _1403_/B _1386_/D _1387_/C vdd gnd OAI22X1
XFILL_1__1571_ vdd gnd FILL
XFILL_3__1507_ vdd gnd FILL
X_1455_ _1682_/Q _1679_/Q _1481_/A vdd gnd NAND2X1
XFILL_1__1640_ vdd gnd FILL
XFILL_3__1438_ vdd gnd FILL
XFILL_3__1369_ vdd gnd FILL
XFILL_2__962_ vdd gnd FILL
XFILL_4__1280_ vdd gnd FILL
XFILL_4__909_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_2__893_ vdd gnd FILL
XFILL_4__1616_ vdd gnd FILL
XFILL_4__1547_ vdd gnd FILL
XFILL_4__1478_ vdd gnd FILL
XFILL_2__1114_ vdd gnd FILL
XFILL_2__1045_ vdd gnd FILL
XFILL103650x39150 vdd gnd FILL
XFILL_3__927_ vdd gnd FILL
XFILL_3__858_ vdd gnd FILL
X_1171_ _982_/A _1549_/A _1245_/B vdd gnd NOR2X1
XFILL_1__980_ vdd gnd FILL
X_1240_ _1297_/A _1288_/A _1265_/A vdd gnd NOR2X1
XFILL_3__1223_ vdd gnd FILL
XFILL_3__1154_ vdd gnd FILL
XFILL_0__1514_ vdd gnd FILL
XFILL_0__1445_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
XFILL_3__1085_ vdd gnd FILL
X_1507_ _1507_/A _1524_/A _1524_/B _1508_/B vdd gnd NAND3X1
XFILL_4__1401_ vdd gnd FILL
XFILL_4__1332_ vdd gnd FILL
X_1438_ _1438_/A _1510_/C _1442_/C vdd gnd AND2X2
X_1369_ _1430_/B _1430_/A _1399_/C vdd gnd NAND2X1
XFILL_4__1263_ vdd gnd FILL
XFILL_1__1623_ vdd gnd FILL
XFILL_1__1554_ vdd gnd FILL
XFILL_4__1194_ vdd gnd FILL
XFILL_1__1485_ vdd gnd FILL
XFILL_2__876_ vdd gnd FILL
X_951_ _951_/D vdd _954_/S _956_/CLK _951_/Q vdd gnd DFFSR
X_882_ _886_/B _884_/B _882_/C _943_/D vdd gnd AOI21X1
XFILL_2__1663_ vdd gnd FILL
XFILL_2__1594_ vdd gnd FILL
XFILL_0__1161_ vdd gnd FILL
XFILL_0__1230_ vdd gnd FILL
XFILL_2__1028_ vdd gnd FILL
XFILL_0__1092_ vdd gnd FILL
X_1223_ _1228_/A _1227_/B _1224_/C vdd gnd NOR2X1
X_1154_ _1691_/Q _1556_/A vdd gnd INVX2
XFILL_1__894_ vdd gnd FILL
XFILL_1__963_ vdd gnd FILL
XFILL_3__1206_ vdd gnd FILL
XFILL_1__1270_ vdd gnd FILL
XFILL_0__1428_ vdd gnd FILL
X_1085_ _1124_/C _1520_/A _1523_/A _1107_/A vdd gnd AOI21X1
XFILL_3__1137_ vdd gnd FILL
XFILL_0__1359_ vdd gnd FILL
XFILL_3__1068_ vdd gnd FILL
XFILL_4__1315_ vdd gnd FILL
XFILL_1__1606_ vdd gnd FILL
XFILL_4__1246_ vdd gnd FILL
XFILL_1__1537_ vdd gnd FILL
XFILL_4__1177_ vdd gnd FILL
XFILL_2__928_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
XFILL_1__1468_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_2__859_ vdd gnd FILL
X_934_ _934_/A _934_/B _934_/C _935_/B vdd gnd NAND3X1
X_865_ _935_/A _937_/B vdd gnd INVX1
XFILL_2__1715_ vdd gnd FILL
XFILL_2__1646_ vdd gnd FILL
XFILL_4__890_ vdd gnd FILL
XFILL_2__1577_ vdd gnd FILL
XFILL_0__1213_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
XFILL_0__1075_ vdd gnd FILL
XFILL102450x43050 vdd gnd FILL
X_1206_ _1243_/A _1208_/B vdd gnd INVX1
XFILL_1__877_ vdd gnd FILL
X_1137_ _1137_/A _1137_/B _1138_/D vdd gnd NOR2X1
XFILL_4__1100_ vdd gnd FILL
XFILL_1__1184_ vdd gnd FILL
XFILL_1__1322_ vdd gnd FILL
XFILL_1__1253_ vdd gnd FILL
X_1068_ _1674_/C _956_/Q _1068_/C _1069_/B vdd gnd OAI21X1
XFILL_2__1500_ vdd gnd FILL
XFILL_2__1431_ vdd gnd FILL
XFILL_4__1229_ vdd gnd FILL
XFILL_2__1362_ vdd gnd FILL
XFILL_2__1293_ vdd gnd FILL
XFILL_0__895_ vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_3__1540_ vdd gnd FILL
X_917_ _935_/A _917_/B _917_/C _951_/D vdd gnd OAI21X1
X_848_ _848_/A _848_/B _894_/A _854_/B vdd gnd AOI21X1
XFILL_3__1471_ vdd gnd FILL
XFILL_2__1629_ vdd gnd FILL
XFILL_4__873_ vdd gnd FILL
XFILL_0__1058_ vdd gnd FILL
XFILL_0__1127_ vdd gnd FILL
X_1686_ _1686_/D vdd _1689_/R _1689_/CLK _1686_/Q vdd gnd DFFSR
XFILL_1__929_ vdd gnd FILL
XFILL_4__1580_ vdd gnd FILL
XFILL_3__1669_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_4__1014_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_3__891_ vdd gnd FILL
XFILL_3__960_ vdd gnd FILL
XFILL_2__1414_ vdd gnd FILL
XFILL_2__1345_ vdd gnd FILL
XFILL_2__1276_ vdd gnd FILL
XFILL_0__878_ vdd gnd FILL
X_1540_ _1540_/A _1595_/B _1540_/C _1544_/D _1686_/D vdd gnd OAI22X1
X_1471_ _1687_/Q _1680_/Q _1498_/A vdd gnd XOR2X1
XFILL_3__1523_ vdd gnd FILL
XFILL_3__1385_ vdd gnd FILL
XFILL_0__1676_ vdd gnd FILL
XFILL_3__1454_ vdd gnd FILL
XFILL_4__925_ vdd gnd FILL
XFILL_4__856_ vdd gnd FILL
XFILL_1__1021_ vdd gnd FILL
XFILL_4__1632_ vdd gnd FILL
X_1669_ _1670_/B _1669_/B _1669_/C _1670_/C vdd gnd NAND3X1
XFILL_4__1494_ vdd gnd FILL
XFILL_3_CLKBUF1_insert9 vdd gnd FILL
XFILL_4__1563_ vdd gnd FILL
XFILL_2__1061_ vdd gnd FILL
XFILL_2__1130_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL_3__874_ vdd gnd FILL
XFILL_3__1170_ vdd gnd FILL
XFILL_0__1530_ vdd gnd FILL
XFILL_0__1461_ vdd gnd FILL
XFILL_2__1328_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2_BUFX2_insert0 vdd gnd FILL
X_1454_ _1489_/A _1462_/B vdd gnd INVX1
X_1523_ _1523_/A _1546_/B _1523_/C _1684_/D vdd gnd OAI21X1
X_1385_ _1386_/D _1403_/B _1583_/A _1615_/C _1387_/A vdd gnd AOI22X1
XFILL_1__1570_ vdd gnd FILL
XFILL_3__1506_ vdd gnd FILL
XFILL_4__908_ vdd gnd FILL
XFILL_3__1437_ vdd gnd FILL
XFILL_3__1368_ vdd gnd FILL
XFILL_2__961_ vdd gnd FILL
XFILL_0__1659_ vdd gnd FILL
XFILL_3__1299_ vdd gnd FILL
XFILL_4__839_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_2__892_ vdd gnd FILL
XFILL_4__1615_ vdd gnd FILL
XFILL_4__1546_ vdd gnd FILL
XFILL_4__1477_ vdd gnd FILL
XFILL_2__1044_ vdd gnd FILL
XFILL_2__1113_ vdd gnd FILL
XFILL_3__926_ vdd gnd FILL
XFILL_3__857_ vdd gnd FILL
X_1170_ _1691_/Q _987_/B _1243_/A vdd gnd NAND2X1
XFILL_3__1153_ vdd gnd FILL
XFILL_0__1375_ vdd gnd FILL
XFILL_3__1222_ vdd gnd FILL
XFILL_0__1513_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
XFILL_3__1084_ vdd gnd FILL
XFILL_4__1400_ vdd gnd FILL
X_1437_ _975_/A _974_/A _1438_/A vdd gnd NOR2X1
X_1506_ _1582_/A _1582_/B _1682_/Q _1508_/C vdd gnd OAI21X1
XFILL_4__1331_ vdd gnd FILL
X_1368_ _1417_/A _1430_/A vdd gnd INVX1
XFILL_4__1262_ vdd gnd FILL
XFILL_1__1622_ vdd gnd FILL
XFILL_1__1484_ vdd gnd FILL
X_1299_ _1299_/A _1299_/B _1300_/B vdd gnd NOR2X1
XFILL_1__1553_ vdd gnd FILL
XFILL_4__1193_ vdd gnd FILL
XFILL_2__875_ vdd gnd FILL
X_950_ _950_/D vdd _954_/S _956_/CLK _990_/A vdd gnd DFFSR
X_881_ _886_/B _884_/B _935_/A _882_/C vdd gnd OAI21X1
XFILL_2__1593_ vdd gnd FILL
XFILL_4__1529_ vdd gnd FILL
XFILL_2__1662_ vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_2__1027_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
XFILL_3__909_ vdd gnd FILL
X_1153_ _1395_/B _1395_/A _1197_/B vdd gnd NAND2X1
X_1222_ _1697_/Q _981_/A _1227_/B vdd gnd NOR2X1
XFILL_1__893_ vdd gnd FILL
X_1084_ _1681_/Q _1682_/Q _1124_/C vdd gnd NOR2X1
XFILL102750x15750 vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_3__1205_ vdd gnd FILL
XFILL_3__1067_ vdd gnd FILL
XFILL_3__1136_ vdd gnd FILL
XFILL_0__1427_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL_4__1176_ vdd gnd FILL
XFILL_4__1245_ vdd gnd FILL
XFILL_1__1605_ vdd gnd FILL
XFILL_1__1467_ vdd gnd FILL
XFILL_1__1536_ vdd gnd FILL
XFILL_4__1314_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_2__858_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
XFILL_2__1714_ vdd gnd FILL
X_933_ _933_/A _933_/B _933_/C _934_/C vdd gnd OAI21X1
X_864_ _964_/A _864_/B _938_/Q _935_/A vdd gnd OAI21X1
XFILL_2__1576_ vdd gnd FILL
XFILL_2__1645_ vdd gnd FILL
XFILL_0__1212_ vdd gnd FILL
XFILL_0__1074_ vdd gnd FILL
XFILL_0__1143_ vdd gnd FILL
XFILL_1__1321_ vdd gnd FILL
XFILL_4__1030_ vdd gnd FILL
X_1205_ _986_/A _1556_/A _1232_/A vdd gnd NAND2X1
XFILL_1__876_ vdd gnd FILL
X_1067_ _1530_/A _1281_/B _1068_/C vdd gnd NOR2X1
X_1136_ _1136_/A _1136_/B _1136_/C _1137_/A vdd gnd NAND3X1
XFILL_1__1183_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_3__1119_ vdd gnd FILL
XFILL_2__1430_ vdd gnd FILL
XFILL_4__1228_ vdd gnd FILL
XFILL_4__1159_ vdd gnd FILL
XFILL_2__1361_ vdd gnd FILL
XFILL_2__1292_ vdd gnd FILL
XFILL_1__1519_ vdd gnd FILL
XFILL_0__894_ vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
X_916_ _928_/B _916_/B _934_/A _917_/B vdd gnd NAND3X1
XFILL_3__1470_ vdd gnd FILL
X_847_ _958_/A _965_/A _848_/B vdd gnd NOR2X1
XFILL_2__1559_ vdd gnd FILL
XFILL_2__1628_ vdd gnd FILL
XFILL_4__872_ vdd gnd FILL
XFILL102750x39150 vdd gnd FILL
XFILL_0__1057_ vdd gnd FILL
XFILL_3_BUFX2_insert11 vdd gnd FILL
X_1685_ _1685_/D vdd _1689_/R _1689_/CLK _1685_/Q vdd gnd DFFSR
XFILL_0__1126_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__859_ vdd gnd FILL
XFILL_3__1599_ vdd gnd FILL
XFILL_3__1668_ vdd gnd FILL
XFILL_4__1013_ vdd gnd FILL
XFILL_1__1235_ vdd gnd FILL
XFILL_1__1304_ vdd gnd FILL
X_1119_ _1544_/A _1121_/B _1689_/Q _1123_/A vdd gnd OAI21X1
XFILL_1__1166_ vdd gnd FILL
XFILL_1__1097_ vdd gnd FILL
XFILL_3__890_ vdd gnd FILL
XFILL_2__1413_ vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL_2__1275_ vdd gnd FILL
XFILL_0__877_ vdd gnd FILL
X_1470_ _1500_/B _1488_/B _1499_/A _1483_/A vdd gnd OAI21X1
XFILL_3__1453_ vdd gnd FILL
XFILL_3__1522_ vdd gnd FILL
XFILL_4__924_ vdd gnd FILL
XFILL_3__1384_ vdd gnd FILL
XFILL_0__1675_ vdd gnd FILL
XFILL_4__855_ vdd gnd FILL
XFILL_1__1020_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
X_1599_ _1599_/A _1599_/B _1677_/A _1600_/B vdd gnd OAI21X1
XFILL_4__1631_ vdd gnd FILL
X_1668_ _1668_/A _1668_/B _1669_/B vdd gnd NAND2X1
XFILL_4__1562_ vdd gnd FILL
XFILL_4__1493_ vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_2__1060_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_3__873_ vdd gnd FILL
XFILL_2__1327_ vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_0__1460_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
XFILL_2__1189_ vdd gnd FILL
XFILL_2__1258_ vdd gnd FILL
XFILL_2_BUFX2_insert1 vdd gnd FILL
X_1453_ _1684_/Q _1680_/Q _1489_/A vdd gnd NOR2X1
X_1522_ _1524_/A _1522_/B _1524_/B _1523_/C vdd gnd NAND3X1
XFILL_3__1436_ vdd gnd FILL
X_1384_ _1420_/B _1420_/A _1387_/B vdd gnd NAND2X1
XFILL_3__1505_ vdd gnd FILL
XFILL_0__1658_ vdd gnd FILL
XFILL_4__907_ vdd gnd FILL
XFILL_3__1367_ vdd gnd FILL
XFILL_2__891_ vdd gnd FILL
XFILL_0__1589_ vdd gnd FILL
XFILL_2__960_ vdd gnd FILL
XFILL_3__1298_ vdd gnd FILL
XFILL_4__838_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_4__1614_ vdd gnd FILL
XFILL_4__1545_ vdd gnd FILL
XFILL_4__1476_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL103650x7950 vdd gnd FILL
XFILL_2__1112_ vdd gnd FILL
XFILL_3__925_ vdd gnd FILL
XFILL_3__856_ vdd gnd FILL
XFILL_0__1512_ vdd gnd FILL
XFILL_3__1221_ vdd gnd FILL
XFILL_3__1152_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
XFILL_3__1083_ vdd gnd FILL
X_1367_ _1367_/A _1367_/B _1367_/C _1417_/A vdd gnd OAI21X1
XFILL_4__1330_ vdd gnd FILL
X_1436_ _953_/Q _952_/Q _1510_/C vdd gnd NOR2X1
XFILL_1__1621_ vdd gnd FILL
X_1505_ _1619_/A _1505_/B _1505_/C _1681_/D vdd gnd OAI21X1
XFILL_4__1192_ vdd gnd FILL
XFILL_3__1419_ vdd gnd FILL
XFILL_4__1261_ vdd gnd FILL
XFILL_1__1552_ vdd gnd FILL
XFILL_1__1483_ vdd gnd FILL
X_1298_ _1681_/Q _1298_/B _1298_/C _1299_/B vdd gnd OAI21X1
XFILL_2__874_ vdd gnd FILL
XFILL_4__1528_ vdd gnd FILL
X_880_ _965_/A _880_/B _884_/B vdd gnd NAND2X1
XFILL_2__1592_ vdd gnd FILL
XFILL_2__1661_ vdd gnd FILL
XFILL_4__1459_ vdd gnd FILL
XFILL_2__1026_ vdd gnd FILL
XFILL_0__1090_ vdd gnd FILL
X_1221_ _975_/A _1604_/A _1228_/A vdd gnd NOR2X1
XFILL_3__908_ vdd gnd FILL
XFILL103050x62550 vdd gnd FILL
XFILL_1__892_ vdd gnd FILL
XFILL_1__961_ vdd gnd FILL
X_1152_ _1348_/B _1605_/B _1395_/A vdd gnd OR2X2
XFILL_3__1204_ vdd gnd FILL
XFILL_3__839_ vdd gnd FILL
X_1083_ _1683_/Q _1520_/A vdd gnd INVX2
XFILL_0__1357_ vdd gnd FILL
XFILL_0__1288_ vdd gnd FILL
XFILL_3__1066_ vdd gnd FILL
XFILL_3__1135_ vdd gnd FILL
XFILL_0__1426_ vdd gnd FILL
X_1419_ _1599_/A _974_/B _981_/B _1604_/A _1425_/B vdd gnd AOI22X1
XFILL_1__1604_ vdd gnd FILL
XFILL_4__1313_ vdd gnd FILL
XFILL_4__1244_ vdd gnd FILL
XFILL_1__1535_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL_1__1466_ vdd gnd FILL
XFILL_2__926_ vdd gnd FILL
XFILL_2__857_ vdd gnd FILL
X_932_ _968_/A _953_/Q _932_/C _934_/B vdd gnd NAND3X1
X_863_ _867_/A _938_/Q _863_/C _939_/D vdd gnd OAI21X1
XFILL_2__1713_ vdd gnd FILL
XFILL_2__1575_ vdd gnd FILL
XFILL_2__1644_ vdd gnd FILL
XFILL_0__1211_ vdd gnd FILL
XFILL_0__1142_ vdd gnd FILL
XFILL_2__1009_ vdd gnd FILL
XFILL_0__1073_ vdd gnd FILL
X_1204_ _1231_/B _1231_/A _1211_/B vdd gnd OR2X2
XFILL_1__875_ vdd gnd FILL
XFILL_1__1320_ vdd gnd FILL
XFILL_1__1251_ vdd gnd FILL
X_1066_ _962_/A _1281_/B vdd gnd INVX1
X_1135_ _962_/B _1135_/B _1136_/A vdd gnd NAND2X1
XFILL_1__1182_ vdd gnd FILL
XFILL_3__1049_ vdd gnd FILL
XFILL_0__1409_ vdd gnd FILL
XFILL_3__1118_ vdd gnd FILL
XFILL_2__1360_ vdd gnd FILL
XFILL_4__1227_ vdd gnd FILL
XFILL_4__1158_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_4__1089_ vdd gnd FILL
XFILL_1__1518_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_2__909_ vdd gnd FILL
XFILL_0__893_ vdd gnd FILL
X_915_ _915_/A _915_/B _925_/A _916_/B vdd gnd OAI21X1
X_846_ _957_/A _960_/A _848_/A vdd gnd NOR2X1
XFILL_2__1627_ vdd gnd FILL
XFILL_4__871_ vdd gnd FILL
XFILL_2__1558_ vdd gnd FILL
XFILL_2__1489_ vdd gnd FILL
XFILL_3_BUFX2_insert12 vdd gnd FILL
XFILL_0__1125_ vdd gnd FILL
XFILL_0__1056_ vdd gnd FILL
X_1684_ _1684_/D vdd _1689_/R _1689_/CLK _1684_/Q vdd gnd DFFSR
XFILL_1__927_ vdd gnd FILL
XFILL_1__858_ vdd gnd FILL
XFILL_3__1598_ vdd gnd FILL
XFILL_3__1667_ vdd gnd FILL
XFILL_4__1012_ vdd gnd FILL
X_1049_ _985_/C _988_/A _1050_/C vdd gnd NAND2X1
XFILL_1__1234_ vdd gnd FILL
XFILL_1__1303_ vdd gnd FILL
X_1118_ _1138_/C _1118_/B _1118_/C _1139_/B vdd gnd AOI21X1
XFILL_1__1165_ vdd gnd FILL
XFILL_1__1096_ vdd gnd FILL
XFILL_4_CLKBUF1_insert4 vdd gnd FILL
XFILL_2__1412_ vdd gnd FILL
XFILL_2__1343_ vdd gnd FILL
XFILL_2__1274_ vdd gnd FILL
XFILL_0__876_ vdd gnd FILL
X_829_ _975_/A _936_/A vdd gnd INVX1
XFILL_3__1383_ vdd gnd FILL
XFILL_0__1674_ vdd gnd FILL
XFILL_3__1452_ vdd gnd FILL
XFILL_3__1521_ vdd gnd FILL
XFILL_4__923_ vdd gnd FILL
XFILL_4__854_ vdd gnd FILL
XFILL_0__1039_ vdd gnd FILL
XFILL_0__1108_ vdd gnd FILL
X_1598_ _1710_/Q _1604_/B _1600_/C vdd gnd NAND2X1
XFILL_4__1561_ vdd gnd FILL
XFILL_3__1719_ vdd gnd FILL
XFILL_4__1492_ vdd gnd FILL
XFILL_4__1630_ vdd gnd FILL
X_1667_ _1667_/A _1668_/A vdd gnd INVX1
XFILL_1__1217_ vdd gnd FILL
XFILL_1__1148_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_3__872_ vdd gnd FILL
XFILL_2__1326_ vdd gnd FILL
XFILL_2__1257_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
XFILL_0__859_ vdd gnd FILL
XFILL_2__1188_ vdd gnd FILL
XFILL_2_BUFX2_insert2 vdd gnd FILL
X_1383_ _1693_/Q _1383_/B _1421_/B _1694_/Q _1420_/A vdd gnd AOI22X1
X_1452_ _1523_/A _1473_/B _1489_/B vdd gnd NOR2X1
X_1521_ _1521_/A _1573_/B _1522_/B vdd gnd NOR2X1
XFILL_3__1366_ vdd gnd FILL
XFILL_0__1657_ vdd gnd FILL
XFILL_3__1435_ vdd gnd FILL
XFILL_3__1504_ vdd gnd FILL
XFILL_4__906_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_2__890_ vdd gnd FILL
XFILL_0__1588_ vdd gnd FILL
XFILL_3__1297_ vdd gnd FILL
X_1719_ _1723_/A rgb[4] vdd gnd BUFX2
XFILL_4__1613_ vdd gnd FILL
XFILL_4__1475_ vdd gnd FILL
XFILL_4__1544_ vdd gnd FILL
XFILL_2__1111_ vdd gnd FILL
XFILL_2__1042_ vdd gnd FILL
XFILL_3__924_ vdd gnd FILL
XFILL_3__1220_ vdd gnd FILL
XFILL_3__855_ vdd gnd FILL
XFILL_0__1511_ vdd gnd FILL
XFILL_3__1151_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
XFILL_3__1082_ vdd gnd FILL
XFILL_2__1309_ vdd gnd FILL
X_1504_ _1504_/A _1524_/A _1524_/B _1505_/B vdd gnd NAND3X1
X_1366_ _1674_/C _1401_/B _1367_/C vdd gnd NAND2X1
XFILL_1__1551_ vdd gnd FILL
X_1435_ _1473_/B _1435_/B _1435_/C _1680_/D vdd gnd OAI21X1
XFILL_1__1620_ vdd gnd FILL
XFILL_4__1191_ vdd gnd FILL
XFILL_3__1349_ vdd gnd FILL
X_1297_ _1297_/A _1297_/B _1300_/A vdd gnd NOR2X1
XFILL_1__1482_ vdd gnd FILL
XFILL_3__1418_ vdd gnd FILL
XFILL_4__1260_ vdd gnd FILL
XFILL_2__873_ vdd gnd FILL
XFILL_2__1660_ vdd gnd FILL
XFILL_4__1527_ vdd gnd FILL
XFILL_2__1591_ vdd gnd FILL
XFILL_4__1458_ vdd gnd FILL
XFILL_4__1389_ vdd gnd FILL
XFILL103650x11850 vdd gnd FILL
XFILL_2__1025_ vdd gnd FILL
XFILL103350x46950 vdd gnd FILL
XFILL103950x93750 vdd gnd FILL
X_1220_ _968_/A _1599_/A _1224_/B vdd gnd NAND2X1
XFILL_3__907_ vdd gnd FILL
X_1151_ _1317_/B _1151_/B _1317_/A _1348_/B vdd gnd NAND3X1
XFILL_3__838_ vdd gnd FILL
XFILL_1__891_ vdd gnd FILL
XFILL_1__960_ vdd gnd FILL
XFILL_3__1203_ vdd gnd FILL
XFILL_0__1425_ vdd gnd FILL
X_1082_ _1684_/Q _1523_/A vdd gnd INVX2
XFILL_0__1356_ vdd gnd FILL
XFILL_3__1065_ vdd gnd FILL
XFILL_3__1134_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
X_1349_ _978_/A _1400_/C _1350_/B vdd gnd NAND2X1
XFILL_4__1243_ vdd gnd FILL
XFILL_1__1603_ vdd gnd FILL
XFILL_1__1534_ vdd gnd FILL
XFILL_4__1312_ vdd gnd FILL
X_1418_ _1418_/A _1432_/A _1677_/B _1435_/B vdd gnd AOI21X1
XFILL_4__1174_ vdd gnd FILL
XFILL_2__925_ vdd gnd FILL
XFILL_1__1396_ vdd gnd FILL
XFILL_1__1465_ vdd gnd FILL
XFILL_2__856_ vdd gnd FILL
X_931_ _938_/D _931_/B _968_/A _935_/C vdd gnd OAI21X1
X_862_ _867_/A _938_/Q _931_/B _863_/C vdd gnd NAND3X1
XFILL_2__1712_ vdd gnd FILL
XFILL_2__1643_ vdd gnd FILL
XFILL_2__1574_ vdd gnd FILL
XFILL_0__1210_ vdd gnd FILL
XFILL_2__1008_ vdd gnd FILL
XFILL103350x58650 vdd gnd FILL
XFILL_0__1141_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
X_1203_ _1210_/C _1209_/A _1231_/B vdd gnd OR2X2
XFILL_1__874_ vdd gnd FILL
X_1134_ _965_/A _1134_/B _1134_/C _1134_/D _1136_/B vdd gnd AOI22X1
XFILL_1__1181_ vdd gnd FILL
XFILL_1__1250_ vdd gnd FILL
X_1065_ _965_/A _1530_/A vdd gnd INVX1
XFILL_3__1117_ vdd gnd FILL
XFILL_0__1408_ vdd gnd FILL
XFILL_3__1048_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
XFILL_4__1226_ vdd gnd FILL
XFILL_1__1517_ vdd gnd FILL
XFILL_2__1290_ vdd gnd FILL
XFILL_2__908_ vdd gnd FILL
XFILL_4__1157_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_0__892_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_4__1088_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_2__839_ vdd gnd FILL
X_914_ _951_/Q _919_/C _928_/B vdd gnd NAND2X1
X_845_ _845_/A _891_/A _894_/A _864_/B vdd gnd AOI21X1
XFILL103650x35250 vdd gnd FILL
XFILL_2__1626_ vdd gnd FILL
XFILL_4__870_ vdd gnd FILL
XFILL_2__1557_ vdd gnd FILL
XFILL_2__1488_ vdd gnd FILL
XFILL_0__1055_ vdd gnd FILL
XFILL_3_BUFX2_insert13 vdd gnd FILL
XFILL_0__1124_ vdd gnd FILL
X_1683_ _1683_/D vdd _1708_/R _1689_/CLK _1683_/Q vdd gnd DFFSR
XFILL_3__1666_ vdd gnd FILL
XFILL_1__926_ vdd gnd FILL
XFILL_1__857_ vdd gnd FILL
XFILL_3__1597_ vdd gnd FILL
X_1117_ _1117_/A _1117_/B _1117_/C _1118_/C vdd gnd OAI21X1
XFILL_1__1164_ vdd gnd FILL
X_1048_ _1048_/A _1048_/B _1060_/A vdd gnd OR2X2
XFILL_4__1011_ vdd gnd FILL
XFILL_1__1233_ vdd gnd FILL
XFILL_4__999_ vdd gnd FILL
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1095_ vdd gnd FILL
XFILL_2__1411_ vdd gnd FILL
XFILL_4_CLKBUF1_insert5 vdd gnd FILL
XFILL_4__1209_ vdd gnd FILL
XFILL_2__1342_ vdd gnd FILL
XFILL_2__1273_ vdd gnd FILL
XFILL_0__875_ vdd gnd FILL
XFILL_3__1520_ vdd gnd FILL
X_828_ _956_/Q _937_/A vdd gnd INVX1
XFILL_3__1382_ vdd gnd FILL
XFILL_2__1609_ vdd gnd FILL
XFILL_0__1673_ vdd gnd FILL
XFILL_3__1451_ vdd gnd FILL
XFILL_4__853_ vdd gnd FILL
XFILL_4__922_ vdd gnd FILL
XFILL_0__1038_ vdd gnd FILL
XFILL102150x62550 vdd gnd FILL
XFILL_0__1107_ vdd gnd FILL
X_1666_ _1666_/A _1673_/A _1666_/C _1668_/B vdd gnd OAI21X1
XFILL_3__1718_ vdd gnd FILL
XFILL_1__909_ vdd gnd FILL
X_1597_ _1597_/A _1599_/B _1597_/C _1604_/B vdd gnd OAI21X1
XFILL_3__1649_ vdd gnd FILL
XFILL_4__1560_ vdd gnd FILL
XFILL_4__1491_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_1__1147_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_3__871_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
XFILL_2__1325_ vdd gnd FILL
XFILL_2__1256_ vdd gnd FILL
XFILL_0__927_ vdd gnd FILL
XFILL_0__858_ vdd gnd FILL
X_1520_ _1520_/A _1546_/B _1520_/C _1683_/D vdd gnd OAI21X1
XFILL_2_BUFX2_insert3 vdd gnd FILL
X_1382_ _1382_/A _1382_/B _1382_/C _1420_/B vdd gnd NAND3X1
XFILL_3__1503_ vdd gnd FILL
X_1451_ _1681_/Q _1678_/Q _1504_/A vdd gnd XOR2X1
XFILL_0__1725_ vdd gnd FILL
XFILL_3__1365_ vdd gnd FILL
XFILL_0__1587_ vdd gnd FILL
XFILL_0__1656_ vdd gnd FILL
XFILL_3__1434_ vdd gnd FILL
XFILL_3__1296_ vdd gnd FILL
XFILL_4__836_ vdd gnd FILL
XFILL_4__905_ vdd gnd FILL
XFILL_1__1001_ vdd gnd FILL
X_1718_ _1724_/A rgb[3] vdd gnd BUFX2
XFILL_4__1612_ vdd gnd FILL
X_1649_ _1649_/A _1655_/C _1656_/A _1650_/C vdd gnd NAND3X1
XFILL_4__1474_ vdd gnd FILL
XFILL_4__1543_ vdd gnd FILL
XFILL_2__1041_ vdd gnd FILL
XFILL_2__1110_ vdd gnd FILL
XFILL_3__923_ vdd gnd FILL
XFILL_3__854_ vdd gnd FILL
XFILL_3__1150_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_0__1510_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
XFILL_2__1308_ vdd gnd FILL
XFILL_3__1081_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
X_1503_ _1503_/A _1503_/B _1524_/A vdd gnd XOR2X1
X_1365_ _1365_/A _1365_/B _1367_/B vdd gnd OR2X2
X_1434_ _1680_/Q _1473_/B vdd gnd INVX2
XFILL_1__1550_ vdd gnd FILL
X_1296_ _1299_/A _1296_/B _1296_/C _1302_/B vdd gnd OAI21X1
XFILL_3__1348_ vdd gnd FILL
XFILL_4__1190_ vdd gnd FILL
XFILL_3__1417_ vdd gnd FILL
XFILL_3__1279_ vdd gnd FILL
XFILL_0__1639_ vdd gnd FILL
XFILL_1__1481_ vdd gnd FILL
XFILL_2__872_ vdd gnd FILL
XFILL_2__1590_ vdd gnd FILL
XFILL_4__1526_ vdd gnd FILL
XFILL_4__1388_ vdd gnd FILL
XFILL_4__1457_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
XFILL_3__837_ vdd gnd FILL
X_1150_ _1604_/A _1599_/A _1151_/B vdd gnd NOR2X1
XFILL_3__906_ vdd gnd FILL
XFILL_1__890_ vdd gnd FILL
XFILL_0_CLKBUF1_insert10 vdd gnd FILL
XFILL_0__1355_ vdd gnd FILL
XFILL_3__1202_ vdd gnd FILL
XFILL_0__1424_ vdd gnd FILL
X_1081_ _1688_/Q _1544_/A vdd gnd INVX2
XFILL_3__1133_ vdd gnd FILL
XFILL_3__1064_ vdd gnd FILL
XFILL_0__1286_ vdd gnd FILL
X_1417_ _1417_/A _1417_/B _1417_/C _1418_/A vdd gnd OAI21X1
X_1348_ _979_/C _1348_/B _1348_/C _1350_/A vdd gnd NAND3X1
XFILL_4__1242_ vdd gnd FILL
XFILL_1__1602_ vdd gnd FILL
XFILL_1__1533_ vdd gnd FILL
XFILL_1__1464_ vdd gnd FILL
X_1279_ _1537_/A _962_/B _1291_/A _1283_/A vdd gnd AOI21X1
XFILL_4__1311_ vdd gnd FILL
XFILL_2__924_ vdd gnd FILL
XFILL_1__1395_ vdd gnd FILL
XFILL_4__1173_ vdd gnd FILL
XFILL_2__855_ vdd gnd FILL
X_930_ _935_/A _930_/B _930_/C _953_/D vdd gnd OAI21X1
X_861_ _964_/A _864_/B _931_/B vdd gnd NOR2X1
XFILL_2__1711_ vdd gnd FILL
XFILL_4__1509_ vdd gnd FILL
XFILL_2__1642_ vdd gnd FILL
XFILL_2__1573_ vdd gnd FILL
XFILL_2__1007_ vdd gnd FILL
XFILL_0__1140_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
X_1202_ _1693_/Q _1512_/B _1209_/A vdd gnd NOR2X1
XFILL_1__873_ vdd gnd FILL
X_1064_ _962_/B _961_/B _1064_/C _1069_/A vdd gnd NAND3X1
X_1133_ _1133_/A _1530_/A _1133_/C _1134_/D vdd gnd AOI21X1
XFILL_0__1338_ vdd gnd FILL
XFILL_1__1180_ vdd gnd FILL
XFILL_3__1047_ vdd gnd FILL
XFILL_0__1407_ vdd gnd FILL
XFILL_3__1116_ vdd gnd FILL
XFILL_0__1269_ vdd gnd FILL
XFILL_4__1225_ vdd gnd FILL
XFILL_4__1156_ vdd gnd FILL
XFILL_1__1516_ vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_2__907_ vdd gnd FILL
XFILL_2__838_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
XFILL_0__891_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL_4__1087_ vdd gnd FILL
X_913_ _925_/C _919_/C vdd gnd INVX1
XFILL103950x19650 vdd gnd FILL
X_844_ _961_/A _894_/A vdd gnd INVX1
XFILL_2__1556_ vdd gnd FILL
XFILL_2__1625_ vdd gnd FILL
XFILL_2__1487_ vdd gnd FILL
XFILL_0__1054_ vdd gnd FILL
X_1682_ _1682_/D vdd _1702_/R _1702_/CLK _1682_/Q vdd gnd DFFSR
XFILL_3_BUFX2_insert14 vdd gnd FILL
XFILL_0__1123_ vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_3__1665_ vdd gnd FILL
XFILL_1__856_ vdd gnd FILL
X_1047_ _998_/A _1512_/B _997_/A _997_/B _1048_/B vdd gnd OAI22X1
XFILL_4__1010_ vdd gnd FILL
XFILL_3__1596_ vdd gnd FILL
X_1116_ _1293_/B _1394_/A _1117_/C vdd gnd NAND2X1
XFILL_1__1301_ vdd gnd FILL
XFILL_1__1163_ vdd gnd FILL
XFILL_1__1232_ vdd gnd FILL
XFILL_4__998_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL_4_CLKBUF1_insert6 vdd gnd FILL
XFILL_2__1410_ vdd gnd FILL
XFILL_2__1341_ vdd gnd FILL
XFILL_4__1208_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_4__1139_ vdd gnd FILL
XFILL_0__874_ vdd gnd FILL
XFILL_3__1450_ vdd gnd FILL
XFILL_4__921_ vdd gnd FILL
XFILL_3__1381_ vdd gnd FILL
XFILL_2__1608_ vdd gnd FILL
XFILL_0__1672_ vdd gnd FILL
XFILL_2__1539_ vdd gnd FILL
XFILL_4__852_ vdd gnd FILL
XFILL102750x11850 vdd gnd FILL
XFILL_0__1037_ vdd gnd FILL
X_1596_ _1696_/Q _1710_/Q _1597_/C vdd gnd NAND2X1
XFILL_0__1106_ vdd gnd FILL
X_1665_ _1666_/C _1667_/A _1665_/C _1669_/C vdd gnd NAND3X1
XFILL_1__908_ vdd gnd FILL
XFILL_3__1648_ vdd gnd FILL
XFILL_3__1579_ vdd gnd FILL
XFILL_3__1717_ vdd gnd FILL
XFILL_4__1490_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL_1__839_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_3__870_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_2__1186_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
XFILL_2__1255_ vdd gnd FILL
XFILL_0__857_ vdd gnd FILL
X_1450_ _1582_/A _1582_/B _1681_/Q _1505_/C vdd gnd OAI21X1
XFILL_0__1724_ vdd gnd FILL
X_1381_ _1381_/A _1381_/B _1381_/C _1382_/C vdd gnd NAND3X1
XFILL_3__999_ vdd gnd FILL
XFILL_3__1433_ vdd gnd FILL
XFILL_3__1502_ vdd gnd FILL
XFILL_4__904_ vdd gnd FILL
XFILL_3__1364_ vdd gnd FILL
XFILL_0__1655_ vdd gnd FILL
XFILL_3__1295_ vdd gnd FILL
XFILL_0__1586_ vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
XFILL_4__835_ vdd gnd FILL
X_1648_ _1648_/A _1650_/A _1670_/B _1703_/D vdd gnd MUX2X1
X_1579_ _1592_/A _1591_/A _1580_/C vdd gnd OR2X2
XFILL_4__1542_ vdd gnd FILL
X_1717_ _1721_/A rgb[2] vdd gnd BUFX2
XFILL_4__1611_ vdd gnd FILL
XFILL_4__1473_ vdd gnd FILL
XFILL_2__1040_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_3__853_ vdd gnd FILL
XFILL_3__922_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_3__1080_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
XFILL_2__1307_ vdd gnd FILL
XFILL_2__1169_ vdd gnd FILL
XFILL_0__909_ vdd gnd FILL
XFILL_2__1238_ vdd gnd FILL
X_1433_ _1433_/A _1435_/B _1435_/C _1679_/D vdd gnd OAI21X1
X_1502_ _1689_/Q _1680_/Q _1503_/B vdd gnd XOR2X1
XFILL_3__1416_ vdd gnd FILL
X_1364_ _1364_/A _1364_/B _1364_/C _1365_/B vdd gnd NAND3X1
X_1295_ _1295_/A _1295_/B _1295_/C _1296_/C vdd gnd AOI21X1
XFILL_1__1480_ vdd gnd FILL
XFILL_3__1347_ vdd gnd FILL
XFILL_2__871_ vdd gnd FILL
XFILL_0__1569_ vdd gnd FILL
XFILL_3__1278_ vdd gnd FILL
XFILL_0__1638_ vdd gnd FILL
XFILL_4__1525_ vdd gnd FILL
XFILL_4__1387_ vdd gnd FILL
XFILL_4__1456_ vdd gnd FILL
XFILL_2__1023_ vdd gnd FILL
XFILL_3__905_ vdd gnd FILL
XFILL_3__836_ vdd gnd FILL
X_1080_ _967_/A _967_/B _1080_/C _1080_/D _1306_/A vdd gnd AOI22X1
XFILL_0__1354_ vdd gnd FILL
XFILL_3__1201_ vdd gnd FILL
XFILL_0__1423_ vdd gnd FILL
XFILL_3__1063_ vdd gnd FILL
XFILL_3__1132_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
X_1416_ _1416_/A _1416_/B _1416_/C _1417_/B vdd gnd AOI21X1
X_1347_ _1347_/A _1347_/B _1358_/A vdd gnd AND2X2
XFILL_1__1601_ vdd gnd FILL
XFILL_4__1172_ vdd gnd FILL
XFILL_4__1241_ vdd gnd FILL
XFILL_1__1532_ vdd gnd FILL
XFILL_1__1463_ vdd gnd FILL
X_1278_ _1686_/Q _1281_/B _1291_/A vdd gnd NOR2X1
XFILL_4__1310_ vdd gnd FILL
XFILL_1__1394_ vdd gnd FILL
XFILL_2__923_ vdd gnd FILL
XFILL_2__854_ vdd gnd FILL
X_860_ _960_/A _867_/A vdd gnd INVX1
XFILL_4__1439_ vdd gnd FILL
XFILL_2__1641_ vdd gnd FILL
XFILL_2__1572_ vdd gnd FILL
XFILL_4__1508_ vdd gnd FILL
XFILL_2__1006_ vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
X_1201_ _951_/Q _1573_/A _1210_/C vdd gnd NOR2X1
XFILL_1__872_ vdd gnd FILL
X_989_ _992_/B _989_/B _996_/B vdd gnd NOR2X1
X_1063_ _961_/A _964_/A _1064_/C vdd gnd NOR2X1
X_1132_ _1683_/Q _1132_/B _1289_/A _1133_/C vdd gnd OAI21X1
XFILL_0__1406_ vdd gnd FILL
XFILL_3__1046_ vdd gnd FILL
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
XFILL_3__1115_ vdd gnd FILL
XFILL_0__1199_ vdd gnd FILL
XFILL_4__1224_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_4__1155_ vdd gnd FILL
XFILL_1__1515_ vdd gnd FILL
XFILL_2__837_ vdd gnd FILL
XFILL_2__906_ vdd gnd FILL
XFILL_0__890_ vdd gnd FILL
XFILL_4__1086_ vdd gnd FILL
X_912_ _938_/D _931_/B _951_/Q _917_/C vdd gnd OAI21X1
X_843_ _965_/A _843_/B _961_/A _849_/C vdd gnd OAI21X1
XFILL_2__1555_ vdd gnd FILL
XFILL_2__1486_ vdd gnd FILL
XFILL_2__1624_ vdd gnd FILL
XFILL_0__1122_ vdd gnd FILL
XFILL_0__1053_ vdd gnd FILL
XFILL_3_BUFX2_insert15 vdd gnd FILL
X_1681_ _1681_/D vdd _1708_/R _1709_/CLK _1681_/Q vdd gnd DFFSR
XFILL_1__924_ vdd gnd FILL
XFILL_1__855_ vdd gnd FILL
XFILL_3__1595_ vdd gnd FILL
XFILL_3__1664_ vdd gnd FILL
XFILL_1__1231_ vdd gnd FILL
X_1046_ _951_/Q _1512_/B vdd gnd INVX1
X_1115_ _1276_/D _1427_/B _1117_/A vdd gnd NAND2X1
XFILL_1__1300_ vdd gnd FILL
XFILL_1__1162_ vdd gnd FILL
XFILL_4__997_ vdd gnd FILL
XFILL_3__1029_ vdd gnd FILL
XFILL_1__1093_ vdd gnd FILL
XFILL_4_CLKBUF1_insert7 vdd gnd FILL
XFILL_2__1340_ vdd gnd FILL
XFILL_4__1207_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_4__1069_ vdd gnd FILL
XFILL_2__1271_ vdd gnd FILL
XFILL_4__1138_ vdd gnd FILL
XFILL_0__873_ vdd gnd FILL
XFILL_2__1607_ vdd gnd FILL
XFILL_0__1671_ vdd gnd FILL
XFILL_4__920_ vdd gnd FILL
XFILL_3__1380_ vdd gnd FILL
XFILL_2__1469_ vdd gnd FILL
XFILL_2__1538_ vdd gnd FILL
XFILL_4__851_ vdd gnd FILL
XFILL_0__1105_ vdd gnd FILL
XFILL_0__1036_ vdd gnd FILL
XFILL_3__1716_ vdd gnd FILL
X_1595_ _1599_/A _1595_/B _1595_/C _1595_/D _1696_/D vdd gnd OAI22X1
X_1664_ _1671_/C _979_/C _1667_/A vdd gnd XOR2X1
XFILL_1__907_ vdd gnd FILL
XFILL_1__838_ vdd gnd FILL
XFILL_3__1647_ vdd gnd FILL
XFILL_3__1578_ vdd gnd FILL
XFILL_1__1214_ vdd gnd FILL
X_1029_ _980_/B _1674_/C _1618_/B vdd gnd XOR2X1
XFILL_1__1145_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_2__1323_ vdd gnd FILL
XFILL_2__1185_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
XFILL_2__1254_ vdd gnd FILL
XFILL_0__856_ vdd gnd FILL
XFILL103050x70350 vdd gnd FILL
X_1380_ _1692_/Q _994_/A _994_/B _1381_/C vdd gnd NAND3X1
XFILL_3__1363_ vdd gnd FILL
XFILL_0__1654_ vdd gnd FILL
XFILL_3__1501_ vdd gnd FILL
XFILL_0__1723_ vdd gnd FILL
XFILL_3__998_ vdd gnd FILL
XFILL_3__1432_ vdd gnd FILL
XFILL_4__903_ vdd gnd FILL
XFILL_4__834_ vdd gnd FILL
XFILL_0__1585_ vdd gnd FILL
XFILL_3__1294_ vdd gnd FILL
X_1716_ _1724_/A rgb[11] vdd gnd BUFX2
XFILL_0__1019_ vdd gnd FILL
X_1647_ _1656_/A _1654_/B _1648_/A vdd gnd XOR2X1
X_1578_ _1591_/A _1592_/A _1583_/C vdd gnd NAND2X1
XFILL_4__1610_ vdd gnd FILL
XFILL_4__1472_ vdd gnd FILL
XFILL_4__1541_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_3__921_ vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_3__852_ vdd gnd FILL
XFILL_2__1237_ vdd gnd FILL
XFILL_2__1306_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
XFILL_0__908_ vdd gnd FILL
XFILL_2__1168_ vdd gnd FILL
XFILL_0__839_ vdd gnd FILL
XFILL_2__1099_ vdd gnd FILL
X_1363_ _1363_/A _1376_/B _1364_/B vdd gnd NOR2X1
X_1501_ _1501_/A _1501_/B _1501_/C _1503_/A vdd gnd AOI21X1
X_1432_ _1432_/A _1675_/B _1432_/C _1435_/C vdd gnd NAND3X1
XFILL_3__1346_ vdd gnd FILL
XFILL_3__1415_ vdd gnd FILL
XFILL_0__1637_ vdd gnd FILL
X_1294_ _1294_/A _1294_/B _1294_/C _1295_/C vdd gnd OAI21X1
XFILL_2__870_ vdd gnd FILL
XFILL_0__1568_ vdd gnd FILL
XFILL_0__1499_ vdd gnd FILL
XFILL_3__1277_ vdd gnd FILL
XFILL_4__1524_ vdd gnd FILL
XFILL_4__1455_ vdd gnd FILL
XFILL_4__1386_ vdd gnd FILL
XFILL_1__1677_ vdd gnd FILL
XFILL_2__1022_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL_3__904_ vdd gnd FILL
XFILL_3__835_ vdd gnd FILL
XFILL_3__1200_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_3__1062_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
XFILL_3__1131_ vdd gnd FILL
X_1346_ _1358_/C _1416_/B _1346_/C _1357_/C vdd gnd NAND3X1
X_1415_ _1415_/A _1415_/B _1416_/C vdd gnd NAND2X1
XFILL_1__1531_ vdd gnd FILL
XFILL_1__1600_ vdd gnd FILL
XFILL_3__1329_ vdd gnd FILL
XFILL_2__922_ vdd gnd FILL
XFILL_4__1171_ vdd gnd FILL
XFILL_4__1240_ vdd gnd FILL
X_1277_ _1277_/A _1277_/B _1295_/A vdd gnd NOR2X1
XFILL_1__1462_ vdd gnd FILL
XFILL_1__1393_ vdd gnd FILL
XFILL_2__853_ vdd gnd FILL
XFILL_2__1640_ vdd gnd FILL
XFILL_4__1438_ vdd gnd FILL
XFILL_2__1571_ vdd gnd FILL
XFILL_4__1507_ vdd gnd FILL
XFILL_4__1369_ vdd gnd FILL
XFILL_2__1005_ vdd gnd FILL
X_1200_ _1248_/A _1248_/B _1231_/A vdd gnd OR2X2
X_988_ _988_/A _989_/B vdd gnd INVX1
XFILL_1__871_ vdd gnd FILL
XFILL_0__1405_ vdd gnd FILL
X_1062_ _1707_/Q _1513_/A _1062_/C _1072_/B vdd gnd OAI21X1
X_1131_ _1683_/Q _959_/B _1289_/A vdd gnd NAND2X1
XFILL_0__1336_ vdd gnd FILL
XFILL_3__1045_ vdd gnd FILL
XFILL_0__1267_ vdd gnd FILL
XFILL_3__1114_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
X_1329_ _971_/A _1411_/B _1329_/C _1358_/C vdd gnd AOI21X1
XFILL_1__1514_ vdd gnd FILL
XFILL_2__905_ vdd gnd FILL
XFILL_4__1154_ vdd gnd FILL
XFILL_1__1376_ vdd gnd FILL
XFILL_1__1445_ vdd gnd FILL
XFILL_4__1085_ vdd gnd FILL
XFILL_2__836_ vdd gnd FILL
X_911_ _935_/A _911_/B _911_/C _950_/D vdd gnd OAI21X1
X_842_ _961_/A _891_/A _845_/A _843_/B vdd gnd NAND3X1
XFILL_2__1623_ vdd gnd FILL
XFILL_2__1485_ vdd gnd FILL
XFILL_2__1554_ vdd gnd FILL
XFILL_0__1052_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
X_1680_ _1680_/D vdd _1702_/R _1702_/CLK _1680_/Q vdd gnd DFFSR
XFILL_1__923_ vdd gnd FILL
XFILL_1__854_ vdd gnd FILL
XFILL_3__1594_ vdd gnd FILL
XFILL_3__1663_ vdd gnd FILL
X_1114_ _961_/B _1276_/D vdd gnd INVX1
XFILL_1__1161_ vdd gnd FILL
XFILL_1__1230_ vdd gnd FILL
X_1045_ _998_/Y _951_/Q _997_/Y _1048_/A vdd gnd OAI21X1
XFILL_4__996_ vdd gnd FILL
XFILL_0__1319_ vdd gnd FILL
XFILL_3__1028_ vdd gnd FILL
XFILL_1__1092_ vdd gnd FILL
XFILL_4_CLKBUF1_insert8 vdd gnd FILL
XFILL_4__1206_ vdd gnd FILL
XFILL_2__1270_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_0__872_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_4__1068_ vdd gnd FILL
XFILL_4__1137_ vdd gnd FILL
XFILL_2__1606_ vdd gnd FILL
XFILL_0__1670_ vdd gnd FILL
XFILL_4__850_ vdd gnd FILL
XFILL_2__1468_ vdd gnd FILL
XFILL_2__1537_ vdd gnd FILL
XFILL_2__1399_ vdd gnd FILL
XFILL_0__1035_ vdd gnd FILL
X_1663_ _1663_/A _1670_/B _1663_/C _1705_/D vdd gnd OAI21X1
XFILL_0__1104_ vdd gnd FILL
X_1594_ _1597_/A _1599_/B _1602_/C _1595_/C vdd gnd OAI21X1
XFILL_3__1715_ vdd gnd FILL
XFILL_1__837_ vdd gnd FILL
XFILL_1__906_ vdd gnd FILL
XFILL_3__1577_ vdd gnd FILL
XFILL_3__1646_ vdd gnd FILL
XFILL_1__1213_ vdd gnd FILL
XFILL_1__1144_ vdd gnd FILL
XFILL_4__979_ vdd gnd FILL
X_1028_ _1707_/Q _1674_/C vdd gnd INVX2
XFILL_1__1075_ vdd gnd FILL
XFILL_2__1322_ vdd gnd FILL
XFILL_2__1253_ vdd gnd FILL
XFILL_2__1184_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_0__855_ vdd gnd FILL
XFILL_3__997_ vdd gnd FILL
XFILL_3__1500_ vdd gnd FILL
XFILL103050x89850 vdd gnd FILL
XFILL_0__1722_ vdd gnd FILL
XFILL_3__1362_ vdd gnd FILL
XFILL_0__1653_ vdd gnd FILL
XFILL_0__1584_ vdd gnd FILL
XFILL_3__1431_ vdd gnd FILL
XFILL_4__833_ vdd gnd FILL
XFILL_4__902_ vdd gnd FILL
XFILL_3__1293_ vdd gnd FILL
XFILL_0__1018_ vdd gnd FILL
X_1715_ _1721_/A rgb[10] vdd gnd BUFX2
X_1646_ _1646_/A _1646_/B _1646_/C _1656_/A vdd gnd OAI21X1
X_1577_ _1577_/A _1577_/B _1577_/C _1592_/A vdd gnd OAI21X1
XFILL_4__1471_ vdd gnd FILL
XFILL_4__1540_ vdd gnd FILL
XFILL_3__1629_ vdd gnd FILL
XFILL_1__1127_ vdd gnd FILL
XFILL_3__920_ vdd gnd FILL
XFILL_3__851_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_4__1669_ vdd gnd FILL
XFILL_2__1236_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL103650x31350 vdd gnd FILL
XFILL_0__907_ vdd gnd FILL
XFILL_0__838_ vdd gnd FILL
XFILL103350x66450 vdd gnd FILL
X_1500_ _1500_/A _1500_/B _1501_/B vdd gnd NOR2X1
XFILL_2__1098_ vdd gnd FILL
X_1362_ _1549_/A _999_/Y _1376_/B vdd gnd NOR2X1
X_1293_ _1688_/Q _1293_/B _1294_/B vdd gnd NOR2X1
X_1431_ _1677_/B _1675_/B vdd gnd INVX1
XFILL_3__1414_ vdd gnd FILL
XFILL_3__1345_ vdd gnd FILL
XFILL_0__1567_ vdd gnd FILL
XFILL_0__1636_ vdd gnd FILL
XFILL_3__1276_ vdd gnd FILL
XFILL_0__1498_ vdd gnd FILL
X_1629_ _1629_/A _984_/B _1674_/B _1700_/D vdd gnd MUX2X1
XFILL_4__1385_ vdd gnd FILL
XFILL_1__1676_ vdd gnd FILL
XFILL_4__1454_ vdd gnd FILL
XFILL_4__1523_ vdd gnd FILL
XFILL_2__1021_ vdd gnd FILL
XFILL_2__998_ vdd gnd FILL
XFILL_3__903_ vdd gnd FILL
XFILL_3__834_ vdd gnd FILL
XFILL103650x43050 vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_3__1130_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
XFILL_2__1219_ vdd gnd FILL
XFILL_3__1061_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
X_1414_ _1414_/A _1414_/B _1414_/C _1416_/A vdd gnd NOR3X1
X_1345_ _1345_/A _1345_/B _1345_/C _1416_/B vdd gnd OAI21X1
XFILL_1__1530_ vdd gnd FILL
X_1276_ _1688_/Q _1293_/B _1687_/Q _1276_/D _1277_/A vdd gnd OAI22X1
XFILL_3__1328_ vdd gnd FILL
XFILL_2__921_ vdd gnd FILL
XFILL_4__1170_ vdd gnd FILL
XFILL_3__1259_ vdd gnd FILL
XFILL_1__1461_ vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_0__1619_ vdd gnd FILL
XFILL_2__852_ vdd gnd FILL
XFILL_4__1437_ vdd gnd FILL
XFILL_4__1368_ vdd gnd FILL
XFILL_2__1570_ vdd gnd FILL
XFILL_1__1659_ vdd gnd FILL
XFILL_4__1506_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
XFILL_4__1299_ vdd gnd FILL
X_987_ _993_/A _987_/B _988_/A vdd gnd NAND2X1
XFILL_1__870_ vdd gnd FILL
X_1130_ _1132_/B _1260_/A _1130_/C _1134_/C vdd gnd NAND3X1
XFILL_0__1404_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
X_1061_ _1061_/A _1061_/B _1062_/C vdd gnd NAND2X1
XFILL_3__1113_ vdd gnd FILL
XFILL_0__1197_ vdd gnd FILL
XFILL_3__1044_ vdd gnd FILL
XFILL_0__1266_ vdd gnd FILL
X_1328_ _1412_/B _1412_/A _1413_/B _1329_/C vdd gnd NAND3X1
XFILL_4__1222_ vdd gnd FILL
XFILL_1__1513_ vdd gnd FILL
XFILL_1__1444_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
X_1259_ _1297_/A _1297_/B _1259_/C _1262_/A vdd gnd OAI21X1
XFILL_2__835_ vdd gnd FILL
XFILL_4__1153_ vdd gnd FILL
XFILL_2__904_ vdd gnd FILL
XFILL_1__1375_ vdd gnd FILL
XFILL_4__1084_ vdd gnd FILL
X_910_ _925_/C _910_/B _934_/A _911_/B vdd gnd NAND3X1
X_841_ _962_/A _962_/B _845_/A vdd gnd NOR2X1
XFILL_2__1622_ vdd gnd FILL
XFILL_2__1553_ vdd gnd FILL
XFILL_2__1484_ vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_0__1120_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
XFILL_3__1662_ vdd gnd FILL
XFILL_1__853_ vdd gnd FILL
X_1044_ _1044_/A _1057_/B _1061_/A vdd gnd NOR2X1
XFILL_3__1593_ vdd gnd FILL
X_1113_ _1293_/B _1394_/A _1117_/B vdd gnd NOR2X1
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1160_ vdd gnd FILL
XFILL_4__995_ vdd gnd FILL
XFILL_1__1091_ vdd gnd FILL
XFILL_0__1249_ vdd gnd FILL
XFILL_3__1027_ vdd gnd FILL
XFILL_4_CLKBUF1_insert9 vdd gnd FILL
XFILL_4__1205_ vdd gnd FILL
XFILL_4__1136_ vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
XFILL_0__871_ vdd gnd FILL
XFILL_4__1067_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_2__1605_ vdd gnd FILL
XFILL_2__1536_ vdd gnd FILL
XFILL_2__1398_ vdd gnd FILL
XFILL_2__1467_ vdd gnd FILL
XFILL_0__1034_ vdd gnd FILL
X_1662_ _1665_/C _1662_/B _1670_/B _1663_/C vdd gnd NAND3X1
XFILL_0__1103_ vdd gnd FILL
XFILL_3__1714_ vdd gnd FILL
XFILL_1__905_ vdd gnd FILL
X_1593_ _1599_/B _1597_/A _1595_/D vdd gnd AND2X2
XFILL_3__1645_ vdd gnd FILL
XFILL_1__836_ vdd gnd FILL
X_1027_ _1079_/C _1074_/B vdd gnd INVX1
XFILL_3__1576_ vdd gnd FILL
XFILL_1__1212_ vdd gnd FILL
XFILL_4__978_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_1__1143_ vdd gnd FILL
XFILL_2__1183_ vdd gnd FILL
XFILL_2__1321_ vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL_4__1119_ vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
XFILL_0__854_ vdd gnd FILL
XFILL_3__996_ vdd gnd FILL
XFILL_0__1721_ vdd gnd FILL
XFILL_3__1361_ vdd gnd FILL
XFILL_4__901_ vdd gnd FILL
XFILL_0__1652_ vdd gnd FILL
XFILL_3__1430_ vdd gnd FILL
XFILL_0__1583_ vdd gnd FILL
XFILL_3__1292_ vdd gnd FILL
XFILL_2__1519_ vdd gnd FILL
XFILL_4__832_ vdd gnd FILL
X_1714_ _1724_/A rgb[1] vdd gnd BUFX2
XFILL_0__1017_ vdd gnd FILL
X_1576_ _1576_/A _1576_/B _1591_/A vdd gnd NOR2X1
X_1645_ _1645_/A _1645_/B _1646_/B vdd gnd NAND2X1
XFILL_3__1559_ vdd gnd FILL
XFILL_4__1470_ vdd gnd FILL
XFILL_3__1628_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
XFILL_3__850_ vdd gnd FILL
XFILL_4__1668_ vdd gnd FILL
XFILL_2__1304_ vdd gnd FILL
XFILL_4__1599_ vdd gnd FILL
XFILL103950x15750 vdd gnd FILL
XFILL_2__1166_ vdd gnd FILL
XFILL_2__1235_ vdd gnd FILL
XFILL_0__906_ vdd gnd FILL
XFILL_0__837_ vdd gnd FILL
X_1430_ _1430_/A _1430_/B _1430_/C _1432_/C vdd gnd AOI21X1
XFILL_2__1097_ vdd gnd FILL
XFILL_3__1413_ vdd gnd FILL
X_1361_ _1361_/A _1361_/B _1361_/C _1365_/A vdd gnd NAND3X1
XFILL_3__979_ vdd gnd FILL
X_1292_ _1688_/Q _1293_/B _1294_/C vdd gnd NAND2X1
XFILL_3__1344_ vdd gnd FILL
XFILL_0__1566_ vdd gnd FILL
XFILL_0__1635_ vdd gnd FILL
XFILL_0__1497_ vdd gnd FILL
XFILL_3__1275_ vdd gnd FILL
X_1559_ _1559_/A _1677_/A _1564_/C vdd gnd NOR2X1
XFILL_4__1522_ vdd gnd FILL
X_1628_ _1628_/A _999_/Y _1629_/A vdd gnd XOR2X1
XFILL_4__1384_ vdd gnd FILL
XFILL_4__1453_ vdd gnd FILL
XFILL_1__1675_ vdd gnd FILL
XFILL_2__997_ vdd gnd FILL
XFILL_2__1020_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_3__833_ vdd gnd FILL
XFILL_3__902_ vdd gnd FILL
XFILL103950x27450 vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_3__1060_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_2__1218_ vdd gnd FILL
XFILL_2__1149_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
X_1413_ _1413_/A _1413_/B _1413_/C _1414_/C vdd gnd NAND3X1
X_1344_ _1344_/A _1344_/B _1345_/C vdd gnd NAND2X1
X_1275_ _1544_/A _961_/A _1294_/A _1277_/B vdd gnd OAI21X1
XFILL_1__1460_ vdd gnd FILL
XFILL_2__920_ vdd gnd FILL
XFILL_3__1327_ vdd gnd FILL
XFILL_3__1189_ vdd gnd FILL
XFILL_2__851_ vdd gnd FILL
XFILL_0__1618_ vdd gnd FILL
XFILL_3__1258_ vdd gnd FILL
XFILL_1__1391_ vdd gnd FILL
XFILL_0__1549_ vdd gnd FILL
XFILL_4__1505_ vdd gnd FILL
XFILL_4__1436_ vdd gnd FILL
XFILL_1__1589_ vdd gnd FILL
XFILL_1__1658_ vdd gnd FILL
XFILL_4__1298_ vdd gnd FILL
XFILL_2__1003_ vdd gnd FILL
XFILL103950x39150 vdd gnd FILL
X_986_ _986_/A _987_/B vdd gnd INVX1
X_1060_ _1060_/A _1060_/B _1061_/B vdd gnd NOR2X1
XFILL_3__1043_ vdd gnd FILL
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1403_ vdd gnd FILL
XFILL_3__1112_ vdd gnd FILL
XFILL_0__1196_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
X_1327_ _1655_/A _1327_/B _1327_/C _1413_/B vdd gnd NAND3X1
X_1189_ _953_/Q _1411_/B _1355_/B _968_/A _1193_/B vdd gnd AOI22X1
XFILL_4__1221_ vdd gnd FILL
XFILL_4__1152_ vdd gnd FILL
XFILL_1__1512_ vdd gnd FILL
XFILL_1__1443_ vdd gnd FILL
X_1258_ _1259_/C _1288_/C _1297_/B vdd gnd NAND2X1
XFILL_1__998_ vdd gnd FILL
XFILL_2__903_ vdd gnd FILL
XFILL_2__834_ vdd gnd FILL
XFILL_1__1374_ vdd gnd FILL
XFILL_4__1083_ vdd gnd FILL
XFILL_4__1419_ vdd gnd FILL
X_840_ _961_/B _891_/A vdd gnd INVX1
XFILL_2__1552_ vdd gnd FILL
XFILL_2__1483_ vdd gnd FILL
XFILL_2__1621_ vdd gnd FILL
XFILL_0__1050_ vdd gnd FILL
XFILL_1__921_ vdd gnd FILL
XFILL_1__852_ vdd gnd FILL
XFILL_3__1592_ vdd gnd FILL
XFILL_3__1661_ vdd gnd FILL
X_1043_ _1055_/B _1043_/B _1043_/C _1044_/A vdd gnd NAND3X1
X_969_ _993_/A _999_/A _992_/B vdd gnd NOR2X1
X_1112_ _1136_/C _1137_/B _1112_/C _1118_/B vdd gnd OAI21X1
XFILL_0__1317_ vdd gnd FILL
XFILL102450x66450 vdd gnd FILL
XFILL_0__1248_ vdd gnd FILL
XFILL_4__994_ vdd gnd FILL
XFILL_3__1026_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_4__1204_ vdd gnd FILL
XFILL_4__1135_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_0__870_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
XFILL_4__1066_ vdd gnd FILL
XFILL_2__1604_ vdd gnd FILL
XFILL_2__1535_ vdd gnd FILL
XFILL_2__1466_ vdd gnd FILL
XFILL_2__1397_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
X_1592_ _1592_/A _1592_/B _1592_/C _1599_/B vdd gnd AOI21X1
XFILL_0__999_ vdd gnd FILL
X_1661_ _1666_/A _1673_/A _1662_/B vdd gnd NAND2X1
XFILL_1__835_ vdd gnd FILL
XFILL_1__904_ vdd gnd FILL
XFILL102750x43050 vdd gnd FILL
XFILL_3__1575_ vdd gnd FILL
XFILL_3__1713_ vdd gnd FILL
XFILL_3__1644_ vdd gnd FILL
XFILL_1__1211_ vdd gnd FILL
X_1026_ _981_/A _981_/B _1424_/D _1513_/A _1079_/C vdd gnd AOI22X1
XFILL_3__1009_ vdd gnd FILL
XFILL_4__977_ vdd gnd FILL
XFILL_1__1073_ vdd gnd FILL
XFILL_1__1142_ vdd gnd FILL
XFILL_2__1320_ vdd gnd FILL
XFILL_2__1182_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_4__1049_ vdd gnd FILL
XFILL_2__1251_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_4__1118_ vdd gnd FILL
XFILL_0__853_ vdd gnd FILL
XFILL_0__1720_ vdd gnd FILL
XFILL_3__995_ vdd gnd FILL
XFILL_0__1651_ vdd gnd FILL
XFILL_4__900_ vdd gnd FILL
XFILL_3__1360_ vdd gnd FILL
XFILL_3__1291_ vdd gnd FILL
XFILL_2__1518_ vdd gnd FILL
XFILL_2__1449_ vdd gnd FILL
XFILL_0__1582_ vdd gnd FILL
XFILL_4__831_ vdd gnd FILL
X_1713_ _1723_/A rgb[0] vdd gnd BUFX2
XFILL_0__1016_ vdd gnd FILL
X_1575_ _1583_/A _1677_/A _1576_/B vdd gnd NOR2X1
X_1644_ _998_/A _997_/A _1672_/B _1646_/C vdd gnd OAI21X1
XFILL_3__1558_ vdd gnd FILL
XFILL_3__1627_ vdd gnd FILL
X_1009_ _1009_/A _1009_/B _1421_/B vdd gnd NAND2X1
XFILL_3__1489_ vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_4__1598_ vdd gnd FILL
XFILL_4__1667_ vdd gnd FILL
XFILL_2__1303_ vdd gnd FILL
XFILL_2__1165_ vdd gnd FILL
XFILL_0__905_ vdd gnd FILL
XFILL_2__1234_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
XFILL_0__836_ vdd gnd FILL
X_1360_ _1360_/A _1360_/B _1361_/C vdd gnd NOR2X1
XFILL_3__1412_ vdd gnd FILL
XFILL_3__1343_ vdd gnd FILL
XFILL_3__978_ vdd gnd FILL
XFILL_0__1634_ vdd gnd FILL
X_1291_ _1291_/A _1291_/B _1291_/C _1295_/B vdd gnd OAI21X1
XFILL_0__1565_ vdd gnd FILL
XFILL_0__1496_ vdd gnd FILL
XFILL_3__1274_ vdd gnd FILL
X_1558_ _1710_/Q _1677_/A vdd gnd INVX2
XFILL_4__1452_ vdd gnd FILL
X_1489_ _1489_/A _1489_/B _1490_/B vdd gnd NOR2X1
X_1627_ _1630_/C _1627_/B _1628_/A vdd gnd NOR2X1
XFILL_4__1521_ vdd gnd FILL
XFILL_4__1383_ vdd gnd FILL
XFILL_1__1674_ vdd gnd FILL
XFILL_2__996_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_3__901_ vdd gnd FILL
XFILL_3__832_ vdd gnd FILL
XFILL_4__1719_ vdd gnd FILL
XFILL_2__1217_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
XFILL_2__1079_ vdd gnd FILL
X_1412_ _1412_/A _1412_/B _1413_/C vdd gnd AND2X2
X_1343_ _1360_/B _1345_/A _1344_/B vdd gnd NOR2X1
XFILL_3__1326_ vdd gnd FILL
XFILL_0__1617_ vdd gnd FILL
X_1274_ _1687_/Q _1276_/D _1294_/A vdd gnd NAND2X1
XFILL_1__1390_ vdd gnd FILL
XFILL_3__1188_ vdd gnd FILL
XFILL_2__850_ vdd gnd FILL
XFILL_3__1257_ vdd gnd FILL
XFILL_0__1479_ vdd gnd FILL
XFILL_0__1548_ vdd gnd FILL
XFILL_4__1435_ vdd gnd FILL
XFILL_4__1504_ vdd gnd FILL
XFILL_4__1366_ vdd gnd FILL
XFILL_1__1588_ vdd gnd FILL
XFILL_4__1297_ vdd gnd FILL
XFILL_1__1657_ vdd gnd FILL
XFILL_2__1002_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
X_985_ _999_/A _985_/B _985_/C _996_/A vdd gnd NAND3X1
XFILL_3__1042_ vdd gnd FILL
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1402_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
XFILL_3__1111_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
X_1326_ _1650_/A _1351_/B _1351_/A _1412_/B vdd gnd NAND3X1
XFILL_1__997_ vdd gnd FILL
XFILL_1__1511_ vdd gnd FILL
X_1188_ _1315_/B _1315_/C _1355_/B vdd gnd NAND2X1
XFILL_4__1220_ vdd gnd FILL
XFILL_4__1151_ vdd gnd FILL
XFILL_1__1442_ vdd gnd FILL
XFILL_1__1373_ vdd gnd FILL
X_1257_ _1682_/Q _959_/A _1288_/C vdd gnd NAND2X1
XFILL_4__1082_ vdd gnd FILL
XFILL_3__1309_ vdd gnd FILL
XFILL_2__833_ vdd gnd FILL
XFILL_2__902_ vdd gnd FILL
XFILL_2__1620_ vdd gnd FILL
XFILL_2__1551_ vdd gnd FILL
XFILL_2__1482_ vdd gnd FILL
XFILL_4__1418_ vdd gnd FILL
XFILL_4__1349_ vdd gnd FILL
XFILL_1__920_ vdd gnd FILL
X_968_ _968_/A _974_/A vdd gnd INVX1
XFILL_1__851_ vdd gnd FILL
XFILL_3__1591_ vdd gnd FILL
XFILL_3__1660_ vdd gnd FILL
X_1042_ _1055_/A _1055_/C _1043_/C vdd gnd NOR2X1
X_899_ _956_/Q _899_/B _934_/A vdd gnd NOR2X1
XFILL_4__993_ vdd gnd FILL
X_1111_ _1111_/A _1112_/C _1137_/B vdd gnd NAND2X1
XFILL_0__1316_ vdd gnd FILL
XFILL_0__1247_ vdd gnd FILL
XFILL_3__1025_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
X_1309_ _1678_/Q _1408_/C vdd gnd INVX1
XFILL_1__1356_ vdd gnd FILL
XFILL_4__1203_ vdd gnd FILL
XFILL_1__1425_ vdd gnd FILL
XFILL_4__1065_ vdd gnd FILL
XFILL_4__1134_ vdd gnd FILL
XFILL_1__1287_ vdd gnd FILL
XFILL_2__1603_ vdd gnd FILL
XFILL_2__1534_ vdd gnd FILL
XFILL_2__1396_ vdd gnd FILL
XFILL_2__1465_ vdd gnd FILL
XFILL_0__1032_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
XFILL_3__1712_ vdd gnd FILL
X_1591_ _1591_/A _1591_/B _1592_/B vdd gnd AND2X2
X_1660_ _1673_/A _1666_/A _1665_/C vdd gnd OR2X2
XFILL_1__903_ vdd gnd FILL
XFILL_1__834_ vdd gnd FILL
XFILL_3__1643_ vdd gnd FILL
XFILL_3__1574_ vdd gnd FILL
XFILL_1__1210_ vdd gnd FILL
XFILL_1__1141_ vdd gnd FILL
X_1025_ _980_/B _1707_/Q _1424_/D vdd gnd XOR2X1
XFILL_4__976_ vdd gnd FILL
XFILL_3__1008_ vdd gnd FILL
XFILL_1__1072_ vdd gnd FILL
XFILL_2__1250_ vdd gnd FILL
XFILL_0__921_ vdd gnd FILL
XFILL_0__852_ vdd gnd FILL
XFILL_2__1181_ vdd gnd FILL
XFILL_4__1048_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_4__1117_ vdd gnd FILL
XFILL_1__1408_ vdd gnd FILL
XFILL_3__994_ vdd gnd FILL
XFILL_0__1650_ vdd gnd FILL
XFILL_4__830_ vdd gnd FILL
XFILL_2__1379_ vdd gnd FILL
XFILL_0__1581_ vdd gnd FILL
XFILL_2__1517_ vdd gnd FILL
XFILL_3__1290_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
X_1712_ _858_/Y p_tick vdd gnd BUFX2
XFILL_0__1015_ vdd gnd FILL
X_1643_ _1649_/A _1655_/C _1654_/B vdd gnd NAND2X1
X_1574_ _1694_/Q _1710_/Q _1576_/A vdd gnd NOR2X1
XFILL_3__1557_ vdd gnd FILL
XFILL_3__1488_ vdd gnd FILL
XFILL_3__1626_ vdd gnd FILL
X_1008_ _1650_/A _992_/B _972_/B _1009_/A vdd gnd NAND3X1
XFILL_4__959_ vdd gnd FILL
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL_4__1597_ vdd gnd FILL
XFILL_4__1666_ vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_2__1302_ vdd gnd FILL
XFILL_0__835_ vdd gnd FILL
XFILL_0__904_ vdd gnd FILL
XFILL_2__1164_ vdd gnd FILL
XFILL_2__1095_ vdd gnd FILL
XFILL_3__977_ vdd gnd FILL
XFILL_3__1411_ vdd gnd FILL
XFILL_3__1342_ vdd gnd FILL
XFILL_0__1564_ vdd gnd FILL
XFILL_0__1633_ vdd gnd FILL
X_1290_ _1298_/C _1290_/B _1290_/C _1296_/B vdd gnd AOI21X1
XFILL_3__1273_ vdd gnd FILL
XFILL_0__1495_ vdd gnd FILL
X_1626_ _984_/B _1671_/C _1630_/C vdd gnd NOR2X1
XFILL_3__1609_ vdd gnd FILL
X_1557_ _1692_/Q _1710_/Q _1560_/A vdd gnd NOR2X1
XFILL_1__1673_ vdd gnd FILL
X_1488_ _1488_/A _1488_/B _1536_/B vdd gnd NAND2X1
XFILL_4__1451_ vdd gnd FILL
XFILL_4__1520_ vdd gnd FILL
XFILL_4__1382_ vdd gnd FILL
XFILL_2__995_ vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_4__1718_ vdd gnd FILL
XFILL_3__831_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_3__900_ vdd gnd FILL
XFILL_4__1649_ vdd gnd FILL
XFILL_2__1216_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_2__1147_ vdd gnd FILL
XFILL_2__1078_ vdd gnd FILL
X_1411_ _971_/A _1411_/B _1413_/A vdd gnd NAND2X1
X_1342_ _997_/A _1342_/B _1360_/B vdd gnd NOR2X1
X_1273_ _1513_/A _1698_/Q _1689_/Q _965_/C _1303_/A vdd gnd AOI22X1
XFILL_3__1325_ vdd gnd FILL
XFILL_0__1616_ vdd gnd FILL
XFILL_0__1547_ vdd gnd FILL
XFILL_3__1256_ vdd gnd FILL
XFILL_3__1187_ vdd gnd FILL
XFILL_4_BUFX2_insert0 vdd gnd FILL
XFILL_0__1478_ vdd gnd FILL
X_1609_ _1674_/C _1655_/A _1609_/C _1623_/B vdd gnd NAND3X1
XFILL_1__1725_ vdd gnd FILL
XFILL_4__1365_ vdd gnd FILL
XFILL_1__1656_ vdd gnd FILL
XFILL_4__1434_ vdd gnd FILL
XFILL_4__1503_ vdd gnd FILL
XFILL_2__1001_ vdd gnd FILL
XFILL_1__1587_ vdd gnd FILL
XFILL_4__1296_ vdd gnd FILL
XFILL_2__978_ vdd gnd FILL
X_984_ _986_/A _984_/B _985_/C vdd gnd NAND2X1
XFILL_0__1401_ vdd gnd FILL
XFILL_3__1110_ vdd gnd FILL
XFILL103050x85950 vdd gnd FILL
XFILL_3__1041_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
XFILL_0__1332_ vdd gnd FILL
XFILL_0__1263_ vdd gnd FILL
X_1325_ _1573_/A _1406_/A _1583_/A _1351_/A vdd gnd OAI21X1
XFILL_1__996_ vdd gnd FILL
XFILL_1__1510_ vdd gnd FILL
X_1256_ _957_/A _1390_/B _1259_/C vdd gnd NAND2X1
X_1187_ _1403_/B _1351_/B _1599_/A _1315_/C vdd gnd OAI21X1
XFILL_4__1150_ vdd gnd FILL
XFILL_2__901_ vdd gnd FILL
XFILL_1__1441_ vdd gnd FILL
XFILL_1__1372_ vdd gnd FILL
XFILL_3__1308_ vdd gnd FILL
XFILL_4__1081_ vdd gnd FILL
XFILL_3__1239_ vdd gnd FILL
XFILL_2__832_ vdd gnd FILL
XFILL_4__1348_ vdd gnd FILL
XFILL_4__1417_ vdd gnd FILL
XFILL_1__1639_ vdd gnd FILL
XFILL_2__1481_ vdd gnd FILL
XFILL_2__1550_ vdd gnd FILL
XFILL_4__1279_ vdd gnd FILL
X_898_ _933_/C _898_/B _936_/A _899_/B vdd gnd OAI21X1
XFILL_1__850_ vdd gnd FILL
XFILL103350x62550 vdd gnd FILL
X_967_ _967_/A _967_/B _967_/Y vdd gnd NAND2X1
XFILL_3__1590_ vdd gnd FILL
X_1110_ _962_/A _1110_/B _1111_/A vdd gnd NAND2X1
X_1041_ _953_/Q _1655_/A _1055_/C vdd gnd NOR2X1
XFILL_4__992_ vdd gnd FILL
XFILL_0__1177_ vdd gnd FILL
XFILL_0__1315_ vdd gnd FILL
XFILL_3__1024_ vdd gnd FILL
XFILL_0__1246_ vdd gnd FILL
XFILL_4__1202_ vdd gnd FILL
XFILL_1__1424_ vdd gnd FILL
XFILL_1__979_ vdd gnd FILL
X_1308_ reset _1308_/Y vdd gnd INVX8
X_1239_ _1681_/Q _1298_/B _1288_/A vdd gnd NOR2X1
XFILL_1__1355_ vdd gnd FILL
XFILL_4__1064_ vdd gnd FILL
XFILL_4__1133_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
XFILL_2__1602_ vdd gnd FILL
XFILL_2__1533_ vdd gnd FILL
XFILL_2__1395_ vdd gnd FILL
XFILL_2__1464_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
XFILL_1__902_ vdd gnd FILL
XFILL_3__1711_ vdd gnd FILL
XFILL_3__1642_ vdd gnd FILL
X_1590_ _1590_/A _1592_/C vdd gnd INVX1
XFILL_1__833_ vdd gnd FILL
X_1024_ _956_/Q _1513_/A vdd gnd INVX2
XFILL_3__1573_ vdd gnd FILL
XFILL_4__975_ vdd gnd FILL
XFILL_1__1140_ vdd gnd FILL
XFILL_0__1229_ vdd gnd FILL
XFILL_3__1007_ vdd gnd FILL
XFILL_1__1071_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_4__1116_ vdd gnd FILL
XFILL_0__920_ vdd gnd FILL
XFILL_0__851_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_4__1047_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_3__993_ vdd gnd FILL
XFILL_2__1516_ vdd gnd FILL
XFILL_0__1580_ vdd gnd FILL
XFILL_2__1378_ vdd gnd FILL
XFILL_2__1447_ vdd gnd FILL
X_1711_ _850_/Y hsync vdd gnd BUFX2
XFILL_0__1014_ vdd gnd FILL
X_1642_ _971_/B _1672_/B _1655_/C vdd gnd NAND2X1
X_1573_ _1573_/A _1573_/B _1573_/C _1693_/D vdd gnd AOI21X1
XFILL_3__1625_ vdd gnd FILL
X_1007_ _1015_/B _1009_/B vdd gnd INVX1
XFILL_3__1556_ vdd gnd FILL
XFILL_3__1487_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_4__889_ vdd gnd FILL
XFILL_4__958_ vdd gnd FILL
XFILL_1__1123_ vdd gnd FILL
XFILL_4__1596_ vdd gnd FILL
XFILL_4__1665_ vdd gnd FILL
XFILL_2__1163_ vdd gnd FILL
XFILL_2__1232_ vdd gnd FILL
XFILL_2__1301_ vdd gnd FILL
XFILL_0__903_ vdd gnd FILL
XFILL_0__834_ vdd gnd FILL
XFILL_2__1094_ vdd gnd FILL
XFILL_3__976_ vdd gnd FILL
XFILL_3__1341_ vdd gnd FILL
XFILL_3__1272_ vdd gnd FILL
XFILL_0__1632_ vdd gnd FILL
XFILL_3__1410_ vdd gnd FILL
XFILL_0__1563_ vdd gnd FILL
XFILL_0__1494_ vdd gnd FILL
X_1556_ _1556_/A _1676_/A _1556_/C _1564_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert11 vdd gnd FILL
X_1625_ _1630_/A _1627_/B vdd gnd INVX1
XFILL_4__1381_ vdd gnd FILL
XFILL_3__1608_ vdd gnd FILL
XFILL_1__1672_ vdd gnd FILL
X_1487_ _1487_/A _1501_/A _1536_/C vdd gnd NAND2X1
XFILL_3__1539_ vdd gnd FILL
XFILL_4__1450_ vdd gnd FILL
XFILL_2__994_ vdd gnd FILL
XFILL_1__1037_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_3__830_ vdd gnd FILL
XFILL_4__1648_ vdd gnd FILL
XFILL_4__1717_ vdd gnd FILL
XFILL_4__1579_ vdd gnd FILL
XFILL_2__1215_ vdd gnd FILL
XFILL_2__1146_ vdd gnd FILL
XFILL_2__1077_ vdd gnd FILL
XFILL_0_CLKBUF1_insert4 vdd gnd FILL
X_1410_ _1545_/A _1410_/B _1432_/A vdd gnd NAND2X1
X_1341_ _1363_/A _1341_/B _1364_/C _1344_/A vdd gnd OAI21X1
XFILL_3__959_ vdd gnd FILL
X_1272_ _964_/A _1397_/B _1303_/C vdd gnd NAND2X1
XFILL_3__1324_ vdd gnd FILL
XFILL_3__1255_ vdd gnd FILL
XFILL_0__1615_ vdd gnd FILL
XFILL_0__1477_ vdd gnd FILL
XFILL_0__1546_ vdd gnd FILL
XFILL_3__1186_ vdd gnd FILL
XFILL_4_BUFX2_insert1 vdd gnd FILL
X_1608_ _971_/B _998_/A _1609_/C vdd gnd NOR2X1
X_1539_ _1539_/A _1621_/A _1540_/C vdd gnd OR2X2
XFILL_4__1502_ vdd gnd FILL
XFILL_1__1724_ vdd gnd FILL
XFILL_4__1364_ vdd gnd FILL
XFILL_1__1655_ vdd gnd FILL
XFILL_4__1433_ vdd gnd FILL
XFILL_4__1295_ vdd gnd FILL
XFILL_1__1586_ vdd gnd FILL
XFILL_2__1000_ vdd gnd FILL
XFILL_2__977_ vdd gnd FILL
X_983_ _993_/A _984_/B vdd gnd INVX2
XFILL_0__1400_ vdd gnd FILL
XFILL_3__1040_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
XFILL_0__1262_ vdd gnd FILL
XFILL_2__1129_ vdd gnd FILL
X_1186_ _1327_/B _1327_/C _1411_/B vdd gnd NAND2X1
X_1324_ _1324_/A _1324_/B _971_/B _1412_/A vdd gnd OAI21X1
XFILL_1__1440_ vdd gnd FILL
XFILL_1__995_ vdd gnd FILL
X_1255_ _1265_/A _1267_/B _1267_/C _1264_/C vdd gnd NAND3X1
XFILL_3__1169_ vdd gnd FILL
XFILL_2__831_ vdd gnd FILL
XFILL_2__900_ vdd gnd FILL
XFILL_4__1080_ vdd gnd FILL
XFILL_1__1371_ vdd gnd FILL
XFILL_0__1529_ vdd gnd FILL
XFILL_3__1307_ vdd gnd FILL
XFILL_3__1238_ vdd gnd FILL
XFILL_4__1416_ vdd gnd FILL
XFILL_4__1347_ vdd gnd FILL
XFILL_1__1569_ vdd gnd FILL
XFILL_4__1278_ vdd gnd FILL
XFILL_2__1480_ vdd gnd FILL
XFILL_1__1638_ vdd gnd FILL
XFILL103950x11850 vdd gnd FILL
XFILL103650x46950 vdd gnd FILL
X_1040_ _952_/Q _1650_/A _1055_/A vdd gnd NOR2X1
X_897_ _968_/A _933_/C vdd gnd INVX1
X_966_ _966_/A _966_/B _967_/B vdd gnd NOR2X1
XFILL_3__1023_ vdd gnd FILL
XFILL_4__991_ vdd gnd FILL
XFILL_0__1314_ vdd gnd FILL
XFILL_0__1176_ vdd gnd FILL
XFILL_0__1245_ vdd gnd FILL
X_1169_ _990_/A _1342_/B _1175_/C vdd gnd NOR2X1
XFILL_4__1201_ vdd gnd FILL
XFILL_1__1423_ vdd gnd FILL
XFILL_1__978_ vdd gnd FILL
X_1307_ _1307_/A _1307_/B _1721_/A vdd gnd NOR2X1
XFILL_4__1132_ vdd gnd FILL
X_1238_ _960_/A _1298_/B vdd gnd INVX1
XFILL_1__1354_ vdd gnd FILL
XFILL_4__1063_ vdd gnd FILL
XFILL_1__1285_ vdd gnd FILL
XFILL_2__1601_ vdd gnd FILL
XFILL_2__1532_ vdd gnd FILL
XFILL_2__1463_ vdd gnd FILL
XFILL_3_CLKBUF1_insert10 vdd gnd FILL
XFILL_2__1394_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL103650x58650 vdd gnd FILL
XFILL_1__832_ vdd gnd FILL
XFILL_1__901_ vdd gnd FILL
XFILL_3__1641_ vdd gnd FILL
XFILL_3__1572_ vdd gnd FILL
X_949_ _949_/D vdd _956_/R _949_/CLK _986_/A vdd gnd DFFSR
X_1023_ _1078_/A _974_/Y _981_/Y _1074_/A vdd gnd AOI21X1
XFILL_0__1228_ vdd gnd FILL
XFILL_3__1006_ vdd gnd FILL
XFILL_4__974_ vdd gnd FILL
XFILL_1__1070_ vdd gnd FILL
XFILL_0__1159_ vdd gnd FILL
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_4__1115_ vdd gnd FILL
XFILL_0__850_ vdd gnd FILL
XFILL_4__1046_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_3__992_ vdd gnd FILL
XFILL_2__1446_ vdd gnd FILL
XFILL_2__1515_ vdd gnd FILL
XFILL103950x35250 vdd gnd FILL
XFILL_2__1377_ vdd gnd FILL
XFILL_0__1013_ vdd gnd FILL
XFILL_0__979_ vdd gnd FILL
X_1710_ _1710_/D vdd _1710_/R _1710_/CLK _1710_/Q vdd gnd DFFSR
X_1641_ _1657_/A _1657_/B _1650_/A _1649_/A vdd gnd OAI21X1
X_1572_ _1572_/A _1572_/B _1572_/C _1573_/C vdd gnd AOI21X1
XFILL_3__1555_ vdd gnd FILL
XFILL_3__1624_ vdd gnd FILL
X_1006_ _992_/B _972_/B _1650_/A _1015_/B vdd gnd AOI21X1
XFILL_3__1486_ vdd gnd FILL
XFILL_1__1053_ vdd gnd FILL
XFILL_4__888_ vdd gnd FILL
XFILL_4__957_ vdd gnd FILL
XFILL_1__1122_ vdd gnd FILL
XFILL_4__1664_ vdd gnd FILL
XFILL_4__1595_ vdd gnd FILL
XFILL_2__1300_ vdd gnd FILL
XFILL_0__902_ vdd gnd FILL
XFILL_2__1162_ vdd gnd FILL
XFILL_2__1231_ vdd gnd FILL
XFILL_4__1029_ vdd gnd FILL
XFILL_2__1093_ vdd gnd FILL
XFILL_0__833_ vdd gnd FILL
XFILL_3__975_ vdd gnd FILL
XFILL_3__1340_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL_3__1271_ vdd gnd FILL
XFILL_0__1631_ vdd gnd FILL
XFILL_0__1493_ vdd gnd FILL
XFILL_0__1562_ vdd gnd FILL
XFILL102450x62550 vdd gnd FILL
XFILL_2_BUFX2_insert12 vdd gnd FILL
X_1555_ _1555_/A _1555_/B _1556_/C vdd gnd NAND2X1
X_1624_ _1657_/A _1657_/B _984_/B _1630_/A vdd gnd OAI21X1
XFILL_4__1380_ vdd gnd FILL
XFILL_3__1607_ vdd gnd FILL
XFILL_1__1671_ vdd gnd FILL
X_1486_ _1488_/B _1501_/A vdd gnd INVX1
XFILL_3__1538_ vdd gnd FILL
XFILL_2__993_ vdd gnd FILL
XFILL_3__1469_ vdd gnd FILL
XFILL_1__1036_ vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_4__1716_ vdd gnd FILL
XFILL_4__1647_ vdd gnd FILL
XFILL_4__1578_ vdd gnd FILL
XFILL_2__1214_ vdd gnd FILL
XFILL_2__1145_ vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
XFILL_0_CLKBUF1_insert5 vdd gnd FILL
X_1340_ _1690_/Q _999_/A _1363_/A vdd gnd NOR2X1
XFILL_0__1614_ vdd gnd FILL
XFILL_3__889_ vdd gnd FILL
XFILL_3__958_ vdd gnd FILL
X_1271_ _1428_/A _1397_/B vdd gnd INVX1
XFILL_3__1185_ vdd gnd FILL
XFILL_3__1323_ vdd gnd FILL
XFILL_4_BUFX2_insert2 vdd gnd FILL
XFILL_3__1254_ vdd gnd FILL
XFILL_0__1476_ vdd gnd FILL
XFILL_0__1545_ vdd gnd FILL
X_1607_ _992_/A _984_/B _1672_/A _1623_/A vdd gnd NAND3X1
XFILL_4__1501_ vdd gnd FILL
X_1469_ _1686_/Q _1685_/Q _1680_/Q _1499_/A vdd gnd OAI21X1
XFILL_1__1723_ vdd gnd FILL
X_1538_ _1602_/C _1621_/A vdd gnd INVX1
XFILL_4__1432_ vdd gnd FILL
XFILL_4__1363_ vdd gnd FILL
XFILL_1__1654_ vdd gnd FILL
XFILL_1__1585_ vdd gnd FILL
XFILL_4__1294_ vdd gnd FILL
XFILL_2__976_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
X_982_ _982_/A _985_/B vdd gnd INVX1
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1261_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_2__1059_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
X_1323_ _1414_/A _1414_/B _1346_/C vdd gnd NOR2X1
XFILL_1__994_ vdd gnd FILL
X_1185_ _1185_/A _1185_/B _1193_/A vdd gnd NAND2X1
X_1254_ _1254_/A _1254_/B _1254_/C _1267_/C vdd gnd OAI21X1
XFILL_3__1306_ vdd gnd FILL
XFILL_1__1370_ vdd gnd FILL
XFILL_2__830_ vdd gnd FILL
XFILL_0__1528_ vdd gnd FILL
XFILL_3__1237_ vdd gnd FILL
XFILL_3__1168_ vdd gnd FILL
XFILL_0__1459_ vdd gnd FILL
XFILL_3__1099_ vdd gnd FILL
XFILL_4__1346_ vdd gnd FILL
XFILL_1__1568_ vdd gnd FILL
XFILL_1__1637_ vdd gnd FILL
XFILL_1__1499_ vdd gnd FILL
XFILL_4__1277_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
X_965_ _965_/A _965_/B _965_/C _966_/B vdd gnd OAI21X1
X_896_ _982_/A _901_/A vdd gnd INVX1
XFILL_2__1677_ vdd gnd FILL
XFILL_4__990_ vdd gnd FILL
XFILL_0__1244_ vdd gnd FILL
XFILL_3__1022_ vdd gnd FILL
XFILL_0__1313_ vdd gnd FILL
XFILL_0__1175_ vdd gnd FILL
X_1306_ _1306_/A _1307_/A _1306_/C _1724_/A vdd gnd AOI21X1
XFILL_1__977_ vdd gnd FILL
XFILL_1__1353_ vdd gnd FILL
X_1237_ _1237_/A _1237_/B _1304_/A vdd gnd NOR2X1
X_1168_ _1332_/B _1332_/A _1342_/B vdd gnd AND2X2
XFILL_4__1200_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
XFILL_4__1062_ vdd gnd FILL
XFILL_4__1131_ vdd gnd FILL
X_1099_ _1099_/A _1099_/B _1099_/C _1138_/C vdd gnd AOI21X1
XFILL_1__1284_ vdd gnd FILL
XFILL_2__1600_ vdd gnd FILL
XFILL_2__1531_ vdd gnd FILL
XFILL_2__1462_ vdd gnd FILL
XFILL_4__1329_ vdd gnd FILL
XFILL_2__1393_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
XFILL_1__831_ vdd gnd FILL
XFILL_1__900_ vdd gnd FILL
X_948_ _948_/D vdd _948_/R _949_/CLK _982_/A vdd gnd DFFSR
XFILL_3__1571_ vdd gnd FILL
XFILL_3__1640_ vdd gnd FILL
X_1022_ _1022_/A _1022_/B _1078_/A vdd gnd NAND2X1
XFILL_4__973_ vdd gnd FILL
X_879_ _962_/B _886_/B vdd gnd INVX1
XFILL_0__1227_ vdd gnd FILL
XFILL_3__1005_ vdd gnd FILL
XFILL_0__1158_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_4__1045_ vdd gnd FILL
XFILL_4__1114_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_3__991_ vdd gnd FILL
XFILL_2__1376_ vdd gnd FILL
XFILL_2__1514_ vdd gnd FILL
XFILL_2__1445_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
XFILL_0__1012_ vdd gnd FILL
X_1571_ _1572_/B _1572_/A _1602_/C _1572_/C vdd gnd OAI21X1
X_1640_ _1640_/A _998_/Y _1670_/B _1702_/D vdd gnd MUX2X1
XFILL_3__1623_ vdd gnd FILL
XFILL_3__1485_ vdd gnd FILL
XFILL_3__1554_ vdd gnd FILL
X_1005_ _971_/B _1650_/A vdd gnd INVX2
XFILL_1__1121_ vdd gnd FILL
XFILL_1__1052_ vdd gnd FILL
XFILL_4__887_ vdd gnd FILL
XFILL_4__1594_ vdd gnd FILL
XFILL_4__1663_ vdd gnd FILL
XFILL_2__1230_ vdd gnd FILL
XFILL_2__1161_ vdd gnd FILL
XFILL_0__832_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_0__901_ vdd gnd FILL
XFILL_4__1028_ vdd gnd FILL
XFILL_2__1092_ vdd gnd FILL
XFILL_3__974_ vdd gnd FILL
XFILL_0__1630_ vdd gnd FILL
XFILL_2__1359_ vdd gnd FILL
XFILL_3__1270_ vdd gnd FILL
XFILL_2__1428_ vdd gnd FILL
XFILL_0__1561_ vdd gnd FILL
XFILL_0__1492_ vdd gnd FILL
XFILL102750x46950 vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
X_1623_ _1623_/A _1623_/B _1657_/B vdd gnd NOR2X1
X_1485_ _1485_/A _1485_/B _1539_/A vdd gnd XNOR2X1
X_1554_ _1709_/Q _1676_/A vdd gnd INVX1
.ends

